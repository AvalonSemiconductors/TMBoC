magic
tech sky130B
magscale 1 2
timestamp 1681305957
<< metal1 >>
rect 397454 700816 397460 700868
rect 397512 700856 397518 700868
rect 445018 700856 445024 700868
rect 397512 700828 445024 700856
rect 397512 700816 397518 700828
rect 445018 700816 445024 700828
rect 445076 700816 445082 700868
rect 364978 700748 364984 700800
rect 365036 700788 365042 700800
rect 446490 700788 446496 700800
rect 365036 700760 446496 700788
rect 365036 700748 365042 700760
rect 446490 700748 446496 700760
rect 446548 700748 446554 700800
rect 332502 700680 332508 700732
rect 332560 700720 332566 700732
rect 444098 700720 444104 700732
rect 332560 700692 444104 700720
rect 332560 700680 332566 700692
rect 444098 700680 444104 700692
rect 444156 700680 444162 700732
rect 218974 700612 218980 700664
rect 219032 700652 219038 700664
rect 418798 700652 418804 700664
rect 219032 700624 418804 700652
rect 219032 700612 219038 700624
rect 418798 700612 418804 700624
rect 418856 700612 418862 700664
rect 235166 700544 235172 700596
rect 235224 700584 235230 700596
rect 446398 700584 446404 700596
rect 235224 700556 446404 700584
rect 235224 700544 235230 700556
rect 446398 700544 446404 700556
rect 446456 700544 446462 700596
rect 202782 700476 202788 700528
rect 202840 700516 202846 700528
rect 446582 700516 446588 700528
rect 202840 700488 446588 700516
rect 202840 700476 202846 700488
rect 446582 700476 446588 700488
rect 446640 700476 446646 700528
rect 154114 700408 154120 700460
rect 154172 700448 154178 700460
rect 418890 700448 418896 700460
rect 154172 700420 418896 700448
rect 154172 700408 154178 700420
rect 418890 700408 418896 700420
rect 418948 700408 418954 700460
rect 447870 700408 447876 700460
rect 447928 700448 447934 700460
rect 478506 700448 478512 700460
rect 447928 700420 478512 700448
rect 447928 700408 447934 700420
rect 478506 700408 478512 700420
rect 478564 700408 478570 700460
rect 170306 700340 170312 700392
rect 170364 700380 170370 700392
rect 449158 700380 449164 700392
rect 170364 700352 449164 700380
rect 170364 700340 170370 700352
rect 449158 700340 449164 700352
rect 449216 700340 449222 700392
rect 40494 700272 40500 700324
rect 40552 700312 40558 700324
rect 446674 700312 446680 700324
rect 40552 700284 446680 700312
rect 40552 700272 40558 700284
rect 446674 700272 446680 700284
rect 446732 700272 446738 700324
rect 447962 700272 447968 700324
rect 448020 700312 448026 700324
rect 494790 700312 494796 700324
rect 448020 700284 494796 700312
rect 448020 700272 448026 700284
rect 494790 700272 494796 700284
rect 494848 700272 494854 700324
rect 576118 696940 576124 696992
rect 576176 696980 576182 696992
rect 580166 696980 580172 696992
rect 576176 696952 580172 696980
rect 576176 696940 576182 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 300118 690616 300124 690668
rect 300176 690656 300182 690668
rect 449250 690656 449256 690668
rect 300176 690628 449256 690656
rect 300176 690616 300182 690628
rect 449250 690616 449256 690628
rect 449308 690616 449314 690668
rect 348786 687896 348792 687948
rect 348844 687936 348850 687948
rect 445110 687936 445116 687948
rect 348844 687908 445116 687936
rect 348844 687896 348850 687908
rect 445110 687896 445116 687908
rect 445168 687896 445174 687948
rect 8110 686468 8116 686520
rect 8168 686508 8174 686520
rect 445202 686508 445208 686520
rect 8168 686480 445208 686508
rect 8168 686468 8174 686480
rect 445202 686468 445208 686480
rect 445260 686468 445266 686520
rect 267642 685244 267648 685296
rect 267700 685284 267706 685296
rect 418982 685284 418988 685296
rect 267700 685256 418988 685284
rect 267700 685244 267706 685256
rect 418982 685244 418988 685256
rect 419040 685244 419046 685296
rect 89162 685176 89168 685228
rect 89220 685216 89226 685228
rect 416038 685216 416044 685228
rect 89220 685188 416044 685216
rect 89220 685176 89226 685188
rect 416038 685176 416044 685188
rect 416096 685176 416102 685228
rect 72970 685108 72976 685160
rect 73028 685148 73034 685160
rect 445294 685148 445300 685160
rect 73028 685120 445300 685148
rect 73028 685108 73034 685120
rect 445294 685108 445300 685120
rect 445352 685108 445358 685160
rect 3786 684632 3792 684684
rect 3844 684672 3850 684684
rect 420270 684672 420276 684684
rect 3844 684644 420276 684672
rect 3844 684632 3850 684644
rect 420270 684632 420276 684644
rect 420328 684632 420334 684684
rect 3418 684564 3424 684616
rect 3476 684604 3482 684616
rect 420178 684604 420184 684616
rect 3476 684576 420184 684604
rect 3476 684564 3482 684576
rect 420178 684564 420184 684576
rect 420236 684564 420242 684616
rect 3970 684496 3976 684548
rect 4028 684536 4034 684548
rect 446858 684536 446864 684548
rect 4028 684508 446864 684536
rect 4028 684496 4034 684508
rect 446858 684496 446864 684508
rect 446916 684496 446922 684548
rect 24118 683680 24124 683732
rect 24176 683720 24182 683732
rect 359458 683720 359464 683732
rect 24176 683692 359464 683720
rect 24176 683680 24182 683692
rect 359458 683680 359464 683692
rect 359516 683680 359522 683732
rect 21450 683612 21456 683664
rect 21508 683652 21514 683664
rect 420822 683652 420828 683664
rect 21508 683624 420828 683652
rect 21508 683612 21514 683624
rect 420822 683612 420828 683624
rect 420880 683612 420886 683664
rect 3878 683544 3884 683596
rect 3936 683584 3942 683596
rect 420362 683584 420368 683596
rect 3936 683556 420368 683584
rect 3936 683544 3942 683556
rect 420362 683544 420368 683556
rect 420420 683544 420426 683596
rect 3602 683476 3608 683528
rect 3660 683516 3666 683528
rect 420638 683516 420644 683528
rect 3660 683488 420644 683516
rect 3660 683476 3666 683488
rect 420638 683476 420644 683488
rect 420696 683476 420702 683528
rect 3694 683408 3700 683460
rect 3752 683448 3758 683460
rect 420730 683448 420736 683460
rect 3752 683420 420736 683448
rect 3752 683408 3758 683420
rect 420730 683408 420736 683420
rect 420788 683408 420794 683460
rect 3326 683340 3332 683392
rect 3384 683380 3390 683392
rect 420546 683380 420552 683392
rect 3384 683352 420552 683380
rect 3384 683340 3390 683352
rect 420546 683340 420552 683352
rect 420604 683340 420610 683392
rect 21358 683272 21364 683324
rect 21416 683312 21422 683324
rect 445478 683312 445484 683324
rect 21416 683284 445484 683312
rect 21416 683272 21422 683284
rect 445478 683272 445484 683284
rect 445536 683272 445542 683324
rect 3510 683204 3516 683256
rect 3568 683244 3574 683256
rect 445386 683244 445392 683256
rect 3568 683216 445392 683244
rect 3568 683204 3574 683216
rect 445386 683204 445392 683216
rect 445444 683204 445450 683256
rect 4062 683136 4068 683188
rect 4120 683176 4126 683188
rect 447042 683176 447048 683188
rect 4120 683148 447048 683176
rect 4120 683136 4126 683148
rect 447042 683136 447048 683148
rect 447100 683136 447106 683188
rect 11054 682728 11060 682780
rect 11112 682768 11118 682780
rect 24118 682768 24124 682780
rect 11112 682740 24124 682768
rect 11112 682728 11118 682740
rect 24118 682728 24124 682740
rect 24176 682728 24182 682780
rect 3234 682660 3240 682712
rect 3292 682700 3298 682712
rect 446306 682700 446312 682712
rect 3292 682672 446312 682700
rect 3292 682660 3298 682672
rect 446306 682660 446312 682672
rect 446364 682660 446370 682712
rect 6914 675792 6920 675844
rect 6972 675832 6978 675844
rect 10962 675832 10968 675844
rect 6972 675804 10968 675832
rect 6972 675792 6978 675804
rect 10962 675792 10968 675804
rect 11020 675792 11026 675844
rect 359458 672052 359464 672104
rect 359516 672092 359522 672104
rect 360838 672092 360844 672104
rect 359516 672064 360844 672092
rect 359516 672052 359522 672064
rect 360838 672052 360844 672064
rect 360896 672052 360902 672104
rect 447778 669944 447784 669996
rect 447836 669984 447842 669996
rect 462314 669984 462320 669996
rect 447836 669956 462320 669984
rect 447836 669944 447842 669956
rect 462314 669944 462320 669956
rect 462372 669944 462378 669996
rect 4798 667904 4804 667956
rect 4856 667944 4862 667956
rect 6822 667944 6828 667956
rect 4856 667916 6828 667944
rect 4856 667904 4862 667916
rect 6822 667904 6828 667916
rect 6880 667904 6886 667956
rect 361758 667904 361764 667956
rect 361816 667944 361822 667956
rect 378778 667944 378784 667956
rect 361816 667916 378784 667944
rect 361816 667904 361822 667916
rect 378778 667904 378784 667916
rect 378836 667904 378842 667956
rect 361758 656888 361764 656940
rect 361816 656928 361822 656940
rect 376018 656928 376024 656940
rect 361816 656900 376024 656928
rect 361816 656888 361822 656900
rect 376018 656888 376024 656900
rect 376076 656888 376082 656940
rect 3510 656140 3516 656192
rect 3568 656180 3574 656192
rect 20898 656180 20904 656192
rect 3568 656152 20904 656180
rect 3568 656140 3574 656152
rect 20898 656140 20904 656152
rect 20956 656140 20962 656192
rect 361758 645872 361764 645924
rect 361816 645912 361822 645924
rect 374730 645912 374736 645924
rect 361816 645884 374736 645912
rect 361816 645872 361822 645884
rect 374730 645872 374736 645884
rect 374788 645872 374794 645924
rect 571978 643084 571984 643136
rect 572036 643124 572042 643136
rect 580166 643124 580172 643136
rect 572036 643096 580172 643124
rect 572036 643084 572042 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 361574 634788 361580 634840
rect 361632 634828 361638 634840
rect 400858 634828 400864 634840
rect 361632 634800 400864 634828
rect 361632 634788 361638 634800
rect 400858 634788 400864 634800
rect 400916 634788 400922 634840
rect 3142 633360 3148 633412
rect 3200 633400 3206 633412
rect 20898 633400 20904 633412
rect 3200 633372 20904 633400
rect 3200 633360 3206 633372
rect 20898 633360 20904 633372
rect 20956 633360 20962 633412
rect 574738 630640 574744 630692
rect 574796 630680 574802 630692
rect 580166 630680 580172 630692
rect 574796 630652 580172 630680
rect 574796 630640 574802 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 361574 623772 361580 623824
rect 361632 623812 361638 623824
rect 371878 623812 371884 623824
rect 361632 623784 371884 623812
rect 361632 623772 361638 623784
rect 371878 623772 371884 623784
rect 371936 623772 371942 623824
rect 570598 616836 570604 616888
rect 570656 616876 570662 616888
rect 580166 616876 580172 616888
rect 570656 616848 580172 616876
rect 570656 616836 570662 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 361574 612824 361580 612876
rect 361632 612864 361638 612876
rect 363598 612864 363604 612876
rect 361632 612836 363604 612864
rect 361632 612824 361638 612836
rect 363598 612824 363604 612836
rect 363656 612824 363662 612876
rect 458634 603984 458640 604036
rect 458692 604024 458698 604036
rect 458910 604024 458916 604036
rect 458692 603996 458916 604024
rect 458692 603984 458698 603996
rect 458910 603984 458916 603996
rect 458968 603984 458974 604036
rect 459002 603712 459008 603764
rect 459060 603752 459066 603764
rect 459462 603752 459468 603764
rect 459060 603724 459468 603752
rect 459060 603712 459066 603724
rect 459462 603712 459468 603724
rect 459520 603712 459526 603764
rect 360838 602284 360844 602336
rect 360896 602324 360902 602336
rect 362954 602324 362960 602336
rect 360896 602296 362960 602324
rect 360896 602284 360902 602296
rect 362954 602284 362960 602296
rect 363012 602284 363018 602336
rect 459830 602080 459836 602132
rect 459888 602120 459894 602132
rect 460106 602120 460112 602132
rect 459888 602092 460112 602120
rect 459888 602080 459894 602092
rect 460106 602080 460112 602092
rect 460164 602080 460170 602132
rect 361758 601672 361764 601724
rect 361816 601712 361822 601724
rect 370498 601712 370504 601724
rect 361816 601684 370504 601712
rect 361816 601672 361822 601684
rect 370498 601672 370504 601684
rect 370556 601672 370562 601724
rect 460106 600244 460112 600296
rect 460164 600284 460170 600296
rect 462314 600284 462320 600296
rect 460164 600256 462320 600284
rect 460164 600244 460170 600256
rect 462314 600244 462320 600256
rect 462372 600244 462378 600296
rect 457806 600176 457812 600228
rect 457864 600216 457870 600228
rect 461578 600216 461584 600228
rect 457864 600188 461584 600216
rect 457864 600176 457870 600188
rect 461578 600176 461584 600188
rect 461636 600176 461642 600228
rect 458726 599768 458732 599820
rect 458784 599808 458790 599820
rect 465074 599808 465080 599820
rect 458784 599780 465080 599808
rect 458784 599768 458790 599780
rect 465074 599768 465080 599780
rect 465132 599768 465138 599820
rect 459002 599700 459008 599752
rect 459060 599740 459066 599752
rect 466454 599740 466460 599752
rect 459060 599712 466460 599740
rect 459060 599700 459066 599712
rect 466454 599700 466460 599712
rect 466512 599700 466518 599752
rect 457346 599632 457352 599684
rect 457404 599672 457410 599684
rect 467098 599672 467104 599684
rect 457404 599644 467104 599672
rect 457404 599632 457410 599644
rect 467098 599632 467104 599644
rect 467156 599632 467162 599684
rect 457254 599564 457260 599616
rect 457312 599604 457318 599616
rect 468478 599604 468484 599616
rect 457312 599576 468484 599604
rect 457312 599564 457318 599576
rect 468478 599564 468484 599576
rect 468536 599564 468542 599616
rect 457438 598748 457444 598800
rect 457496 598788 457502 598800
rect 461670 598788 461676 598800
rect 457496 598760 461676 598788
rect 457496 598748 457502 598760
rect 461670 598748 461676 598760
rect 461728 598748 461734 598800
rect 459462 598408 459468 598460
rect 459520 598448 459526 598460
rect 463694 598448 463700 598460
rect 459520 598420 463700 598448
rect 459520 598408 459526 598420
rect 463694 598408 463700 598420
rect 463752 598408 463758 598460
rect 362954 598340 362960 598392
rect 363012 598380 363018 598392
rect 365438 598380 365444 598392
rect 363012 598352 365444 598380
rect 363012 598340 363018 598352
rect 365438 598340 365444 598352
rect 365496 598340 365502 598392
rect 488626 598272 488632 598324
rect 488684 598312 488690 598324
rect 494330 598312 494336 598324
rect 488684 598284 494336 598312
rect 488684 598272 488690 598284
rect 494330 598272 494336 598284
rect 494388 598272 494394 598324
rect 460198 598204 460204 598256
rect 460256 598244 460262 598256
rect 467926 598244 467932 598256
rect 460256 598216 467932 598244
rect 460256 598204 460262 598216
rect 467926 598204 467932 598216
rect 467984 598204 467990 598256
rect 493318 598204 493324 598256
rect 493376 598244 493382 598256
rect 526714 598244 526720 598256
rect 493376 598216 526720 598244
rect 493376 598204 493382 598216
rect 526714 598204 526720 598216
rect 526772 598204 526778 598256
rect 457530 597524 457536 597576
rect 457588 597564 457594 597576
rect 462958 597564 462964 597576
rect 457588 597536 462964 597564
rect 457588 597524 457594 597536
rect 462958 597524 462964 597536
rect 463016 597524 463022 597576
rect 459830 596980 459836 597032
rect 459888 597020 459894 597032
rect 466546 597020 466552 597032
rect 459888 596992 466552 597020
rect 459888 596980 459894 596992
rect 466546 596980 466552 596992
rect 466604 596980 466610 597032
rect 457622 596912 457628 596964
rect 457680 596952 457686 596964
rect 464338 596952 464344 596964
rect 457680 596924 464344 596952
rect 457680 596912 457686 596924
rect 464338 596912 464344 596924
rect 464396 596912 464402 596964
rect 458634 596844 458640 596896
rect 458692 596884 458698 596896
rect 469398 596884 469404 596896
rect 458692 596856 469404 596884
rect 458692 596844 458698 596856
rect 469398 596844 469404 596856
rect 469456 596844 469462 596896
rect 450538 596776 450544 596828
rect 450596 596816 450602 596828
rect 494974 596816 494980 596828
rect 450596 596788 494980 596816
rect 450596 596776 450602 596788
rect 494974 596776 494980 596788
rect 495032 596776 495038 596828
rect 457714 595416 457720 595468
rect 457772 595456 457778 595468
rect 468570 595456 468576 595468
rect 457772 595428 468576 595456
rect 457772 595416 457778 595428
rect 468570 595416 468576 595428
rect 468628 595416 468634 595468
rect 459922 594056 459928 594108
rect 459980 594096 459986 594108
rect 463786 594096 463792 594108
rect 459980 594068 463792 594096
rect 459980 594056 459986 594068
rect 463786 594056 463792 594068
rect 463844 594056 463850 594108
rect 460014 592628 460020 592680
rect 460072 592668 460078 592680
rect 465166 592668 465172 592680
rect 460072 592640 465172 592668
rect 460072 592628 460078 592640
rect 465166 592628 465172 592640
rect 465224 592628 465230 592680
rect 361574 590792 361580 590844
rect 361632 590832 361638 590844
rect 363690 590832 363696 590844
rect 361632 590804 363696 590832
rect 361632 590792 361638 590804
rect 363690 590792 363696 590804
rect 363748 590792 363754 590844
rect 519538 590656 519544 590708
rect 519596 590696 519602 590708
rect 579614 590696 579620 590708
rect 519596 590668 579620 590696
rect 519596 590656 519602 590668
rect 579614 590656 579620 590668
rect 579672 590656 579678 590708
rect 365438 590588 365444 590640
rect 365496 590628 365502 590640
rect 367738 590628 367744 590640
rect 365496 590600 367744 590628
rect 365496 590588 365502 590600
rect 367738 590588 367744 590600
rect 367796 590588 367802 590640
rect 459186 587120 459192 587172
rect 459244 587160 459250 587172
rect 470594 587160 470600 587172
rect 459244 587132 470600 587160
rect 459244 587120 459250 587132
rect 470594 587120 470600 587132
rect 470652 587120 470658 587172
rect 459278 584400 459284 584452
rect 459336 584440 459342 584452
rect 470686 584440 470692 584452
rect 459336 584412 470692 584440
rect 459336 584400 459342 584412
rect 470686 584400 470692 584412
rect 470744 584400 470750 584452
rect 367738 582836 367744 582888
rect 367796 582876 367802 582888
rect 371234 582876 371240 582888
rect 367796 582848 371240 582876
rect 367796 582836 367802 582848
rect 371234 582836 371240 582848
rect 371292 582836 371298 582888
rect 361758 579640 361764 579692
rect 361816 579680 361822 579692
rect 367738 579680 367744 579692
rect 361816 579652 367744 579680
rect 361816 579640 361822 579652
rect 367738 579640 367744 579652
rect 367796 579640 367802 579692
rect 371234 578892 371240 578944
rect 371292 578932 371298 578944
rect 373994 578932 374000 578944
rect 371292 578904 374000 578932
rect 371292 578892 371298 578904
rect 373994 578892 374000 578904
rect 374052 578892 374058 578944
rect 511258 576852 511264 576904
rect 511316 576892 511322 576904
rect 579614 576892 579620 576904
rect 511316 576864 579620 576892
rect 511316 576852 511322 576864
rect 579614 576852 579620 576864
rect 579672 576852 579678 576904
rect 373994 575492 374000 575544
rect 374052 575532 374058 575544
rect 374052 575504 376800 575532
rect 374052 575492 374058 575504
rect 376772 575464 376800 575504
rect 378134 575464 378140 575476
rect 376772 575436 378140 575464
rect 378134 575424 378140 575436
rect 378192 575424 378198 575476
rect 378134 569848 378140 569900
rect 378192 569888 378198 569900
rect 380342 569888 380348 569900
rect 378192 569860 380348 569888
rect 378192 569848 378198 569860
rect 380342 569848 380348 569860
rect 380400 569848 380406 569900
rect 361574 568760 361580 568812
rect 361632 568800 361638 568812
rect 363782 568800 363788 568812
rect 361632 568772 363788 568800
rect 361632 568760 361638 568772
rect 363782 568760 363788 568772
rect 363840 568760 363846 568812
rect 515398 563048 515404 563100
rect 515456 563088 515462 563100
rect 579890 563088 579896 563100
rect 515456 563060 579896 563088
rect 515456 563048 515462 563060
rect 579890 563048 579896 563060
rect 579948 563048 579954 563100
rect 380342 562980 380348 563032
rect 380400 563020 380406 563032
rect 382274 563020 382280 563032
rect 380400 562992 382280 563020
rect 380400 562980 380406 562992
rect 382274 562980 382280 562992
rect 382332 562980 382338 563032
rect 382274 559716 382280 559768
rect 382332 559756 382338 559768
rect 385034 559756 385040 559768
rect 382332 559728 385040 559756
rect 382332 559716 382338 559728
rect 385034 559716 385040 559728
rect 385092 559716 385098 559768
rect 361666 557540 361672 557592
rect 361724 557580 361730 557592
rect 403618 557580 403624 557592
rect 361724 557552 403624 557580
rect 361724 557540 361730 557552
rect 403618 557540 403624 557552
rect 403676 557540 403682 557592
rect 385034 555568 385040 555620
rect 385092 555608 385098 555620
rect 387058 555608 387064 555620
rect 385092 555580 387064 555608
rect 385092 555568 385098 555580
rect 387058 555568 387064 555580
rect 387116 555568 387122 555620
rect 387058 553392 387064 553444
rect 387116 553432 387122 553444
rect 387116 553404 387840 553432
rect 387116 553392 387122 553404
rect 387812 553364 387840 553404
rect 389818 553364 389824 553376
rect 387812 553336 389824 553364
rect 389818 553324 389824 553336
rect 389876 553324 389882 553376
rect 457898 551284 457904 551336
rect 457956 551324 457962 551336
rect 467190 551324 467196 551336
rect 457956 551296 467196 551324
rect 457956 551284 457962 551296
rect 467190 551284 467196 551296
rect 467248 551284 467254 551336
rect 361758 546456 361764 546508
rect 361816 546496 361822 546508
rect 419074 546496 419080 546508
rect 361816 546468 419080 546496
rect 361816 546456 361822 546468
rect 419074 546456 419080 546468
rect 419132 546456 419138 546508
rect 389818 540948 389824 541000
rect 389876 540988 389882 541000
rect 389876 540960 390600 540988
rect 389876 540948 389882 540960
rect 390572 540920 390600 540960
rect 392302 540920 392308 540932
rect 390572 540892 392308 540920
rect 392302 540880 392308 540892
rect 392360 540880 392366 540932
rect 392302 536800 392308 536852
rect 392360 536840 392366 536852
rect 392360 536812 393314 536840
rect 392360 536800 392366 536812
rect 393286 536772 393314 536812
rect 394694 536772 394700 536784
rect 393286 536744 394700 536772
rect 394694 536732 394700 536744
rect 394752 536732 394758 536784
rect 361758 535440 361764 535492
rect 361816 535480 361822 535492
rect 406378 535480 406384 535492
rect 361816 535452 406384 535480
rect 361816 535440 361822 535452
rect 406378 535440 406384 535452
rect 406436 535440 406442 535492
rect 394694 529864 394700 529916
rect 394752 529904 394758 529916
rect 396718 529904 396724 529916
rect 394752 529876 396724 529904
rect 394752 529864 394758 529876
rect 396718 529864 396724 529876
rect 396776 529864 396782 529916
rect 361758 524424 361764 524476
rect 361816 524464 361822 524476
rect 407758 524464 407764 524476
rect 361816 524436 407764 524464
rect 361816 524424 361822 524436
rect 407758 524424 407764 524436
rect 407816 524424 407822 524476
rect 457990 523676 457996 523728
rect 458048 523716 458054 523728
rect 465718 523716 465724 523728
rect 458048 523688 465724 523716
rect 458048 523676 458054 523688
rect 465718 523676 465724 523688
rect 465776 523676 465782 523728
rect 482922 520888 482928 520940
rect 482980 520928 482986 520940
rect 520274 520928 520280 520940
rect 482980 520900 520280 520928
rect 482980 520888 482986 520900
rect 520274 520888 520280 520900
rect 520332 520888 520338 520940
rect 461762 520276 461768 520328
rect 461820 520316 461826 520328
rect 488626 520316 488632 520328
rect 461820 520288 488632 520316
rect 461820 520276 461826 520288
rect 488626 520276 488632 520288
rect 488684 520276 488690 520328
rect 459370 519528 459376 519580
rect 459428 519568 459434 519580
rect 469306 519568 469312 519580
rect 459428 519540 469312 519568
rect 459428 519528 459434 519540
rect 469306 519528 469312 519540
rect 469364 519528 469370 519580
rect 458082 518236 458088 518288
rect 458140 518276 458146 518288
rect 464430 518276 464436 518288
rect 458140 518248 464436 518276
rect 458140 518236 458146 518248
rect 464430 518236 464436 518248
rect 464488 518236 464494 518288
rect 449802 518168 449808 518220
rect 449860 518208 449866 518220
rect 469858 518208 469864 518220
rect 449860 518180 469864 518208
rect 449860 518168 449866 518180
rect 469858 518168 469864 518180
rect 469916 518208 469922 518220
rect 494238 518208 494244 518220
rect 469916 518180 494244 518208
rect 469916 518168 469922 518180
rect 494238 518168 494244 518180
rect 494296 518168 494302 518220
rect 476022 517556 476028 517608
rect 476080 517596 476086 517608
rect 494146 517596 494152 517608
rect 476080 517568 494152 517596
rect 476080 517556 476086 517568
rect 494146 517556 494152 517568
rect 494204 517556 494210 517608
rect 450354 517488 450360 517540
rect 450412 517528 450418 517540
rect 494330 517528 494336 517540
rect 450412 517500 494336 517528
rect 450412 517488 450418 517500
rect 494330 517488 494336 517500
rect 494388 517488 494394 517540
rect 482278 517420 482284 517472
rect 482336 517420 482342 517472
rect 450630 516808 450636 516860
rect 450688 516848 450694 516860
rect 476022 516848 476028 516860
rect 450688 516820 476028 516848
rect 450688 516808 450694 516820
rect 476022 516808 476028 516820
rect 476080 516808 476086 516860
rect 449986 516740 449992 516792
rect 450044 516780 450050 516792
rect 482296 516780 482324 517420
rect 492122 516780 492128 516792
rect 450044 516752 492128 516780
rect 450044 516740 450050 516752
rect 492122 516740 492128 516752
rect 492180 516740 492186 516792
rect 3970 514768 3976 514820
rect 4028 514808 4034 514820
rect 4798 514808 4804 514820
rect 4028 514780 4804 514808
rect 4028 514768 4034 514780
rect 4798 514768 4804 514780
rect 4856 514768 4862 514820
rect 502242 514020 502248 514072
rect 502300 514060 502306 514072
rect 545114 514060 545120 514072
rect 502300 514032 545120 514060
rect 502300 514020 502306 514032
rect 545114 514020 545120 514032
rect 545172 514020 545178 514072
rect 361758 513340 361764 513392
rect 361816 513380 361822 513392
rect 410518 513380 410524 513392
rect 361816 513352 410524 513380
rect 361816 513340 361822 513352
rect 410518 513340 410524 513352
rect 410576 513340 410582 513392
rect 492122 512592 492128 512644
rect 492180 512632 492186 512644
rect 535454 512632 535460 512644
rect 492180 512604 535460 512632
rect 492180 512592 492186 512604
rect 535454 512592 535460 512604
rect 535512 512592 535518 512644
rect 396718 511912 396724 511964
rect 396776 511952 396782 511964
rect 400950 511952 400956 511964
rect 396776 511924 400956 511952
rect 396776 511912 396782 511924
rect 400950 511912 400956 511924
rect 401008 511912 401014 511964
rect 519630 510620 519636 510672
rect 519688 510660 519694 510672
rect 579614 510660 579620 510672
rect 519688 510632 579620 510660
rect 519688 510620 519694 510632
rect 579614 510620 579620 510632
rect 579672 510620 579678 510672
rect 494330 509872 494336 509924
rect 494388 509912 494394 509924
rect 538214 509912 538220 509924
rect 494388 509884 538220 509912
rect 494388 509872 494394 509884
rect 538214 509872 538220 509884
rect 538272 509872 538278 509924
rect 494146 508512 494152 508564
rect 494204 508552 494210 508564
rect 532694 508552 532700 508564
rect 494204 508524 532700 508552
rect 494204 508512 494210 508524
rect 532694 508512 532700 508524
rect 532752 508512 532758 508564
rect 495066 505724 495072 505776
rect 495124 505764 495130 505776
rect 529934 505764 529940 505776
rect 495124 505736 529940 505764
rect 495124 505724 495130 505736
rect 529934 505724 529940 505736
rect 529992 505724 529998 505776
rect 361758 502324 361764 502376
rect 361816 502364 361822 502376
rect 411898 502364 411904 502376
rect 361816 502336 411904 502364
rect 361816 502324 361822 502336
rect 411898 502324 411904 502336
rect 411956 502324 411962 502376
rect 461854 497700 461860 497752
rect 461912 497740 461918 497752
rect 482646 497740 482652 497752
rect 461912 497712 482652 497740
rect 461912 497700 461918 497712
rect 482646 497700 482652 497712
rect 482704 497700 482710 497752
rect 457622 497632 457628 497684
rect 457680 497672 457686 497684
rect 480254 497672 480260 497684
rect 457680 497644 480260 497672
rect 457680 497632 457686 497644
rect 480254 497632 480260 497644
rect 480312 497632 480318 497684
rect 457438 497564 457444 497616
rect 457496 497604 457502 497616
rect 483842 497604 483848 497616
rect 457496 497576 483848 497604
rect 457496 497564 457502 497576
rect 483842 497564 483848 497576
rect 483900 497564 483906 497616
rect 458818 497496 458824 497548
rect 458876 497536 458882 497548
rect 485038 497536 485044 497548
rect 458876 497508 485044 497536
rect 458876 497496 458882 497508
rect 485038 497496 485044 497508
rect 485096 497496 485102 497548
rect 453298 497428 453304 497480
rect 453356 497468 453362 497480
rect 481634 497468 481640 497480
rect 453356 497440 481640 497468
rect 453356 497428 453362 497440
rect 481634 497428 481640 497440
rect 481692 497428 481698 497480
rect 455322 497020 455328 497072
rect 455380 497060 455386 497072
rect 459554 497060 459560 497072
rect 455380 497032 459560 497060
rect 455380 497020 455386 497032
rect 459554 497020 459560 497032
rect 459612 497020 459618 497072
rect 456518 496952 456524 497004
rect 456576 496992 456582 497004
rect 461026 496992 461032 497004
rect 456576 496964 461032 496992
rect 456576 496952 456582 496964
rect 461026 496952 461032 496964
rect 461084 496952 461090 497004
rect 455138 496884 455144 496936
rect 455196 496924 455202 496936
rect 458082 496924 458088 496936
rect 455196 496896 458088 496924
rect 455196 496884 455202 496896
rect 458082 496884 458088 496896
rect 458140 496884 458146 496936
rect 452562 496816 452568 496868
rect 452620 496856 452626 496868
rect 453666 496856 453672 496868
rect 452620 496828 453672 496856
rect 452620 496816 452626 496828
rect 453666 496816 453672 496828
rect 453724 496816 453730 496868
rect 453942 496816 453948 496868
rect 454000 496856 454006 496868
rect 456610 496856 456616 496868
rect 454000 496828 456616 496856
rect 454000 496816 454006 496828
rect 456610 496816 456616 496828
rect 456668 496816 456674 496868
rect 400950 495456 400956 495508
rect 401008 495496 401014 495508
rect 402238 495496 402244 495508
rect 401008 495468 402244 495496
rect 401008 495456 401014 495468
rect 402238 495456 402244 495468
rect 402296 495456 402302 495508
rect 361758 491308 361764 491360
rect 361816 491348 361822 491360
rect 381538 491348 381544 491360
rect 361816 491320 381544 491348
rect 361816 491308 361822 491320
rect 381538 491308 381544 491320
rect 381596 491308 381602 491360
rect 518158 484372 518164 484424
rect 518216 484412 518222 484424
rect 580166 484412 580172 484424
rect 518216 484384 580172 484412
rect 518216 484372 518222 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 361758 480224 361764 480276
rect 361816 480264 361822 480276
rect 419166 480264 419172 480276
rect 361816 480236 419172 480264
rect 361816 480224 361822 480236
rect 419166 480224 419172 480236
rect 419224 480224 419230 480276
rect 515490 470568 515496 470620
rect 515548 470608 515554 470620
rect 579982 470608 579988 470620
rect 515548 470580 579988 470608
rect 515548 470568 515554 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 361758 469208 361764 469260
rect 361816 469248 361822 469260
rect 396718 469248 396724 469260
rect 361816 469220 396724 469248
rect 361816 469208 361822 469220
rect 396718 469208 396724 469220
rect 396776 469208 396782 469260
rect 494698 462408 494704 462460
rect 494756 462448 494762 462460
rect 527634 462448 527640 462460
rect 494756 462420 527640 462448
rect 494756 462408 494762 462420
rect 527634 462408 527640 462420
rect 527692 462408 527698 462460
rect 402238 462340 402244 462392
rect 402296 462380 402302 462392
rect 404998 462380 405004 462392
rect 402296 462352 405004 462380
rect 402296 462340 402302 462352
rect 404998 462340 405004 462352
rect 405056 462340 405062 462392
rect 450538 462340 450544 462392
rect 450596 462380 450602 462392
rect 542354 462380 542360 462392
rect 450596 462352 542360 462380
rect 450596 462340 450602 462352
rect 542354 462340 542360 462352
rect 542412 462340 542418 462392
rect 448974 461048 448980 461100
rect 449032 461088 449038 461100
rect 524690 461088 524696 461100
rect 449032 461060 524696 461088
rect 449032 461048 449038 461060
rect 524690 461048 524696 461060
rect 524748 461048 524754 461100
rect 468662 460980 468668 461032
rect 468720 461020 468726 461032
rect 553854 461020 553860 461032
rect 468720 460992 553860 461020
rect 468720 460980 468726 460992
rect 553854 460980 553860 460992
rect 553912 460980 553918 461032
rect 458910 460912 458916 460964
rect 458968 460952 458974 460964
rect 550910 460952 550916 460964
rect 458968 460924 550916 460952
rect 458968 460912 458974 460924
rect 550910 460912 550916 460924
rect 550968 460912 550974 460964
rect 361758 458192 361764 458244
rect 361816 458232 361822 458244
rect 414658 458232 414664 458244
rect 361816 458204 414664 458232
rect 361816 458192 361822 458204
rect 414658 458192 414664 458204
rect 414716 458192 414722 458244
rect 449618 457444 449624 457496
rect 449676 457484 449682 457496
rect 489914 457484 489920 457496
rect 449676 457456 489920 457484
rect 449676 457444 449682 457456
rect 489914 457444 489920 457456
rect 489972 457444 489978 457496
rect 569218 456764 569224 456816
rect 569276 456804 569282 456816
rect 580166 456804 580172 456816
rect 569276 456776 580172 456804
rect 569276 456764 569282 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 488258 456016 488264 456068
rect 488316 456056 488322 456068
rect 494698 456056 494704 456068
rect 488316 456028 494704 456056
rect 488316 456016 488322 456028
rect 494698 456016 494704 456028
rect 494756 456016 494762 456068
rect 452010 455472 452016 455524
rect 452068 455512 452074 455524
rect 480990 455512 480996 455524
rect 452068 455484 480996 455512
rect 452068 455472 452074 455484
rect 480990 455472 480996 455484
rect 481048 455472 481054 455524
rect 454678 455404 454684 455456
rect 454736 455444 454742 455456
rect 488258 455444 488264 455456
rect 454736 455416 488264 455444
rect 454736 455404 454742 455416
rect 488258 455404 488264 455416
rect 488316 455404 488322 455456
rect 449710 454724 449716 454776
rect 449768 454764 449774 454776
rect 485774 454764 485780 454776
rect 449768 454736 485780 454764
rect 449768 454724 449774 454736
rect 485774 454724 485780 454736
rect 485832 454724 485838 454776
rect 449526 454656 449532 454708
rect 449584 454696 449590 454708
rect 487154 454696 487160 454708
rect 449584 454668 487160 454696
rect 449584 454656 449590 454668
rect 487154 454656 487160 454668
rect 487212 454656 487218 454708
rect 459002 454044 459008 454096
rect 459060 454084 459066 454096
rect 473722 454084 473728 454096
rect 459060 454056 473728 454084
rect 459060 454044 459066 454056
rect 473722 454044 473728 454056
rect 473780 454044 473786 454096
rect 404998 453976 405004 454028
rect 405056 454016 405062 454028
rect 408402 454016 408408 454028
rect 405056 453988 408408 454016
rect 405056 453976 405062 453988
rect 408402 453976 408408 453988
rect 408460 453976 408466 454028
rect 408402 448536 408408 448588
rect 408460 448576 408466 448588
rect 408460 448548 408540 448576
rect 408460 448536 408466 448548
rect 408512 448508 408540 448548
rect 410426 448508 410432 448520
rect 408512 448480 410432 448508
rect 410426 448468 410432 448480
rect 410484 448468 410490 448520
rect 447318 447924 447324 447976
rect 447376 447964 447382 447976
rect 448422 447964 448428 447976
rect 447376 447936 448428 447964
rect 447376 447924 447382 447936
rect 448422 447924 448428 447936
rect 448480 447964 448486 447976
rect 459002 447964 459008 447976
rect 448480 447936 459008 447964
rect 448480 447924 448486 447936
rect 459002 447924 459008 447936
rect 459060 447924 459066 447976
rect 447226 447856 447232 447908
rect 447284 447896 447290 447908
rect 448054 447896 448060 447908
rect 447284 447868 448060 447896
rect 447284 447856 447290 447868
rect 448054 447856 448060 447868
rect 448112 447896 448118 447908
rect 458910 447896 458916 447908
rect 448112 447868 458916 447896
rect 448112 447856 448118 447868
rect 458910 447856 458916 447868
rect 458968 447856 458974 447908
rect 447134 447788 447140 447840
rect 447192 447828 447198 447840
rect 447686 447828 447692 447840
rect 447192 447800 447692 447828
rect 447192 447788 447198 447800
rect 447686 447788 447692 447800
rect 447744 447828 447750 447840
rect 468662 447828 468668 447840
rect 447744 447800 468668 447828
rect 447744 447788 447750 447800
rect 468662 447788 468668 447800
rect 468720 447788 468726 447840
rect 422478 447380 422484 447432
rect 422536 447420 422542 447432
rect 447318 447420 447324 447432
rect 422536 447392 447324 447420
rect 422536 447380 422542 447392
rect 447318 447380 447324 447392
rect 447376 447380 447382 447432
rect 437382 447312 437388 447364
rect 437440 447352 437446 447364
rect 447134 447352 447140 447364
rect 437440 447324 447140 447352
rect 437440 447312 437446 447324
rect 447134 447312 447140 447324
rect 447192 447312 447198 447364
rect 432414 447244 432420 447296
rect 432472 447284 432478 447296
rect 447226 447284 447232 447296
rect 432472 447256 447232 447284
rect 432472 447244 432478 447256
rect 447226 447244 447232 447256
rect 447284 447244 447290 447296
rect 427446 447176 427452 447228
rect 427504 447216 427510 447228
rect 445662 447216 445668 447228
rect 427504 447188 445668 447216
rect 427504 447176 427510 447188
rect 445662 447176 445668 447188
rect 445720 447176 445726 447228
rect 361758 447108 361764 447160
rect 361816 447148 361822 447160
rect 399478 447148 399484 447160
rect 361816 447120 399484 447148
rect 361816 447108 361822 447120
rect 399478 447108 399484 447120
rect 399536 447108 399542 447160
rect 410426 445680 410432 445732
rect 410484 445720 410490 445732
rect 413278 445720 413284 445732
rect 410484 445692 413284 445720
rect 410484 445680 410490 445692
rect 413278 445680 413284 445692
rect 413336 445680 413342 445732
rect 429838 445000 429844 445052
rect 429896 445040 429902 445052
rect 447134 445040 447140 445052
rect 429896 445012 447140 445040
rect 429896 445000 429902 445012
rect 447134 445000 447140 445012
rect 447192 445000 447198 445052
rect 442626 444320 442632 444372
rect 442684 444360 442690 444372
rect 446214 444360 446220 444372
rect 442684 444332 446220 444360
rect 442684 444320 442690 444332
rect 446214 444320 446220 444332
rect 446272 444320 446278 444372
rect 361758 436092 361764 436144
rect 361816 436132 361822 436144
rect 416130 436132 416136 436144
rect 361816 436104 416136 436132
rect 361816 436092 361822 436104
rect 416130 436092 416136 436104
rect 416188 436092 416194 436144
rect 413278 433236 413284 433288
rect 413336 433276 413342 433288
rect 414750 433276 414756 433288
rect 413336 433248 414756 433276
rect 413336 433236 413342 433248
rect 414750 433236 414756 433248
rect 414808 433236 414814 433288
rect 573358 430584 573364 430636
rect 573416 430624 573422 430636
rect 579614 430624 579620 430636
rect 573416 430596 579620 430624
rect 573416 430584 573422 430596
rect 579614 430584 579620 430596
rect 579672 430584 579678 430636
rect 458082 429972 458088 430024
rect 458140 430012 458146 430024
rect 474274 430012 474280 430024
rect 458140 429984 474280 430012
rect 458140 429972 458146 429984
rect 474274 429972 474280 429984
rect 474332 429972 474338 430024
rect 459370 429904 459376 429956
rect 459428 429944 459434 429956
rect 476942 429944 476948 429956
rect 459428 429916 476948 429944
rect 459428 429904 459434 429916
rect 476942 429904 476948 429916
rect 477000 429904 477006 429956
rect 459462 429836 459468 429888
rect 459520 429876 459526 429888
rect 479610 429876 479616 429888
rect 459520 429848 479616 429876
rect 459520 429836 459526 429848
rect 479610 429836 479616 429848
rect 479668 429836 479674 429888
rect 480898 429156 480904 429208
rect 480956 429196 480962 429208
rect 482278 429196 482284 429208
rect 480956 429168 482284 429196
rect 480956 429156 480962 429168
rect 482278 429156 482284 429168
rect 482336 429156 482342 429208
rect 483658 429156 483664 429208
rect 483716 429196 483722 429208
rect 484946 429196 484952 429208
rect 483716 429168 484952 429196
rect 483716 429156 483722 429168
rect 484946 429156 484952 429168
rect 485004 429156 485010 429208
rect 457530 428408 457536 428460
rect 457588 428448 457594 428460
rect 471606 428448 471612 428460
rect 457588 428420 471612 428448
rect 457588 428408 457594 428420
rect 471606 428408 471612 428420
rect 471664 428408 471670 428460
rect 361758 425076 361764 425128
rect 361816 425116 361822 425128
rect 417418 425116 417424 425128
rect 361816 425088 417424 425116
rect 361816 425076 361822 425088
rect 417418 425076 417424 425088
rect 417476 425076 417482 425128
rect 529198 423580 529204 423632
rect 529256 423620 529262 423632
rect 530210 423620 530216 423632
rect 529256 423592 530216 423620
rect 529256 423580 529262 423592
rect 530210 423580 530216 423592
rect 530268 423580 530274 423632
rect 530578 423580 530584 423632
rect 530636 423620 530642 423632
rect 532786 423620 532792 423632
rect 530636 423592 532792 423620
rect 530636 423580 530642 423592
rect 532786 423580 532792 423592
rect 532844 423580 532850 423632
rect 511350 423512 511356 423564
rect 511408 423552 511414 423564
rect 523770 423552 523776 423564
rect 511408 423524 523776 423552
rect 511408 423512 511414 423524
rect 523770 423512 523776 423524
rect 523828 423512 523834 423564
rect 522298 423444 522304 423496
rect 522356 423484 522362 423496
rect 549530 423484 549536 423496
rect 522356 423456 549536 423484
rect 522356 423444 522362 423456
rect 549530 423444 549536 423456
rect 549588 423444 549594 423496
rect 502978 423376 502984 423428
rect 503036 423416 503042 423428
rect 522482 423416 522488 423428
rect 503036 423388 522488 423416
rect 503036 423376 503042 423388
rect 522482 423376 522488 423388
rect 522540 423376 522546 423428
rect 523678 423376 523684 423428
rect 523736 423416 523742 423428
rect 552106 423416 552112 423428
rect 523736 423388 552112 423416
rect 523736 423376 523742 423388
rect 552106 423376 552112 423388
rect 552164 423376 552170 423428
rect 487062 423308 487068 423360
rect 487120 423348 487126 423360
rect 526346 423348 526352 423360
rect 487120 423320 526352 423348
rect 487120 423308 487126 423320
rect 526346 423308 526352 423320
rect 526404 423308 526410 423360
rect 526438 423308 526444 423360
rect 526496 423348 526502 423360
rect 554682 423348 554688 423360
rect 526496 423320 554688 423348
rect 526496 423308 526502 423320
rect 554682 423308 554688 423320
rect 554740 423308 554746 423360
rect 488258 423240 488264 423292
rect 488316 423280 488322 423292
rect 528922 423280 528928 423292
rect 488316 423252 528928 423280
rect 488316 423240 488322 423252
rect 528922 423240 528928 423252
rect 528980 423240 528986 423292
rect 489638 423172 489644 423224
rect 489696 423212 489702 423224
rect 531498 423212 531504 423224
rect 489696 423184 531504 423212
rect 489696 423172 489702 423184
rect 531498 423172 531504 423184
rect 531556 423172 531562 423224
rect 498102 423104 498108 423156
rect 498160 423144 498166 423156
rect 545666 423144 545672 423156
rect 498160 423116 545672 423144
rect 498160 423104 498166 423116
rect 545666 423104 545672 423116
rect 545724 423104 545730 423156
rect 499298 423036 499304 423088
rect 499356 423076 499362 423088
rect 548242 423076 548248 423088
rect 499356 423048 548248 423076
rect 499356 423036 499362 423048
rect 548242 423036 548248 423048
rect 548300 423036 548306 423088
rect 500678 422968 500684 423020
rect 500736 423008 500742 423020
rect 550818 423008 550824 423020
rect 500736 422980 550824 423008
rect 500736 422968 500742 422980
rect 550818 422968 550824 422980
rect 550876 422968 550882 423020
rect 444282 422900 444288 422952
rect 444340 422940 444346 422952
rect 447962 422940 447968 422952
rect 444340 422912 447968 422940
rect 444340 422900 444346 422912
rect 447962 422900 447968 422912
rect 448020 422900 448026 422952
rect 502242 422900 502248 422952
rect 502300 422940 502306 422952
rect 553394 422940 553400 422952
rect 502300 422912 553400 422940
rect 502300 422900 502306 422912
rect 553394 422900 553400 422912
rect 553452 422900 553458 422952
rect 484302 421540 484308 421592
rect 484360 421580 484366 421592
rect 521194 421580 521200 421592
rect 484360 421552 521200 421580
rect 484360 421540 484366 421552
rect 521194 421540 521200 421552
rect 521252 421540 521258 421592
rect 414750 420928 414756 420980
rect 414808 420968 414814 420980
rect 414808 420940 418200 420968
rect 414808 420928 414814 420940
rect 418172 420900 418200 420940
rect 420914 420900 420920 420912
rect 418172 420872 420920 420900
rect 420914 420860 420920 420872
rect 420972 420860 420978 420912
rect 495342 420180 495348 420232
rect 495400 420220 495406 420232
rect 541802 420220 541808 420232
rect 495400 420192 541808 420220
rect 495400 420180 495406 420192
rect 541802 420180 541808 420192
rect 541860 420180 541866 420232
rect 442810 419500 442816 419552
rect 442868 419540 442874 419552
rect 447870 419540 447876 419552
rect 442868 419512 447876 419540
rect 442868 419500 442874 419512
rect 447870 419500 447876 419512
rect 447928 419500 447934 419552
rect 424686 417732 424692 417784
rect 424744 417772 424750 417784
rect 506474 417772 506480 417784
rect 424744 417744 506480 417772
rect 424744 417732 424750 417744
rect 506474 417732 506480 417744
rect 506532 417732 506538 417784
rect 421466 417664 421472 417716
rect 421524 417704 421530 417716
rect 503714 417704 503720 417716
rect 421524 417676 503720 417704
rect 421524 417664 421530 417676
rect 503714 417664 503720 417676
rect 503772 417664 503778 417716
rect 425974 417596 425980 417648
rect 426032 417636 426038 417648
rect 507854 417636 507860 417648
rect 426032 417608 507860 417636
rect 426032 417596 426038 417608
rect 507854 417596 507860 417608
rect 507912 417596 507918 417648
rect 420914 417528 420920 417580
rect 420972 417568 420978 417580
rect 425054 417568 425060 417580
rect 420972 417540 425060 417568
rect 420972 417528 420978 417540
rect 425054 417528 425060 417540
rect 425112 417528 425118 417580
rect 425330 417528 425336 417580
rect 425388 417568 425394 417580
rect 507946 417568 507952 417580
rect 425388 417540 507952 417568
rect 425388 417528 425394 417540
rect 507946 417528 507952 417540
rect 508004 417528 508010 417580
rect 422110 417460 422116 417512
rect 422168 417500 422174 417512
rect 503990 417500 503996 417512
rect 422168 417472 503996 417500
rect 422168 417460 422174 417472
rect 503990 417460 503996 417472
rect 504048 417460 504054 417512
rect 424042 417392 424048 417444
rect 424100 417432 424106 417444
rect 506566 417432 506572 417444
rect 424100 417404 506572 417432
rect 424100 417392 424106 417404
rect 506566 417392 506572 417404
rect 506624 417392 506630 417444
rect 423122 416304 423128 416356
rect 423180 416344 423186 416356
rect 423582 416344 423588 416356
rect 423180 416316 423588 416344
rect 423180 416304 423186 416316
rect 423582 416304 423588 416316
rect 423640 416304 423646 416356
rect 486970 416032 486976 416084
rect 487028 416072 487034 416084
rect 527634 416072 527640 416084
rect 487028 416044 527640 416072
rect 487028 416032 487034 416044
rect 527634 416032 527640 416044
rect 527692 416032 527698 416084
rect 361574 413992 361580 414044
rect 361632 414032 361638 414044
rect 443638 414032 443644 414044
rect 361632 414004 443644 414032
rect 361632 413992 361638 414004
rect 443638 413992 443644 414004
rect 443696 413992 443702 414044
rect 425054 413924 425060 413976
rect 425112 413964 425118 413976
rect 427078 413964 427084 413976
rect 425112 413936 427084 413964
rect 425112 413924 425118 413936
rect 427078 413924 427084 413936
rect 427136 413924 427142 413976
rect 361574 402976 361580 403028
rect 361632 403016 361638 403028
rect 439498 403016 439504 403028
rect 361632 402988 439504 403016
rect 361632 402976 361638 402988
rect 439498 402976 439504 402988
rect 439556 402976 439562 403028
rect 503438 402228 503444 402280
rect 503496 402268 503502 402280
rect 557534 402268 557540 402280
rect 503496 402240 557540 402268
rect 503496 402228 503502 402240
rect 557534 402228 557540 402240
rect 557592 402228 557598 402280
rect 497918 400868 497924 400920
rect 497976 400908 497982 400920
rect 546494 400908 546500 400920
rect 497976 400880 546500 400908
rect 497976 400868 497982 400880
rect 546494 400868 546500 400880
rect 546552 400868 546558 400920
rect 494606 399440 494612 399492
rect 494664 399480 494670 399492
rect 539594 399480 539600 399492
rect 494664 399452 539600 399480
rect 494664 399440 494670 399452
rect 539594 399440 539600 399452
rect 539652 399440 539658 399492
rect 493962 398080 493968 398132
rect 494020 398120 494026 398132
rect 538214 398120 538220 398132
rect 494020 398092 538220 398120
rect 494020 398080 494026 398092
rect 538214 398080 538220 398092
rect 538272 398080 538278 398132
rect 427078 397400 427084 397452
rect 427136 397440 427142 397452
rect 428458 397440 428464 397452
rect 427136 397412 428464 397440
rect 427136 397400 427142 397412
rect 428458 397400 428464 397412
rect 428516 397400 428522 397452
rect 493134 396720 493140 396772
rect 493192 396760 493198 396772
rect 536834 396760 536840 396772
rect 493192 396732 536840 396760
rect 493192 396720 493198 396732
rect 536834 396720 536840 396732
rect 536892 396720 536898 396772
rect 460750 395292 460756 395344
rect 460808 395332 460814 395344
rect 483658 395332 483664 395344
rect 460808 395304 483664 395332
rect 460808 395292 460814 395304
rect 483658 395292 483664 395304
rect 483716 395292 483722 395344
rect 492398 395292 492404 395344
rect 492456 395332 492462 395344
rect 535454 395332 535460 395344
rect 492456 395304 535460 395332
rect 492456 395292 492462 395304
rect 535454 395292 535460 395304
rect 535512 395292 535518 395344
rect 496722 394000 496728 394052
rect 496780 394040 496786 394052
rect 543734 394040 543740 394052
rect 496780 394012 543740 394040
rect 496780 394000 496786 394012
rect 543734 394000 543740 394012
rect 543792 394000 543798 394052
rect 423490 393932 423496 393984
rect 423548 393972 423554 393984
rect 505554 393972 505560 393984
rect 423548 393944 505560 393972
rect 423548 393932 423554 393944
rect 505554 393932 505560 393944
rect 505612 393932 505618 393984
rect 463602 392572 463608 392624
rect 463660 392612 463666 392624
rect 487154 392612 487160 392624
rect 463660 392584 487160 392612
rect 463660 392572 463666 392584
rect 487154 392572 487160 392584
rect 487212 392572 487218 392624
rect 491570 392572 491576 392624
rect 491628 392612 491634 392624
rect 534166 392612 534172 392624
rect 491628 392584 534172 392612
rect 491628 392572 491634 392584
rect 534166 392572 534172 392584
rect 534224 392572 534230 392624
rect 361574 391960 361580 392012
rect 361632 392000 361638 392012
rect 443730 392000 443736 392012
rect 361632 391972 443736 392000
rect 361632 391960 361638 391972
rect 443730 391960 443736 391972
rect 443788 391960 443794 392012
rect 495710 391280 495716 391332
rect 495768 391320 495774 391332
rect 542354 391320 542360 391332
rect 495768 391292 542360 391320
rect 495768 391280 495774 391292
rect 542354 391280 542360 391292
rect 542412 391280 542418 391332
rect 423582 391212 423588 391264
rect 423640 391252 423646 391264
rect 505278 391252 505284 391264
rect 423640 391224 505284 391252
rect 423640 391212 423646 391224
rect 505278 391212 505284 391224
rect 505336 391212 505342 391264
rect 459646 389852 459652 389904
rect 459704 389892 459710 389904
rect 480898 389892 480904 389904
rect 459704 389864 480904 389892
rect 459704 389852 459710 389864
rect 480898 389852 480904 389864
rect 480956 389852 480962 389904
rect 464890 389784 464896 389836
rect 464948 389824 464954 389836
rect 489914 389824 489920 389836
rect 464948 389796 489920 389824
rect 464948 389784 464954 389796
rect 489914 389784 489920 389796
rect 489972 389784 489978 389836
rect 490558 389784 490564 389836
rect 490616 389824 490622 389836
rect 534074 389824 534080 389836
rect 490616 389796 534080 389824
rect 490616 389784 490622 389796
rect 534074 389784 534080 389796
rect 534132 389784 534138 389836
rect 465074 389240 465080 389292
rect 465132 389280 465138 389292
rect 465902 389280 465908 389292
rect 465132 389252 465908 389280
rect 465132 389240 465138 389252
rect 465902 389240 465908 389252
rect 465960 389240 465966 389292
rect 466454 389240 466460 389292
rect 466512 389280 466518 389292
rect 467374 389280 467380 389292
rect 466512 389252 467380 389280
rect 466512 389240 466518 389252
rect 467374 389240 467380 389252
rect 467432 389240 467438 389292
rect 470594 389240 470600 389292
rect 470652 389280 470658 389292
rect 471054 389280 471060 389292
rect 470652 389252 471060 389280
rect 470652 389240 470658 389252
rect 471054 389240 471060 389252
rect 471112 389240 471118 389292
rect 486418 389240 486424 389292
rect 486476 389280 486482 389292
rect 487062 389280 487068 389292
rect 486476 389252 487068 389280
rect 486476 389240 486482 389252
rect 487062 389240 487068 389252
rect 487120 389240 487126 389292
rect 497458 389240 497464 389292
rect 497516 389280 497522 389292
rect 498102 389280 498108 389292
rect 497516 389252 498108 389280
rect 497516 389240 497522 389252
rect 498102 389240 498108 389252
rect 498160 389240 498166 389292
rect 506474 389240 506480 389292
rect 506532 389280 506538 389292
rect 507118 389280 507124 389292
rect 506532 389252 507124 389280
rect 506532 389240 506538 389252
rect 507118 389240 507124 389252
rect 507176 389240 507182 389292
rect 507854 389240 507860 389292
rect 507912 389280 507918 389292
rect 508590 389280 508596 389292
rect 507912 389252 508596 389280
rect 507912 389240 507918 389252
rect 508590 389240 508596 389252
rect 508648 389240 508654 389292
rect 453022 389104 453028 389156
rect 453080 389144 453086 389156
rect 454034 389144 454040 389156
rect 453080 389116 454040 389144
rect 453080 389104 453086 389116
rect 454034 389104 454040 389116
rect 454092 389104 454098 389156
rect 456702 389104 456708 389156
rect 456760 389144 456766 389156
rect 457530 389144 457536 389156
rect 456760 389116 457536 389144
rect 456760 389104 456766 389116
rect 457530 389104 457536 389116
rect 457588 389104 457594 389156
rect 468478 389036 468484 389088
rect 468536 389076 468542 389088
rect 474366 389076 474372 389088
rect 468536 389048 474372 389076
rect 468536 389036 468542 389048
rect 474366 389036 474372 389048
rect 474424 389036 474430 389088
rect 467098 388968 467104 389020
rect 467156 389008 467162 389020
rect 475102 389008 475108 389020
rect 467156 388980 475108 389008
rect 467156 388968 467162 388980
rect 475102 388968 475108 388980
rect 475160 388968 475166 389020
rect 461118 388900 461124 388952
rect 461176 388940 461182 388952
rect 463602 388940 463608 388952
rect 461176 388912 463608 388940
rect 461176 388900 461182 388912
rect 463602 388900 463608 388912
rect 463660 388900 463666 388952
rect 468570 388900 468576 388952
rect 468628 388940 468634 388952
rect 478782 388940 478788 388952
rect 468628 388912 478788 388940
rect 468628 388900 468634 388912
rect 478782 388900 478788 388912
rect 478840 388900 478846 388952
rect 502334 388900 502340 388952
rect 502392 388940 502398 388952
rect 502392 388912 509234 388940
rect 502392 388900 502398 388912
rect 467190 388832 467196 388884
rect 467248 388872 467254 388884
rect 480254 388872 480260 388884
rect 467248 388844 480260 388872
rect 467248 388832 467254 388844
rect 480254 388832 480260 388844
rect 480312 388832 480318 388884
rect 483934 388832 483940 388884
rect 483992 388872 483998 388884
rect 502978 388872 502984 388884
rect 483992 388844 502984 388872
rect 483992 388832 483998 388844
rect 502978 388832 502984 388844
rect 503036 388832 503042 388884
rect 509206 388872 509234 388912
rect 526438 388872 526444 388884
rect 509206 388844 526444 388872
rect 526438 388832 526444 388844
rect 526496 388832 526502 388884
rect 461670 388764 461676 388816
rect 461728 388804 461734 388816
rect 475838 388804 475844 388816
rect 461728 388776 475844 388804
rect 461728 388764 461734 388776
rect 475838 388764 475844 388776
rect 475896 388764 475902 388816
rect 499390 388764 499396 388816
rect 499448 388804 499454 388816
rect 522298 388804 522304 388816
rect 499448 388776 522304 388804
rect 499448 388764 499454 388776
rect 522298 388764 522304 388776
rect 522356 388764 522362 388816
rect 464338 388696 464344 388748
rect 464396 388736 464402 388748
rect 478046 388736 478052 388748
rect 464396 388708 478052 388736
rect 464396 388696 464402 388708
rect 478046 388696 478052 388708
rect 478104 388696 478110 388748
rect 500862 388696 500868 388748
rect 500920 388736 500926 388748
rect 523678 388736 523684 388748
rect 500920 388708 523684 388736
rect 500920 388696 500926 388708
rect 523678 388696 523684 388708
rect 523736 388696 523742 388748
rect 462958 388628 462964 388680
rect 463016 388668 463022 388680
rect 476574 388668 476580 388680
rect 463016 388640 476580 388668
rect 463016 388628 463022 388640
rect 476574 388628 476580 388640
rect 476632 388628 476638 388680
rect 484670 388628 484676 388680
rect 484728 388668 484734 388680
rect 511350 388668 511356 388680
rect 484728 388640 511356 388668
rect 484728 388628 484734 388640
rect 511350 388628 511356 388640
rect 511408 388628 511414 388680
rect 465718 388560 465724 388612
rect 465776 388600 465782 388612
rect 480990 388600 480996 388612
rect 465776 388572 480996 388600
rect 465776 388560 465782 388572
rect 480990 388560 480996 388572
rect 481048 388560 481054 388612
rect 485406 388560 485412 388612
rect 485464 388600 485470 388612
rect 524414 388600 524420 388612
rect 485464 388572 524420 388600
rect 485464 388560 485470 388572
rect 524414 388560 524420 388572
rect 524472 388560 524478 388612
rect 447870 388492 447876 388544
rect 447928 388532 447934 388544
rect 458818 388532 458824 388544
rect 447928 388504 458824 388532
rect 447928 388492 447934 388504
rect 458818 388492 458824 388504
rect 458876 388492 458882 388544
rect 464522 388492 464528 388544
rect 464580 388532 464586 388544
rect 481726 388532 481732 388544
rect 464580 388504 481732 388532
rect 464580 388492 464586 388504
rect 481726 388492 481732 388504
rect 481784 388492 481790 388544
rect 489822 388492 489828 388544
rect 489880 388532 489886 388544
rect 530578 388532 530584 388544
rect 489880 388504 530584 388532
rect 489880 388492 489886 388504
rect 530578 388492 530584 388504
rect 530636 388492 530642 388544
rect 448330 388424 448336 388476
rect 448388 388464 448394 388476
rect 461762 388464 461768 388476
rect 448388 388436 461768 388464
rect 448388 388424 448394 388436
rect 461762 388424 461768 388436
rect 461820 388424 461826 388476
rect 463050 388424 463056 388476
rect 463108 388464 463114 388476
rect 482462 388464 482468 388476
rect 463108 388436 482468 388464
rect 463108 388424 463114 388436
rect 482462 388424 482468 388436
rect 482520 388424 482526 388476
rect 488350 388424 488356 388476
rect 488408 388464 488414 388476
rect 529198 388464 529204 388476
rect 488408 388436 529204 388464
rect 488408 388424 488414 388436
rect 529198 388424 529204 388436
rect 529256 388424 529262 388476
rect 461578 388016 461584 388068
rect 461636 388056 461642 388068
rect 462590 388056 462596 388068
rect 461636 388028 462596 388056
rect 461636 388016 461642 388028
rect 462590 388016 462596 388028
rect 462648 388016 462654 388068
rect 462130 387812 462136 387864
rect 462188 387852 462194 387864
rect 464890 387852 464896 387864
rect 462188 387824 464896 387852
rect 462188 387812 462194 387824
rect 464890 387812 464896 387824
rect 464948 387812 464954 387864
rect 428458 387744 428464 387796
rect 428516 387784 428522 387796
rect 431218 387784 431224 387796
rect 428516 387756 431224 387784
rect 428516 387744 428522 387756
rect 431218 387744 431224 387756
rect 431276 387744 431282 387796
rect 442718 387744 442724 387796
rect 442776 387784 442782 387796
rect 447134 387784 447140 387796
rect 442776 387756 447140 387784
rect 442776 387744 442782 387756
rect 447134 387744 447140 387756
rect 447192 387744 447198 387796
rect 450722 387336 450728 387388
rect 450780 387376 450786 387388
rect 454678 387376 454684 387388
rect 450780 387348 454684 387376
rect 450780 387336 450786 387348
rect 454678 387336 454684 387348
rect 454736 387336 454742 387388
rect 447410 387268 447416 387320
rect 447468 387308 447474 387320
rect 457438 387308 457444 387320
rect 447468 387280 457444 387308
rect 447468 387268 447474 387280
rect 457438 387268 457444 387280
rect 457496 387268 457502 387320
rect 447594 387200 447600 387252
rect 447652 387240 447658 387252
rect 461854 387240 461860 387252
rect 447652 387212 461860 387240
rect 447652 387200 447658 387212
rect 461854 387200 461860 387212
rect 461912 387200 461918 387252
rect 449802 387132 449808 387184
rect 449860 387172 449866 387184
rect 491294 387172 491300 387184
rect 449860 387144 491300 387172
rect 449860 387132 449866 387144
rect 491294 387132 491300 387144
rect 491352 387132 491358 387184
rect 441522 387064 441528 387116
rect 441580 387104 441586 387116
rect 447778 387104 447784 387116
rect 441580 387076 447784 387104
rect 441580 387064 441586 387076
rect 447778 387064 447784 387076
rect 447836 387064 447842 387116
rect 449434 387064 449440 387116
rect 449492 387104 449498 387116
rect 513374 387104 513380 387116
rect 449492 387076 513380 387104
rect 449492 387064 449498 387076
rect 513374 387064 513380 387076
rect 513432 387064 513438 387116
rect 448422 386588 448428 386640
rect 448480 386628 448486 386640
rect 553946 386628 553952 386640
rect 448480 386600 553952 386628
rect 448480 386588 448486 386600
rect 553946 386588 553952 386600
rect 554004 386588 554010 386640
rect 382918 386520 382924 386572
rect 382976 386560 382982 386572
rect 512086 386560 512092 386572
rect 382976 386532 512092 386560
rect 382976 386520 382982 386532
rect 512086 386520 512092 386532
rect 512144 386520 512150 386572
rect 374638 386452 374644 386504
rect 374696 386492 374702 386504
rect 512270 386492 512276 386504
rect 374696 386464 512276 386492
rect 374696 386452 374702 386464
rect 512270 386452 512276 386464
rect 512328 386452 512334 386504
rect 369118 386384 369124 386436
rect 369176 386424 369182 386436
rect 511994 386424 512000 386436
rect 369176 386396 512000 386424
rect 369176 386384 369182 386396
rect 511994 386384 512000 386396
rect 512052 386384 512058 386436
rect 448146 385976 448152 386028
rect 448204 386016 448210 386028
rect 453298 386016 453304 386028
rect 448204 385988 453304 386016
rect 448204 385976 448210 385988
rect 453298 385976 453304 385988
rect 453356 385976 453362 386028
rect 447962 385636 447968 385688
rect 448020 385676 448026 385688
rect 457346 385676 457352 385688
rect 448020 385648 457352 385676
rect 448020 385636 448026 385648
rect 457346 385636 457352 385648
rect 457404 385636 457410 385688
rect 448238 385364 448244 385416
rect 448296 385404 448302 385416
rect 452010 385404 452016 385416
rect 448296 385376 452016 385404
rect 448296 385364 448302 385376
rect 452010 385364 452016 385376
rect 452068 385364 452074 385416
rect 449342 385092 449348 385144
rect 449400 385132 449406 385144
rect 563422 385132 563428 385144
rect 449400 385104 563428 385132
rect 449400 385092 449406 385104
rect 563422 385092 563428 385104
rect 563480 385092 563486 385144
rect 373258 385024 373264 385076
rect 373316 385064 373322 385076
rect 512178 385064 512184 385076
rect 373316 385036 512184 385064
rect 373316 385024 373322 385036
rect 512178 385024 512184 385036
rect 512236 385024 512242 385076
rect 513282 383732 513288 383784
rect 513340 383772 513346 383784
rect 530578 383772 530584 383784
rect 513340 383744 530584 383772
rect 513340 383732 513346 383744
rect 530578 383732 530584 383744
rect 530636 383732 530642 383784
rect 512454 383664 512460 383716
rect 512512 383704 512518 383716
rect 548518 383704 548524 383716
rect 512512 383676 548524 383704
rect 512512 383664 512518 383676
rect 548518 383664 548524 383676
rect 548576 383664 548582 383716
rect 362218 383596 362224 383648
rect 362276 383636 362282 383648
rect 447134 383636 447140 383648
rect 362276 383608 447140 383636
rect 362276 383596 362282 383608
rect 447134 383596 447140 383608
rect 447192 383596 447198 383648
rect 378778 383528 378784 383580
rect 378836 383568 378842 383580
rect 447226 383568 447232 383580
rect 378836 383540 447232 383568
rect 378836 383528 378842 383540
rect 447226 383528 447232 383540
rect 447284 383528 447290 383580
rect 512638 382984 512644 383036
rect 512696 383024 512702 383036
rect 519722 383024 519728 383036
rect 512696 382996 519728 383024
rect 512696 382984 512702 382996
rect 519722 382984 519728 382996
rect 519780 382984 519786 383036
rect 513282 382576 513288 382628
rect 513340 382616 513346 382628
rect 518250 382616 518256 382628
rect 513340 382588 518256 382616
rect 513340 382576 513346 382588
rect 518250 382576 518256 382588
rect 518308 382576 518314 382628
rect 512454 382440 512460 382492
rect 512512 382480 512518 382492
rect 515582 382480 515588 382492
rect 512512 382452 515588 382480
rect 512512 382440 512518 382452
rect 515582 382440 515588 382452
rect 515640 382440 515646 382492
rect 374730 382168 374736 382220
rect 374788 382208 374794 382220
rect 447226 382208 447232 382220
rect 374788 382180 447232 382208
rect 374788 382168 374794 382180
rect 447226 382168 447232 382180
rect 447284 382168 447290 382220
rect 376018 382100 376024 382152
rect 376076 382140 376082 382152
rect 447134 382140 447140 382152
rect 376076 382112 447140 382140
rect 376076 382100 376082 382112
rect 447134 382100 447140 382112
rect 447192 382100 447198 382152
rect 361574 380876 361580 380928
rect 361632 380916 361638 380928
rect 443822 380916 443828 380928
rect 361632 380888 443828 380916
rect 361632 380876 361638 380888
rect 443822 380876 443828 380888
rect 443880 380876 443886 380928
rect 512454 380876 512460 380928
rect 512512 380916 512518 380928
rect 547138 380916 547144 380928
rect 512512 380888 547144 380916
rect 512512 380876 512518 380888
rect 547138 380876 547144 380888
rect 547196 380876 547202 380928
rect 363598 380808 363604 380860
rect 363656 380848 363662 380860
rect 447502 380848 447508 380860
rect 363656 380820 447508 380848
rect 363656 380808 363662 380820
rect 447502 380808 447508 380820
rect 447560 380808 447566 380860
rect 371878 380740 371884 380792
rect 371936 380780 371942 380792
rect 447134 380780 447140 380792
rect 371936 380752 447140 380780
rect 371936 380740 371942 380752
rect 447134 380740 447140 380752
rect 447192 380740 447198 380792
rect 400858 380672 400864 380724
rect 400916 380712 400922 380724
rect 447226 380712 447232 380724
rect 400916 380684 447232 380712
rect 400916 380672 400922 380684
rect 447226 380672 447232 380684
rect 447284 380672 447290 380724
rect 512546 379720 512552 379772
rect 512604 379760 512610 379772
rect 515674 379760 515680 379772
rect 512604 379732 515680 379760
rect 512604 379720 512610 379732
rect 515674 379720 515680 379732
rect 515732 379720 515738 379772
rect 513282 379516 513288 379568
rect 513340 379556 513346 379568
rect 549898 379556 549904 379568
rect 513340 379528 549904 379556
rect 513340 379516 513346 379528
rect 549898 379516 549904 379528
rect 549956 379516 549962 379568
rect 363690 379448 363696 379500
rect 363748 379488 363754 379500
rect 447318 379488 447324 379500
rect 363748 379460 447324 379488
rect 363748 379448 363754 379460
rect 447318 379448 447324 379460
rect 447376 379448 447382 379500
rect 370498 379380 370504 379432
rect 370556 379420 370562 379432
rect 447134 379420 447140 379432
rect 370556 379392 447140 379420
rect 370556 379380 370562 379392
rect 447134 379380 447140 379392
rect 447192 379380 447198 379432
rect 513282 378292 513288 378344
rect 513340 378332 513346 378344
rect 522298 378332 522304 378344
rect 513340 378304 522304 378332
rect 513340 378292 513346 378304
rect 522298 378292 522304 378304
rect 522356 378292 522362 378344
rect 512822 378224 512828 378276
rect 512880 378264 512886 378276
rect 547230 378264 547236 378276
rect 512880 378236 547236 378264
rect 512880 378224 512886 378236
rect 547230 378224 547236 378236
rect 547288 378224 547294 378276
rect 514018 378156 514024 378208
rect 514076 378196 514082 378208
rect 580166 378196 580172 378208
rect 514076 378168 580172 378196
rect 514076 378156 514082 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 363782 378088 363788 378140
rect 363840 378128 363846 378140
rect 447226 378128 447232 378140
rect 363840 378100 447232 378128
rect 363840 378088 363846 378100
rect 447226 378088 447232 378100
rect 447284 378088 447290 378140
rect 367738 378020 367744 378072
rect 367796 378060 367802 378072
rect 447134 378060 447140 378072
rect 367796 378032 447140 378060
rect 367796 378020 367802 378032
rect 447134 378020 447140 378032
rect 447192 378020 447198 378072
rect 513190 377408 513196 377460
rect 513248 377448 513254 377460
rect 548610 377448 548616 377460
rect 513248 377420 548616 377448
rect 513248 377408 513254 377420
rect 548610 377408 548616 377420
rect 548668 377408 548674 377460
rect 512822 376728 512828 376780
rect 512880 376768 512886 376780
rect 516226 376768 516232 376780
rect 512880 376740 516232 376768
rect 512880 376728 512886 376740
rect 516226 376728 516232 376740
rect 516284 376728 516290 376780
rect 403618 376660 403624 376712
rect 403676 376700 403682 376712
rect 447134 376700 447140 376712
rect 403676 376672 447140 376700
rect 403676 376660 403682 376672
rect 447134 376660 447140 376672
rect 447192 376660 447198 376712
rect 419074 376592 419080 376644
rect 419132 376632 419138 376644
rect 447226 376632 447232 376644
rect 419132 376604 447232 376632
rect 419132 376592 419138 376604
rect 447226 376592 447232 376604
rect 447284 376592 447290 376644
rect 513098 375980 513104 376032
rect 513156 376020 513162 376032
rect 544378 376020 544384 376032
rect 513156 375992 544384 376020
rect 513156 375980 513162 375992
rect 544378 375980 544384 375992
rect 544436 375980 544442 376032
rect 513282 375912 513288 375964
rect 513340 375952 513346 375964
rect 518894 375952 518900 375964
rect 513340 375924 518900 375952
rect 513340 375912 513346 375924
rect 518894 375912 518900 375924
rect 518952 375912 518958 375964
rect 513282 375368 513288 375420
rect 513340 375408 513346 375420
rect 518342 375408 518348 375420
rect 513340 375380 518348 375408
rect 513340 375368 513346 375380
rect 518342 375368 518348 375380
rect 518400 375368 518406 375420
rect 406378 375300 406384 375352
rect 406436 375340 406442 375352
rect 447134 375340 447140 375352
rect 406436 375312 447140 375340
rect 406436 375300 406442 375312
rect 447134 375300 447140 375312
rect 447192 375300 447198 375352
rect 407758 375232 407764 375284
rect 407816 375272 407822 375284
rect 447226 375272 447232 375284
rect 407816 375244 447232 375272
rect 407816 375232 407822 375244
rect 447226 375232 447232 375244
rect 447284 375232 447290 375284
rect 512086 374008 512092 374060
rect 512144 374048 512150 374060
rect 520274 374048 520280 374060
rect 512144 374020 520280 374048
rect 512144 374008 512150 374020
rect 520274 374008 520280 374020
rect 520332 374008 520338 374060
rect 410518 373940 410524 373992
rect 410576 373980 410582 373992
rect 447134 373980 447140 373992
rect 410576 373952 447140 373980
rect 410576 373940 410582 373952
rect 447134 373940 447140 373952
rect 447192 373940 447198 373992
rect 411898 373872 411904 373924
rect 411956 373912 411962 373924
rect 447226 373912 447232 373924
rect 411956 373884 447232 373912
rect 411956 373872 411962 373884
rect 447226 373872 447232 373884
rect 447284 373872 447290 373924
rect 512454 372716 512460 372768
rect 512512 372756 512518 372768
rect 521654 372756 521660 372768
rect 512512 372728 521660 372756
rect 512512 372716 512518 372728
rect 521654 372716 521660 372728
rect 521712 372716 521718 372768
rect 512086 372648 512092 372700
rect 512144 372688 512150 372700
rect 514754 372688 514760 372700
rect 512144 372660 514760 372688
rect 512144 372648 512150 372660
rect 514754 372648 514760 372660
rect 514812 372648 514818 372700
rect 511994 372580 512000 372632
rect 512052 372620 512058 372632
rect 514846 372620 514852 372632
rect 512052 372592 514852 372620
rect 512052 372580 512058 372592
rect 514846 372580 514852 372592
rect 514904 372580 514910 372632
rect 381538 372512 381544 372564
rect 381596 372552 381602 372564
rect 447134 372552 447140 372564
rect 381596 372524 447140 372552
rect 381596 372512 381602 372524
rect 447134 372512 447140 372524
rect 447192 372512 447198 372564
rect 419166 372444 419172 372496
rect 419224 372484 419230 372496
rect 447226 372484 447232 372496
rect 419224 372456 447232 372484
rect 419224 372444 419230 372456
rect 447226 372444 447232 372456
rect 447284 372444 447290 372496
rect 512454 371900 512460 371952
rect 512512 371940 512518 371952
rect 516318 371940 516324 371952
rect 512512 371912 516324 371940
rect 512512 371900 512518 371912
rect 516318 371900 516324 371912
rect 516376 371900 516382 371952
rect 396718 371152 396724 371204
rect 396776 371192 396782 371204
rect 447134 371192 447140 371204
rect 396776 371164 447140 371192
rect 396776 371152 396782 371164
rect 447134 371152 447140 371164
rect 447192 371152 447198 371204
rect 414658 371084 414664 371136
rect 414716 371124 414722 371136
rect 447226 371124 447232 371136
rect 414716 371096 447232 371124
rect 414716 371084 414722 371096
rect 447226 371084 447232 371096
rect 447284 371084 447290 371136
rect 512454 370336 512460 370388
rect 512512 370376 512518 370388
rect 517606 370376 517612 370388
rect 512512 370348 517612 370376
rect 512512 370336 512518 370348
rect 517606 370336 517612 370348
rect 517664 370336 517670 370388
rect 512822 369928 512828 369980
rect 512880 369968 512886 369980
rect 516870 369968 516876 369980
rect 512880 369940 516876 369968
rect 512880 369928 512886 369940
rect 516870 369928 516876 369940
rect 516928 369928 516934 369980
rect 361574 369860 361580 369912
rect 361632 369900 361638 369912
rect 409874 369900 409880 369912
rect 361632 369872 409880 369900
rect 361632 369860 361638 369872
rect 409874 369860 409880 369872
rect 409932 369860 409938 369912
rect 513282 369860 513288 369912
rect 513340 369900 513346 369912
rect 523034 369900 523040 369912
rect 513340 369872 523040 369900
rect 513340 369860 513346 369872
rect 523034 369860 523040 369872
rect 523092 369860 523098 369912
rect 399478 369792 399484 369844
rect 399536 369832 399542 369844
rect 447134 369832 447140 369844
rect 399536 369804 447140 369832
rect 399536 369792 399542 369804
rect 447134 369792 447140 369804
rect 447192 369792 447198 369844
rect 416130 369724 416136 369776
rect 416188 369764 416194 369776
rect 447226 369764 447232 369776
rect 416188 369736 447232 369764
rect 416188 369724 416194 369736
rect 447226 369724 447232 369736
rect 447284 369724 447290 369776
rect 431218 369656 431224 369708
rect 431276 369696 431282 369708
rect 432874 369696 432880 369708
rect 431276 369668 432880 369696
rect 431276 369656 431282 369668
rect 432874 369656 432880 369668
rect 432932 369656 432938 369708
rect 512822 368568 512828 368620
rect 512880 368608 512886 368620
rect 516410 368608 516416 368620
rect 512880 368580 516416 368608
rect 512880 368568 512886 368580
rect 516410 368568 516416 368580
rect 516468 368568 516474 368620
rect 513282 368500 513288 368552
rect 513340 368540 513346 368552
rect 520366 368540 520372 368552
rect 513340 368512 520372 368540
rect 513340 368500 513346 368512
rect 520366 368500 520372 368512
rect 520424 368500 520430 368552
rect 417418 368432 417424 368484
rect 417476 368472 417482 368484
rect 447134 368472 447140 368484
rect 417476 368444 447140 368472
rect 417476 368432 417482 368444
rect 447134 368432 447140 368444
rect 447192 368432 447198 368484
rect 443638 368364 443644 368416
rect 443696 368404 443702 368416
rect 447226 368404 447232 368416
rect 443696 368376 447232 368404
rect 443696 368364 443702 368376
rect 447226 368364 447232 368376
rect 447284 368364 447290 368416
rect 513282 367208 513288 367260
rect 513340 367248 513346 367260
rect 517974 367248 517980 367260
rect 513340 367220 517980 367248
rect 513340 367208 513346 367220
rect 517974 367208 517980 367220
rect 518032 367208 518038 367260
rect 511994 367072 512000 367124
rect 512052 367112 512058 367124
rect 514110 367112 514116 367124
rect 512052 367084 514116 367112
rect 512052 367072 512058 367084
rect 514110 367072 514116 367084
rect 514168 367072 514174 367124
rect 439498 367004 439504 367056
rect 439556 367044 439562 367056
rect 447134 367044 447140 367056
rect 439556 367016 447140 367044
rect 439556 367004 439562 367016
rect 447134 367004 447140 367016
rect 447192 367004 447198 367056
rect 443730 366936 443736 366988
rect 443788 366976 443794 366988
rect 447226 366976 447232 366988
rect 443788 366948 447232 366976
rect 443788 366936 443794 366948
rect 447226 366936 447232 366948
rect 447284 366936 447290 366988
rect 511994 365848 512000 365900
rect 512052 365888 512058 365900
rect 514202 365888 514208 365900
rect 512052 365860 514208 365888
rect 512052 365848 512058 365860
rect 514202 365848 514208 365860
rect 514260 365848 514266 365900
rect 513282 365712 513288 365764
rect 513340 365752 513346 365764
rect 521746 365752 521752 365764
rect 513340 365724 521752 365752
rect 513340 365712 513346 365724
rect 521746 365712 521752 365724
rect 521804 365712 521810 365764
rect 409874 365644 409880 365696
rect 409932 365684 409938 365696
rect 447134 365684 447140 365696
rect 409932 365656 447140 365684
rect 409932 365644 409938 365656
rect 447134 365644 447140 365656
rect 447192 365644 447198 365696
rect 443822 365576 443828 365628
rect 443880 365616 443886 365628
rect 447226 365616 447232 365628
rect 443880 365588 447232 365616
rect 443880 365576 443886 365588
rect 447226 365576 447232 365588
rect 447284 365576 447290 365628
rect 512638 365168 512644 365220
rect 512696 365208 512702 365220
rect 520458 365208 520464 365220
rect 512696 365180 520464 365208
rect 512696 365168 512702 365180
rect 520458 365168 520464 365180
rect 520516 365168 520522 365220
rect 513282 364352 513288 364404
rect 513340 364392 513346 364404
rect 523126 364392 523132 364404
rect 513340 364364 523132 364392
rect 513340 364352 513346 364364
rect 523126 364352 523132 364364
rect 523184 364352 523190 364404
rect 576210 364352 576216 364404
rect 576268 364392 576274 364404
rect 580166 364392 580172 364404
rect 576268 364364 580172 364392
rect 576268 364352 576274 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 432690 362992 432696 363044
rect 432748 363032 432754 363044
rect 447134 363032 447140 363044
rect 432748 363004 447140 363032
rect 432748 362992 432754 363004
rect 447134 362992 447140 363004
rect 447192 362992 447198 363044
rect 512454 362992 512460 363044
rect 512512 363032 512518 363044
rect 521838 363032 521844 363044
rect 512512 363004 521844 363032
rect 512512 362992 512518 363004
rect 521838 362992 521844 363004
rect 521896 362992 521902 363044
rect 432782 362924 432788 362976
rect 432840 362964 432846 362976
rect 447226 362964 447232 362976
rect 432840 362936 447232 362964
rect 432840 362924 432846 362936
rect 447226 362924 447232 362936
rect 447284 362924 447290 362976
rect 511994 362312 512000 362364
rect 512052 362352 512058 362364
rect 513650 362352 513656 362364
rect 512052 362324 513656 362352
rect 512052 362312 512058 362324
rect 513650 362312 513656 362324
rect 513708 362312 513714 362364
rect 442258 361632 442264 361684
rect 442316 361672 442322 361684
rect 447226 361672 447232 361684
rect 442316 361644 447232 361672
rect 442316 361632 442322 361644
rect 447226 361632 447232 361644
rect 447284 361632 447290 361684
rect 432598 361564 432604 361616
rect 432656 361604 432662 361616
rect 447134 361604 447140 361616
rect 432656 361576 447140 361604
rect 432656 361564 432662 361576
rect 447134 361564 447140 361576
rect 447192 361564 447198 361616
rect 513006 361564 513012 361616
rect 513064 361604 513070 361616
rect 520550 361604 520556 361616
rect 513064 361576 520556 361604
rect 513064 361564 513070 361576
rect 520550 361564 520556 361576
rect 520608 361564 520614 361616
rect 512914 360952 512920 361004
rect 512972 360992 512978 361004
rect 518986 360992 518992 361004
rect 512972 360964 518992 360992
rect 512972 360952 512978 360964
rect 518986 360952 518992 360964
rect 519044 360952 519050 361004
rect 512362 360680 512368 360732
rect 512420 360720 512426 360732
rect 515030 360720 515036 360732
rect 512420 360692 515036 360720
rect 512420 360680 512426 360692
rect 515030 360680 515036 360692
rect 515088 360680 515094 360732
rect 513190 360544 513196 360596
rect 513248 360584 513254 360596
rect 517698 360584 517704 360596
rect 513248 360556 517704 360584
rect 513248 360544 513254 360556
rect 517698 360544 517704 360556
rect 517756 360544 517762 360596
rect 439774 360272 439780 360324
rect 439832 360312 439838 360324
rect 447226 360312 447232 360324
rect 439832 360284 447232 360312
rect 439832 360272 439838 360284
rect 447226 360272 447232 360284
rect 447284 360272 447290 360324
rect 436922 360204 436928 360256
rect 436980 360244 436986 360256
rect 447134 360244 447140 360256
rect 436980 360216 447140 360244
rect 436980 360204 436986 360216
rect 447134 360204 447140 360216
rect 447192 360204 447198 360256
rect 547230 360136 547236 360188
rect 547288 360176 547294 360188
rect 552014 360176 552020 360188
rect 547288 360148 552020 360176
rect 547288 360136 547294 360148
rect 552014 360136 552020 360148
rect 552072 360136 552078 360188
rect 530578 360068 530584 360120
rect 530636 360108 530642 360120
rect 566734 360108 566740 360120
rect 530636 360080 566740 360108
rect 530636 360068 530642 360080
rect 566734 360068 566740 360080
rect 566792 360068 566798 360120
rect 522298 360000 522304 360052
rect 522356 360040 522362 360052
rect 550634 360040 550640 360052
rect 522356 360012 550640 360040
rect 522356 360000 522362 360012
rect 550634 360000 550640 360012
rect 550692 360000 550698 360052
rect 549898 359932 549904 359984
rect 549956 359972 549962 359984
rect 554958 359972 554964 359984
rect 549956 359944 554964 359972
rect 549956 359932 549962 359944
rect 554958 359932 554964 359944
rect 555016 359932 555022 359984
rect 565262 359972 565268 359984
rect 563026 359944 565268 359972
rect 547138 359864 547144 359916
rect 547196 359904 547202 359916
rect 558178 359904 558184 359916
rect 547196 359876 558184 359904
rect 547196 359864 547202 359876
rect 558178 359864 558184 359876
rect 558236 359864 558242 359916
rect 515674 359796 515680 359848
rect 515732 359836 515738 359848
rect 553762 359836 553768 359848
rect 515732 359808 553768 359836
rect 515732 359796 515738 359808
rect 553762 359796 553768 359808
rect 553820 359796 553826 359848
rect 548518 359728 548524 359780
rect 548576 359768 548582 359780
rect 563026 359768 563054 359944
rect 565262 359932 565268 359944
rect 565320 359932 565326 359984
rect 548576 359740 563054 359768
rect 548576 359728 548582 359740
rect 443822 358844 443828 358896
rect 443880 358884 443886 358896
rect 447226 358884 447232 358896
rect 443880 358856 447232 358884
rect 443880 358844 443886 358856
rect 447226 358844 447232 358856
rect 447284 358844 447290 358896
rect 435450 358776 435456 358828
rect 435508 358816 435514 358828
rect 447134 358816 447140 358828
rect 435508 358788 447140 358816
rect 435508 358776 435514 358788
rect 447134 358776 447140 358788
rect 447192 358776 447198 358828
rect 512730 358776 512736 358828
rect 512788 358816 512794 358828
rect 517882 358816 517888 358828
rect 512788 358788 517888 358816
rect 512788 358776 512794 358788
rect 517882 358776 517888 358788
rect 517940 358776 517946 358828
rect 548610 358708 548616 358760
rect 548668 358748 548674 358760
rect 556706 358748 556712 358760
rect 548668 358720 556712 358748
rect 548668 358708 548674 358720
rect 556706 358708 556712 358720
rect 556764 358708 556770 358760
rect 518250 358640 518256 358692
rect 518308 358680 518314 358692
rect 562594 358680 562600 358692
rect 518308 358652 562600 358680
rect 518308 358640 518314 358652
rect 562594 358640 562600 358652
rect 562652 358640 562658 358692
rect 519722 358572 519728 358624
rect 519780 358612 519786 358624
rect 564066 358612 564072 358624
rect 519780 358584 564072 358612
rect 519780 358572 519786 358584
rect 564066 358572 564072 358584
rect 564124 358572 564130 358624
rect 544378 358504 544384 358556
rect 544436 358544 544442 358556
rect 559650 358544 559656 358556
rect 544436 358516 559656 358544
rect 544436 358504 544442 358516
rect 559650 358504 559656 358516
rect 559708 358504 559714 358556
rect 515582 358436 515588 358488
rect 515640 358476 515646 358488
rect 561122 358476 561128 358488
rect 515640 358448 561128 358476
rect 515640 358436 515646 358448
rect 561122 358436 561128 358448
rect 561180 358436 561186 358488
rect 513282 357824 513288 357876
rect 513340 357864 513346 357876
rect 519078 357864 519084 357876
rect 513340 357836 519084 357864
rect 513340 357824 513346 357836
rect 519078 357824 519084 357836
rect 519136 357824 519142 357876
rect 513282 356056 513288 356108
rect 513340 356096 513346 356108
rect 523218 356096 523224 356108
rect 513340 356068 523224 356096
rect 513340 356056 513346 356068
rect 523218 356056 523224 356068
rect 523276 356056 523282 356108
rect 513282 354968 513288 355020
rect 513340 355008 513346 355020
rect 519170 355008 519176 355020
rect 513340 354980 519176 355008
rect 513340 354968 513346 354980
rect 519170 354968 519176 354980
rect 519228 354968 519234 355020
rect 511994 353948 512000 354000
rect 512052 353988 512058 354000
rect 513742 353988 513748 354000
rect 512052 353960 513748 353988
rect 512052 353948 512058 353960
rect 513742 353948 513748 353960
rect 513800 353948 513806 354000
rect 513282 353472 513288 353524
rect 513340 353512 513346 353524
rect 517790 353512 517796 353524
rect 513340 353484 517796 353512
rect 513340 353472 513346 353484
rect 517790 353472 517796 353484
rect 517848 353472 517854 353524
rect 445662 353268 445668 353320
rect 445720 353308 445726 353320
rect 447870 353308 447876 353320
rect 445720 353280 447876 353308
rect 445720 353268 445726 353280
rect 447870 353268 447876 353280
rect 447928 353268 447934 353320
rect 446214 353064 446220 353116
rect 446272 353104 446278 353116
rect 447778 353104 447784 353116
rect 446272 353076 447784 353104
rect 446272 353064 446278 353076
rect 447778 353064 447784 353076
rect 447836 353064 447842 353116
rect 511994 352384 512000 352436
rect 512052 352424 512058 352436
rect 515122 352424 515128 352436
rect 512052 352396 515128 352424
rect 512052 352384 512058 352396
rect 515122 352384 515128 352396
rect 515180 352384 515186 352436
rect 513282 351908 513288 351960
rect 513340 351948 513346 351960
rect 521930 351948 521936 351960
rect 513340 351920 521936 351948
rect 513340 351908 513346 351920
rect 521930 351908 521936 351920
rect 521988 351908 521994 351960
rect 512638 350888 512644 350940
rect 512696 350928 512702 350940
rect 519354 350928 519360 350940
rect 512696 350900 519360 350928
rect 512696 350888 512702 350900
rect 519354 350888 519360 350900
rect 519412 350888 519418 350940
rect 512546 350616 512552 350668
rect 512604 350656 512610 350668
rect 515214 350656 515220 350668
rect 512604 350628 515220 350656
rect 512604 350616 512610 350628
rect 515214 350616 515220 350628
rect 515272 350616 515278 350668
rect 407022 350548 407028 350600
rect 407080 350588 407086 350600
rect 447134 350588 447140 350600
rect 407080 350560 447140 350588
rect 407080 350548 407086 350560
rect 447134 350548 447140 350560
rect 447192 350548 447198 350600
rect 513282 349528 513288 349580
rect 513340 349568 513346 349580
rect 519446 349568 519452 349580
rect 513340 349540 519452 349568
rect 513340 349528 513346 349540
rect 519446 349528 519452 349540
rect 519504 349528 519510 349580
rect 511994 349392 512000 349444
rect 512052 349432 512058 349444
rect 514938 349432 514944 349444
rect 512052 349404 514944 349432
rect 512052 349392 512058 349404
rect 514938 349392 514944 349404
rect 514996 349392 515002 349444
rect 511994 349256 512000 349308
rect 512052 349296 512058 349308
rect 513834 349296 513840 349308
rect 512052 349268 513840 349296
rect 512052 349256 512058 349268
rect 513834 349256 513840 349268
rect 513892 349256 513898 349308
rect 432874 349052 432880 349104
rect 432932 349092 432938 349104
rect 437014 349092 437020 349104
rect 432932 349064 437020 349092
rect 432932 349052 432938 349064
rect 437014 349052 437020 349064
rect 437072 349052 437078 349104
rect 512914 348032 512920 348084
rect 512972 348072 512978 348084
rect 516502 348072 516508 348084
rect 512972 348044 516508 348072
rect 512972 348032 512978 348044
rect 516502 348032 516508 348044
rect 516560 348032 516566 348084
rect 361758 347760 361764 347812
rect 361816 347800 361822 347812
rect 402238 347800 402244 347812
rect 361816 347772 402244 347800
rect 361816 347760 361822 347772
rect 402238 347760 402244 347772
rect 402296 347760 402302 347812
rect 513282 347760 513288 347812
rect 513340 347800 513346 347812
rect 523310 347800 523316 347812
rect 513340 347772 523316 347800
rect 513340 347760 513346 347772
rect 523310 347760 523316 347772
rect 523368 347760 523374 347812
rect 362218 347692 362224 347744
rect 362276 347732 362282 347744
rect 447134 347732 447140 347744
rect 362276 347704 447140 347732
rect 362276 347692 362282 347704
rect 447134 347692 447140 347704
rect 447192 347692 447198 347744
rect 513282 346944 513288 346996
rect 513340 346984 513346 346996
rect 519262 346984 519268 346996
rect 513340 346956 519268 346984
rect 513340 346944 513346 346956
rect 519262 346944 519268 346956
rect 519320 346944 519326 346996
rect 512546 346536 512552 346588
rect 512604 346576 512610 346588
rect 515306 346576 515312 346588
rect 512604 346548 515312 346576
rect 512604 346536 512610 346548
rect 515306 346536 515312 346548
rect 515364 346536 515370 346588
rect 513282 346468 513288 346520
rect 513340 346508 513346 346520
rect 518066 346508 518072 346520
rect 513340 346480 518072 346508
rect 513340 346468 513346 346480
rect 518066 346468 518072 346480
rect 518124 346468 518130 346520
rect 513006 343816 513012 343868
rect 513064 343856 513070 343868
rect 516686 343856 516692 343868
rect 513064 343828 516692 343856
rect 513064 343816 513070 343828
rect 516686 343816 516692 343828
rect 516744 343816 516750 343868
rect 512822 343748 512828 343800
rect 512880 343788 512886 343800
rect 517514 343788 517520 343800
rect 512880 343760 517520 343788
rect 512880 343748 512886 343760
rect 517514 343748 517520 343760
rect 517572 343748 517578 343800
rect 513006 342320 513012 342372
rect 513064 342360 513070 342372
rect 516778 342360 516784 342372
rect 513064 342332 516784 342360
rect 513064 342320 513070 342332
rect 516778 342320 516784 342332
rect 516836 342320 516842 342372
rect 513282 341368 513288 341420
rect 513340 341408 513346 341420
rect 520642 341408 520648 341420
rect 513340 341380 520648 341408
rect 513340 341368 513346 341380
rect 520642 341368 520648 341380
rect 520700 341368 520706 341420
rect 513282 341096 513288 341148
rect 513340 341136 513346 341148
rect 518250 341136 518256 341148
rect 513340 341108 518256 341136
rect 513340 341096 513346 341108
rect 518250 341096 518256 341108
rect 518308 341096 518314 341148
rect 444190 340960 444196 341012
rect 444248 341000 444254 341012
rect 447226 341000 447232 341012
rect 444248 340972 447232 341000
rect 444248 340960 444254 340972
rect 447226 340960 447232 340972
rect 447284 340960 447290 341012
rect 361758 340892 361764 340944
rect 361816 340932 361822 340944
rect 447134 340932 447140 340944
rect 361816 340904 447140 340932
rect 361816 340892 361822 340904
rect 447134 340892 447140 340904
rect 447192 340892 447198 340944
rect 512638 339736 512644 339788
rect 512696 339776 512702 339788
rect 516134 339776 516140 339788
rect 512696 339748 516140 339776
rect 512696 339736 512702 339748
rect 516134 339736 516140 339748
rect 516192 339736 516198 339788
rect 431218 339532 431224 339584
rect 431276 339572 431282 339584
rect 447134 339572 447140 339584
rect 431276 339544 447140 339572
rect 431276 339532 431282 339544
rect 447134 339532 447140 339544
rect 447192 339532 447198 339584
rect 371878 339464 371884 339516
rect 371936 339504 371942 339516
rect 447226 339504 447232 339516
rect 371936 339476 447232 339504
rect 371936 339464 371942 339476
rect 447226 339464 447232 339476
rect 447284 339464 447290 339516
rect 512638 339464 512644 339516
rect 512696 339504 512702 339516
rect 515582 339504 515588 339516
rect 512696 339476 515588 339504
rect 512696 339464 512702 339476
rect 515582 339464 515588 339476
rect 515640 339464 515646 339516
rect 513006 338376 513012 338428
rect 513064 338416 513070 338428
rect 516594 338416 516600 338428
rect 513064 338388 516600 338416
rect 513064 338376 513070 338388
rect 516594 338376 516600 338388
rect 516652 338376 516658 338428
rect 436830 338172 436836 338224
rect 436888 338212 436894 338224
rect 447134 338212 447140 338224
rect 436888 338184 447140 338212
rect 436888 338172 436894 338184
rect 447134 338172 447140 338184
rect 447192 338172 447198 338224
rect 435358 338104 435364 338156
rect 435416 338144 435422 338156
rect 447226 338144 447232 338156
rect 435416 338116 447232 338144
rect 435416 338104 435422 338116
rect 447226 338104 447232 338116
rect 447284 338104 447290 338156
rect 450078 337968 450084 338020
rect 450136 338008 450142 338020
rect 450354 338008 450360 338020
rect 450136 337980 450360 338008
rect 450136 337968 450142 337980
rect 450354 337968 450360 337980
rect 450412 337968 450418 338020
rect 402238 337356 402244 337408
rect 402296 337396 402302 337408
rect 447870 337396 447876 337408
rect 402296 337368 447876 337396
rect 402296 337356 402302 337368
rect 447870 337356 447876 337368
rect 447928 337396 447934 337408
rect 448422 337396 448428 337408
rect 447928 337368 448428 337396
rect 447928 337356 447934 337368
rect 448422 337356 448428 337368
rect 448480 337356 448486 337408
rect 513190 337288 513196 337340
rect 513248 337328 513254 337340
rect 519722 337328 519728 337340
rect 513248 337300 519728 337328
rect 513248 337288 513254 337300
rect 519722 337288 519728 337300
rect 519780 337288 519786 337340
rect 513282 337152 513288 337204
rect 513340 337192 513346 337204
rect 520918 337192 520924 337204
rect 513340 337164 520924 337192
rect 513340 337152 513346 337164
rect 520918 337152 520924 337164
rect 520976 337152 520982 337204
rect 440878 336948 440884 337000
rect 440936 336988 440942 337000
rect 447134 336988 447140 337000
rect 440936 336960 447140 336988
rect 440936 336948 440942 336960
rect 447134 336948 447140 336960
rect 447192 336948 447198 337000
rect 416774 336880 416780 336932
rect 416832 336920 416838 336932
rect 450354 336920 450360 336932
rect 416832 336892 450360 336920
rect 416832 336880 416838 336892
rect 450354 336880 450360 336892
rect 450412 336880 450418 336932
rect 413094 336812 413100 336864
rect 413152 336852 413158 336864
rect 450170 336852 450176 336864
rect 413152 336824 450176 336852
rect 413152 336812 413158 336824
rect 450170 336812 450176 336824
rect 450228 336812 450234 336864
rect 409414 336744 409420 336796
rect 409472 336784 409478 336796
rect 450722 336784 450728 336796
rect 409472 336756 450728 336784
rect 409472 336744 409478 336756
rect 450722 336744 450728 336756
rect 450780 336744 450786 336796
rect 418890 336336 418896 336388
rect 418948 336376 418954 336388
rect 440970 336376 440976 336388
rect 418948 336348 440976 336376
rect 418948 336336 418954 336348
rect 440970 336336 440976 336348
rect 441028 336336 441034 336388
rect 418982 336268 418988 336320
rect 419040 336308 419046 336320
rect 441246 336308 441252 336320
rect 419040 336280 441252 336308
rect 419040 336268 419046 336280
rect 441246 336268 441252 336280
rect 441304 336268 441310 336320
rect 418798 336200 418804 336252
rect 418856 336240 418862 336252
rect 441154 336240 441160 336252
rect 418856 336212 441160 336240
rect 418856 336200 418862 336212
rect 441154 336200 441160 336212
rect 441212 336200 441218 336252
rect 416038 336132 416044 336184
rect 416096 336172 416102 336184
rect 441062 336172 441068 336184
rect 416096 336144 441068 336172
rect 416096 336132 416102 336144
rect 441062 336132 441068 336144
rect 441120 336132 441126 336184
rect 413646 336064 413652 336116
rect 413704 336104 413710 336116
rect 449434 336104 449440 336116
rect 413704 336076 449440 336104
rect 413704 336064 413710 336076
rect 449434 336064 449440 336076
rect 449492 336064 449498 336116
rect 362218 335996 362224 336048
rect 362276 336036 362282 336048
rect 444190 336036 444196 336048
rect 362276 336008 444196 336036
rect 362276 335996 362282 336008
rect 444190 335996 444196 336008
rect 444248 335996 444254 336048
rect 443730 335656 443736 335708
rect 443788 335696 443794 335708
rect 447226 335696 447232 335708
rect 443788 335668 447232 335696
rect 443788 335656 443794 335668
rect 447226 335656 447232 335668
rect 447284 335656 447290 335708
rect 399478 335316 399484 335368
rect 399536 335356 399542 335368
rect 447134 335356 447140 335368
rect 399536 335328 447140 335356
rect 399536 335316 399542 335328
rect 447134 335316 447140 335328
rect 447192 335316 447198 335368
rect 439682 335044 439688 335096
rect 439740 335084 439746 335096
rect 447502 335084 447508 335096
rect 439740 335056 447508 335084
rect 439740 335044 439746 335056
rect 447502 335044 447508 335056
rect 447560 335044 447566 335096
rect 420546 334976 420552 335028
rect 420604 335016 420610 335028
rect 439866 335016 439872 335028
rect 420604 334988 439872 335016
rect 420604 334976 420610 334988
rect 439866 334976 439872 334988
rect 439924 334976 439930 335028
rect 420822 334908 420828 334960
rect 420880 334948 420886 334960
rect 442350 334948 442356 334960
rect 420880 334920 442356 334948
rect 420880 334908 420886 334920
rect 442350 334908 442356 334920
rect 442408 334908 442414 334960
rect 420270 334840 420276 334892
rect 420328 334880 420334 334892
rect 442442 334880 442448 334892
rect 420328 334852 442448 334880
rect 420328 334840 420334 334852
rect 442442 334840 442448 334852
rect 442500 334840 442506 334892
rect 513282 334840 513288 334892
rect 513340 334880 513346 334892
rect 520734 334880 520740 334892
rect 513340 334852 520740 334880
rect 513340 334840 513346 334852
rect 520734 334840 520740 334852
rect 520792 334840 520798 334892
rect 420178 334772 420184 334824
rect 420236 334812 420242 334824
rect 444926 334812 444932 334824
rect 420236 334784 444932 334812
rect 420236 334772 420242 334784
rect 444926 334772 444932 334784
rect 444984 334772 444990 334824
rect 420270 334704 420276 334756
rect 420328 334744 420334 334756
rect 445662 334744 445668 334756
rect 420328 334716 445668 334744
rect 420328 334704 420334 334716
rect 445662 334704 445668 334716
rect 445720 334704 445726 334756
rect 513006 334704 513012 334756
rect 513064 334744 513070 334756
rect 520826 334744 520832 334756
rect 513064 334716 520832 334744
rect 513064 334704 513070 334716
rect 520826 334704 520832 334716
rect 520884 334704 520890 334756
rect 420638 334636 420644 334688
rect 420696 334676 420702 334688
rect 449526 334676 449532 334688
rect 420696 334648 449532 334676
rect 420696 334636 420702 334648
rect 449526 334636 449532 334648
rect 449584 334636 449590 334688
rect 420730 334568 420736 334620
rect 420788 334608 420794 334620
rect 449618 334608 449624 334620
rect 420788 334580 449624 334608
rect 420788 334568 420794 334580
rect 449618 334568 449624 334580
rect 449676 334568 449682 334620
rect 443638 334024 443644 334076
rect 443696 334064 443702 334076
rect 447226 334064 447232 334076
rect 443696 334036 447232 334064
rect 443696 334024 443702 334036
rect 447226 334024 447232 334036
rect 447284 334024 447290 334076
rect 364058 333956 364064 334008
rect 364116 333996 364122 334008
rect 447134 333996 447140 334008
rect 364116 333968 447140 333996
rect 364116 333956 364122 333968
rect 447134 333956 447140 333968
rect 447192 333956 447198 334008
rect 439590 332664 439596 332716
rect 439648 332704 439654 332716
rect 447226 332704 447232 332716
rect 439648 332676 447232 332704
rect 439648 332664 439654 332676
rect 447226 332664 447232 332676
rect 447284 332664 447290 332716
rect 436738 332596 436744 332648
rect 436796 332636 436802 332648
rect 447134 332636 447140 332648
rect 436796 332608 447140 332636
rect 436796 332596 436802 332608
rect 447134 332596 447140 332608
rect 447192 332596 447198 332648
rect 512638 331304 512644 331356
rect 512696 331344 512702 331356
rect 513926 331344 513932 331356
rect 512696 331316 513932 331344
rect 512696 331304 512702 331316
rect 513926 331304 513932 331316
rect 513984 331304 513990 331356
rect 447134 330488 447140 330540
rect 447192 330528 447198 330540
rect 447870 330528 447876 330540
rect 447192 330500 447876 330528
rect 447192 330488 447198 330500
rect 447870 330488 447876 330500
rect 447928 330488 447934 330540
rect 450078 330488 450084 330540
rect 450136 330528 450142 330540
rect 450722 330528 450728 330540
rect 450136 330500 450728 330528
rect 450136 330488 450142 330500
rect 450722 330488 450728 330500
rect 450780 330488 450786 330540
rect 439498 330420 439504 330472
rect 439556 330460 439562 330472
rect 447410 330460 447416 330472
rect 439556 330432 447416 330460
rect 439556 330420 439562 330432
rect 447410 330420 447416 330432
rect 447468 330460 447474 330472
rect 448054 330460 448060 330472
rect 447468 330432 448060 330460
rect 447468 330420 447474 330432
rect 448054 330420 448060 330432
rect 448112 330420 448118 330472
rect 442902 330352 442908 330404
rect 442960 330392 442966 330404
rect 447226 330392 447232 330404
rect 442960 330364 447232 330392
rect 442960 330352 442966 330364
rect 447226 330352 447232 330364
rect 447284 330352 447290 330404
rect 432782 330216 432788 330268
rect 432840 330256 432846 330268
rect 439774 330256 439780 330268
rect 432840 330228 439780 330256
rect 432840 330216 432846 330228
rect 439774 330216 439780 330228
rect 439832 330216 439838 330268
rect 512638 328584 512644 328636
rect 512696 328624 512702 328636
rect 516962 328624 516968 328636
rect 512696 328596 516968 328624
rect 512696 328584 512702 328596
rect 516962 328584 516968 328596
rect 517020 328584 517026 328636
rect 436002 328516 436008 328568
rect 436060 328556 436066 328568
rect 449894 328556 449900 328568
rect 436060 328528 449900 328556
rect 436060 328516 436066 328528
rect 449894 328516 449900 328528
rect 449952 328516 449958 328568
rect 431862 328448 431868 328500
rect 431920 328488 431926 328500
rect 450446 328488 450452 328500
rect 431920 328460 450452 328488
rect 431920 328448 431926 328460
rect 450446 328448 450452 328460
rect 450504 328448 450510 328500
rect 446306 327428 446312 327480
rect 446364 327468 446370 327480
rect 449710 327468 449716 327480
rect 446364 327440 449716 327468
rect 446364 327428 446370 327440
rect 449710 327428 449716 327440
rect 449768 327428 449774 327480
rect 509326 326408 509332 326460
rect 509384 326448 509390 326460
rect 509970 326448 509976 326460
rect 509384 326420 509976 326448
rect 509384 326408 509390 326420
rect 509970 326408 509976 326420
rect 510028 326408 510034 326460
rect 509418 326340 509424 326392
rect 509476 326380 509482 326392
rect 509694 326380 509700 326392
rect 509476 326352 509700 326380
rect 509476 326340 509482 326352
rect 509694 326340 509700 326352
rect 509752 326340 509758 326392
rect 437014 324980 437020 325032
rect 437072 325020 437078 325032
rect 439314 325020 439320 325032
rect 437072 324992 439320 325020
rect 437072 324980 437078 324992
rect 439314 324980 439320 324992
rect 439372 324980 439378 325032
rect 432874 324912 432880 324964
rect 432932 324952 432938 324964
rect 442258 324952 442264 324964
rect 432932 324924 442264 324952
rect 432932 324912 432938 324924
rect 442258 324912 442264 324924
rect 442316 324912 442322 324964
rect 510430 324912 510436 324964
rect 510488 324952 510494 324964
rect 580626 324952 580632 324964
rect 510488 324924 580632 324952
rect 510488 324912 510494 324924
rect 580626 324912 580632 324924
rect 580684 324912 580690 324964
rect 511902 323620 511908 323672
rect 511960 323660 511966 323672
rect 580166 323660 580172 323672
rect 511960 323632 580172 323660
rect 511960 323620 511966 323632
rect 580166 323620 580172 323632
rect 580224 323620 580230 323672
rect 510522 323552 510528 323604
rect 510580 323592 510586 323604
rect 580534 323592 580540 323604
rect 510580 323564 580540 323592
rect 510580 323552 510586 323564
rect 580534 323552 580540 323564
rect 580592 323552 580598 323604
rect 459940 323088 463694 323116
rect 432598 322940 432604 322992
rect 432656 322980 432662 322992
rect 436922 322980 436928 322992
rect 432656 322952 436928 322980
rect 432656 322940 432662 322952
rect 436922 322940 436928 322952
rect 436980 322940 436986 322992
rect 445570 322736 445576 322788
rect 445628 322776 445634 322788
rect 445628 322748 451274 322776
rect 445628 322736 445634 322748
rect 451246 322640 451274 322748
rect 459646 322668 459652 322720
rect 459704 322708 459710 322720
rect 459940 322708 459968 323088
rect 461320 323020 462820 323048
rect 461320 322720 461348 323020
rect 462792 322844 462820 323020
rect 463666 322912 463694 323088
rect 473326 323020 473860 323048
rect 473326 322912 473354 323020
rect 473832 322912 473860 323020
rect 570598 322912 570604 322924
rect 463666 322884 473354 322912
rect 473464 322884 473768 322912
rect 473832 322884 570604 322912
rect 473464 322844 473492 322884
rect 462792 322816 473492 322844
rect 473740 322844 473768 322884
rect 570598 322872 570604 322884
rect 570656 322872 570662 322924
rect 569218 322844 569224 322856
rect 473740 322816 569224 322844
rect 569218 322804 569224 322816
rect 569276 322804 569282 322856
rect 473308 322776 473314 322788
rect 462700 322748 473314 322776
rect 459704 322680 459968 322708
rect 459704 322668 459710 322680
rect 461302 322668 461308 322720
rect 461360 322668 461366 322720
rect 462700 322640 462728 322748
rect 473308 322736 473314 322748
rect 473366 322736 473372 322788
rect 571978 322776 571984 322788
rect 480640 322748 571984 322776
rect 480640 322720 480668 322748
rect 571978 322736 571984 322748
rect 572036 322736 572042 322788
rect 473446 322708 473452 322720
rect 451246 322612 462728 322640
rect 462884 322680 473452 322708
rect 459094 322532 459100 322584
rect 459152 322572 459158 322584
rect 462884 322572 462912 322680
rect 473446 322668 473452 322680
rect 473504 322668 473510 322720
rect 480622 322668 480628 322720
rect 480680 322668 480686 322720
rect 519630 322708 519636 322720
rect 482986 322680 519636 322708
rect 462958 322600 462964 322652
rect 463016 322640 463022 322652
rect 478138 322640 478144 322652
rect 463016 322612 478144 322640
rect 463016 322600 463022 322612
rect 478138 322600 478144 322612
rect 478196 322600 478202 322652
rect 480898 322600 480904 322652
rect 480956 322640 480962 322652
rect 482986 322640 483014 322680
rect 519630 322668 519636 322680
rect 519688 322668 519694 322720
rect 515398 322640 515404 322652
rect 480956 322612 483014 322640
rect 485746 322612 515404 322640
rect 480956 322600 480962 322612
rect 459152 322544 462912 322572
rect 459152 322532 459158 322544
rect 469030 322532 469036 322584
rect 469088 322572 469094 322584
rect 469088 322544 473124 322572
rect 469088 322532 469094 322544
rect 445018 322464 445024 322516
rect 445076 322504 445082 322516
rect 473096 322504 473124 322544
rect 473464 322544 474044 322572
rect 473464 322504 473492 322544
rect 445076 322476 471284 322504
rect 473096 322476 473492 322504
rect 474016 322504 474044 322544
rect 480622 322532 480628 322584
rect 480680 322572 480686 322584
rect 485746 322572 485774 322612
rect 515398 322600 515404 322612
rect 515456 322600 515462 322652
rect 515490 322572 515496 322584
rect 480680 322544 485774 322572
rect 495406 322544 515496 322572
rect 480680 322532 480686 322544
rect 495406 322504 495434 322544
rect 515490 322532 515496 322544
rect 515548 322532 515554 322584
rect 474016 322476 495434 322504
rect 445076 322464 445082 322476
rect 446582 322396 446588 322448
rect 446640 322436 446646 322448
rect 471256 322436 471284 322476
rect 507394 322464 507400 322516
rect 507452 322504 507458 322516
rect 509878 322504 509884 322516
rect 507452 322476 509884 322504
rect 507452 322464 507458 322476
rect 509878 322464 509884 322476
rect 509936 322464 509942 322516
rect 473446 322436 473452 322448
rect 446640 322408 471192 322436
rect 471256 322408 473452 322436
rect 446640 322396 446646 322408
rect 439866 322328 439872 322380
rect 439924 322368 439930 322380
rect 471164 322368 471192 322408
rect 473446 322396 473452 322408
rect 473504 322396 473510 322448
rect 482278 322368 482284 322380
rect 439924 322340 466454 322368
rect 471164 322340 482284 322368
rect 439924 322328 439930 322340
rect 442350 322260 442356 322312
rect 442408 322300 442414 322312
rect 463786 322300 463792 322312
rect 442408 322272 463792 322300
rect 442408 322260 442414 322272
rect 463786 322260 463792 322272
rect 463844 322260 463850 322312
rect 466426 322300 466454 322340
rect 482278 322328 482284 322340
rect 482336 322328 482342 322380
rect 473446 322300 473452 322312
rect 466426 322272 473452 322300
rect 473446 322260 473452 322272
rect 473504 322260 473510 322312
rect 478138 322260 478144 322312
rect 478196 322300 478202 322312
rect 480622 322300 480628 322312
rect 478196 322272 480628 322300
rect 478196 322260 478202 322272
rect 480622 322260 480628 322272
rect 480680 322260 480686 322312
rect 506934 322260 506940 322312
rect 506992 322300 506998 322312
rect 511442 322300 511448 322312
rect 506992 322272 511448 322300
rect 506992 322260 506998 322272
rect 511442 322260 511448 322272
rect 511500 322260 511506 322312
rect 439314 322192 439320 322244
rect 439372 322232 439378 322244
rect 474274 322232 474280 322244
rect 439372 322204 474280 322232
rect 439372 322192 439378 322204
rect 474274 322192 474280 322204
rect 474332 322192 474338 322244
rect 475102 322192 475108 322244
rect 475160 322232 475166 322244
rect 475378 322232 475384 322244
rect 475160 322204 475384 322232
rect 475160 322192 475166 322204
rect 475378 322192 475384 322204
rect 475436 322192 475442 322244
rect 490282 322192 490288 322244
rect 490340 322232 490346 322244
rect 490558 322232 490564 322244
rect 490340 322204 490564 322232
rect 490340 322192 490346 322204
rect 490558 322192 490564 322204
rect 490616 322192 490622 322244
rect 442442 322124 442448 322176
rect 442500 322164 442506 322176
rect 484210 322164 484216 322176
rect 442500 322136 473354 322164
rect 442500 322124 442506 322136
rect 459370 322056 459376 322108
rect 459428 322096 459434 322108
rect 462958 322096 462964 322108
rect 459428 322068 462964 322096
rect 459428 322056 459434 322068
rect 462958 322056 462964 322068
rect 463016 322056 463022 322108
rect 473326 322028 473354 322136
rect 482986 322136 484216 322164
rect 482986 322028 483014 322136
rect 484210 322124 484216 322136
rect 484268 322124 484274 322176
rect 473326 322000 483014 322028
rect 509418 321988 509424 322040
rect 509476 322028 509482 322040
rect 509970 322028 509976 322040
rect 509476 322000 509976 322028
rect 509476 321988 509482 322000
rect 509970 321988 509976 322000
rect 510028 321988 510034 322040
rect 507486 321784 507492 321836
rect 507544 321824 507550 321836
rect 511166 321824 511172 321836
rect 507544 321796 511172 321824
rect 507544 321784 507550 321796
rect 511166 321784 511172 321796
rect 511224 321784 511230 321836
rect 458082 321512 458088 321564
rect 458140 321552 458146 321564
rect 580810 321552 580816 321564
rect 458140 321524 580816 321552
rect 458140 321512 458146 321524
rect 580810 321512 580816 321524
rect 580868 321512 580874 321564
rect 458358 321444 458364 321496
rect 458416 321484 458422 321496
rect 580718 321484 580724 321496
rect 458416 321456 580724 321484
rect 458416 321444 458422 321456
rect 580718 321444 580724 321456
rect 580776 321444 580782 321496
rect 446490 321376 446496 321428
rect 446548 321416 446554 321428
rect 460842 321416 460848 321428
rect 446548 321388 460848 321416
rect 446548 321376 446554 321388
rect 460842 321376 460848 321388
rect 460900 321376 460906 321428
rect 468570 321376 468576 321428
rect 468628 321416 468634 321428
rect 576210 321416 576216 321428
rect 468628 321388 576216 321416
rect 468628 321376 468634 321388
rect 576210 321376 576216 321388
rect 576268 321376 576274 321428
rect 449158 321308 449164 321360
rect 449216 321348 449222 321360
rect 461670 321348 461676 321360
rect 449216 321320 461676 321348
rect 449216 321308 449222 321320
rect 461670 321308 461676 321320
rect 461728 321308 461734 321360
rect 469950 321308 469956 321360
rect 470008 321348 470014 321360
rect 574738 321348 574744 321360
rect 470008 321320 574744 321348
rect 470008 321308 470014 321320
rect 574738 321308 574744 321320
rect 574796 321308 574802 321360
rect 479334 321240 479340 321292
rect 479392 321280 479398 321292
rect 573358 321280 573364 321292
rect 479392 321252 573364 321280
rect 479392 321240 479398 321252
rect 573358 321240 573364 321252
rect 573416 321240 573422 321292
rect 444926 321172 444932 321224
rect 444984 321212 444990 321224
rect 484578 321212 484584 321224
rect 444984 321184 484584 321212
rect 444984 321172 444990 321184
rect 484578 321172 484584 321184
rect 484636 321172 484642 321224
rect 507670 321172 507676 321224
rect 507728 321212 507734 321224
rect 509970 321212 509976 321224
rect 507728 321184 509976 321212
rect 507728 321172 507734 321184
rect 509970 321172 509976 321184
rect 510028 321172 510034 321224
rect 447502 321104 447508 321156
rect 447560 321144 447566 321156
rect 463326 321144 463332 321156
rect 447560 321116 463332 321144
rect 447560 321104 447566 321116
rect 463326 321104 463332 321116
rect 463384 321104 463390 321156
rect 479058 321104 479064 321156
rect 479116 321144 479122 321156
rect 514018 321144 514024 321156
rect 479116 321116 514024 321144
rect 479116 321104 479122 321116
rect 514018 321104 514024 321116
rect 514076 321104 514082 321156
rect 447042 321036 447048 321088
rect 447100 321076 447106 321088
rect 484026 321076 484032 321088
rect 447100 321048 484032 321076
rect 447100 321036 447106 321048
rect 484026 321036 484032 321048
rect 484084 321036 484090 321088
rect 507302 321036 507308 321088
rect 507360 321076 507366 321088
rect 517514 321076 517520 321088
rect 507360 321048 517520 321076
rect 507360 321036 507366 321048
rect 517514 321036 517520 321048
rect 517572 321036 517578 321088
rect 460658 320968 460664 321020
rect 460716 321008 460722 321020
rect 516134 321008 516140 321020
rect 460716 320980 516140 321008
rect 460716 320968 460722 320980
rect 516134 320968 516140 320980
rect 516192 320968 516198 321020
rect 441154 320900 441160 320952
rect 441212 320940 441218 320952
rect 471882 320940 471888 320952
rect 441212 320912 471888 320940
rect 441212 320900 441218 320912
rect 471882 320900 471888 320912
rect 471940 320900 471946 320952
rect 502242 320900 502248 320952
rect 502300 320940 502306 320952
rect 580258 320940 580264 320952
rect 502300 320912 580264 320940
rect 502300 320900 502306 320912
rect 580258 320900 580264 320912
rect 580316 320900 580322 320952
rect 446398 320832 446404 320884
rect 446456 320872 446462 320884
rect 451826 320872 451832 320884
rect 446456 320844 451832 320872
rect 446456 320832 446462 320844
rect 451826 320832 451832 320844
rect 451884 320832 451890 320884
rect 451936 320844 456794 320872
rect 444098 320764 444104 320816
rect 444156 320804 444162 320816
rect 451936 320804 451964 320844
rect 444156 320776 451964 320804
rect 456766 320804 456794 320844
rect 459922 320832 459928 320884
rect 459980 320872 459986 320884
rect 580350 320872 580356 320884
rect 459980 320844 580356 320872
rect 459980 320832 459986 320844
rect 580350 320832 580356 320844
rect 580408 320832 580414 320884
rect 481818 320804 481824 320816
rect 456766 320776 481824 320804
rect 444156 320764 444162 320776
rect 481818 320764 481824 320776
rect 481876 320764 481882 320816
rect 507578 320764 507584 320816
rect 507636 320804 507642 320816
rect 507636 320776 511304 320804
rect 507636 320764 507642 320776
rect 451918 320696 451924 320748
rect 451976 320736 451982 320748
rect 461394 320736 461400 320748
rect 451976 320708 461400 320736
rect 451976 320696 451982 320708
rect 461394 320696 461400 320708
rect 461452 320696 461458 320748
rect 507118 320696 507124 320748
rect 507176 320736 507182 320748
rect 511276 320736 511304 320776
rect 512638 320764 512644 320816
rect 512696 320804 512702 320816
rect 512822 320804 512828 320816
rect 512696 320776 512828 320804
rect 512696 320764 512702 320776
rect 512822 320764 512828 320776
rect 512880 320764 512886 320816
rect 513374 320736 513380 320748
rect 507176 320708 509234 320736
rect 511276 320708 513380 320736
rect 507176 320696 507182 320708
rect 441062 320628 441068 320680
rect 441120 320668 441126 320680
rect 472434 320668 472440 320680
rect 441120 320640 448744 320668
rect 441120 320628 441126 320640
rect 446858 320560 446864 320612
rect 446916 320600 446922 320612
rect 447502 320600 447508 320612
rect 446916 320572 447508 320600
rect 446916 320560 446922 320572
rect 447502 320560 447508 320572
rect 447560 320560 447566 320612
rect 448716 320600 448744 320640
rect 448900 320640 472440 320668
rect 448900 320600 448928 320640
rect 472434 320628 472440 320640
rect 472492 320628 472498 320680
rect 509206 320668 509234 320708
rect 513374 320696 513380 320708
rect 513432 320696 513438 320748
rect 513466 320668 513472 320680
rect 509206 320640 513472 320668
rect 513466 320628 513472 320640
rect 513524 320628 513530 320680
rect 448716 320572 448928 320600
rect 449710 320560 449716 320612
rect 449768 320600 449774 320612
rect 463050 320600 463056 320612
rect 449768 320572 463056 320600
rect 449768 320560 449774 320572
rect 463050 320560 463056 320572
rect 463108 320560 463114 320612
rect 441246 320492 441252 320544
rect 441304 320532 441310 320544
rect 482094 320532 482100 320544
rect 441304 320504 482100 320532
rect 441304 320492 441310 320504
rect 482094 320492 482100 320504
rect 482152 320492 482158 320544
rect 441522 320424 441528 320476
rect 441580 320464 441586 320476
rect 481266 320464 481272 320476
rect 441580 320436 481272 320464
rect 441580 320424 441586 320436
rect 481266 320424 481272 320436
rect 481324 320424 481330 320476
rect 507762 320220 507768 320272
rect 507820 320260 507826 320272
rect 511074 320260 511080 320272
rect 507820 320232 511080 320260
rect 507820 320220 507826 320232
rect 511074 320220 511080 320232
rect 511132 320220 511138 320272
rect 479886 320084 479892 320136
rect 479944 320124 479950 320136
rect 580442 320124 580448 320136
rect 479944 320096 580448 320124
rect 479944 320084 479950 320096
rect 580442 320084 580448 320096
rect 580500 320084 580506 320136
rect 442718 320016 442724 320068
rect 442776 320056 442782 320068
rect 460566 320056 460572 320068
rect 442776 320028 460572 320056
rect 442776 320016 442782 320028
rect 460566 320016 460572 320028
rect 460624 320016 460630 320068
rect 480714 320016 480720 320068
rect 480772 320056 480778 320068
rect 576118 320056 576124 320068
rect 480772 320028 576124 320056
rect 480772 320016 480778 320028
rect 576118 320016 576124 320028
rect 576176 320016 576182 320068
rect 444282 319948 444288 320000
rect 444340 319988 444346 320000
rect 460290 319988 460296 320000
rect 444340 319960 460296 319988
rect 444340 319948 444346 319960
rect 460290 319948 460296 319960
rect 460348 319948 460354 320000
rect 469674 319948 469680 320000
rect 469732 319988 469738 320000
rect 511258 319988 511264 320000
rect 469732 319960 511264 319988
rect 469732 319948 469738 319960
rect 511258 319948 511264 319960
rect 511316 319948 511322 320000
rect 449618 319880 449624 319932
rect 449676 319920 449682 319932
rect 463602 319920 463608 319932
rect 449676 319892 463608 319920
rect 449676 319880 449682 319892
rect 463602 319880 463608 319892
rect 463660 319880 463666 319932
rect 468846 319880 468852 319932
rect 468904 319920 468910 319932
rect 510430 319920 510436 319932
rect 468904 319892 510436 319920
rect 468904 319880 468910 319892
rect 510430 319880 510436 319892
rect 510488 319880 510494 319932
rect 449250 319812 449256 319864
rect 449308 319852 449314 319864
rect 461118 319852 461124 319864
rect 449308 319824 461124 319852
rect 449308 319812 449314 319824
rect 461118 319812 461124 319824
rect 461176 319812 461182 319864
rect 469398 319812 469404 319864
rect 469456 319852 469462 319864
rect 510522 319852 510528 319864
rect 469456 319824 510528 319852
rect 469456 319812 469462 319824
rect 510522 319812 510528 319824
rect 510580 319812 510586 319864
rect 449434 319744 449440 319796
rect 449492 319784 449498 319796
rect 471054 319784 471060 319796
rect 449492 319756 471060 319784
rect 449492 319744 449498 319756
rect 471054 319744 471060 319756
rect 471112 319744 471118 319796
rect 480162 319744 480168 319796
rect 480220 319784 480226 319796
rect 519538 319784 519544 319796
rect 480220 319756 519544 319784
rect 480220 319744 480226 319756
rect 519538 319744 519544 319756
rect 519596 319744 519602 319796
rect 445110 319676 445116 319728
rect 445168 319716 445174 319728
rect 471330 319716 471336 319728
rect 445168 319688 471336 319716
rect 445168 319676 445174 319688
rect 471330 319676 471336 319688
rect 471388 319676 471394 319728
rect 479610 319676 479616 319728
rect 479668 319716 479674 319728
rect 518158 319716 518164 319728
rect 479668 319688 518164 319716
rect 479668 319676 479674 319688
rect 518158 319676 518164 319688
rect 518216 319676 518222 319728
rect 449526 319608 449532 319660
rect 449584 319648 449590 319660
rect 474090 319648 474096 319660
rect 449584 319620 474096 319648
rect 449584 319608 449590 319620
rect 474090 319608 474096 319620
rect 474148 319608 474154 319660
rect 478782 319608 478788 319660
rect 478840 319648 478846 319660
rect 511902 319648 511908 319660
rect 478840 319620 511908 319648
rect 478840 319608 478846 319620
rect 511902 319608 511908 319620
rect 511960 319608 511966 319660
rect 445478 319540 445484 319592
rect 445536 319580 445542 319592
rect 462774 319580 462780 319592
rect 445536 319552 462780 319580
rect 445536 319540 445542 319552
rect 462774 319540 462780 319552
rect 462832 319540 462838 319592
rect 470226 319540 470232 319592
rect 470284 319580 470290 319592
rect 502242 319580 502248 319592
rect 470284 319552 502248 319580
rect 470284 319540 470290 319552
rect 502242 319540 502248 319552
rect 502300 319540 502306 319592
rect 502794 319540 502800 319592
rect 502852 319580 502858 319592
rect 533338 319580 533344 319592
rect 502852 319552 533344 319580
rect 502852 319540 502858 319552
rect 533338 319540 533344 319552
rect 533396 319540 533402 319592
rect 445386 319472 445392 319524
rect 445444 319512 445450 319524
rect 483474 319512 483480 319524
rect 445444 319484 483480 319512
rect 445444 319472 445450 319484
rect 483474 319472 483480 319484
rect 483532 319472 483538 319524
rect 498654 319472 498660 319524
rect 498712 319512 498718 319524
rect 534718 319512 534724 319524
rect 498712 319484 534724 319512
rect 498712 319472 498718 319484
rect 534718 319472 534724 319484
rect 534776 319472 534782 319524
rect 460290 319404 460296 319456
rect 460348 319444 460354 319456
rect 476298 319444 476304 319456
rect 460348 319416 476304 319444
rect 460348 319404 460354 319416
rect 476298 319404 476304 319416
rect 476356 319404 476362 319456
rect 502150 319404 502156 319456
rect 502208 319444 502214 319456
rect 538858 319444 538864 319456
rect 502208 319416 538864 319444
rect 502208 319404 502214 319416
rect 538858 319404 538864 319416
rect 538916 319404 538922 319456
rect 440970 319336 440976 319388
rect 441028 319376 441034 319388
rect 472158 319376 472164 319388
rect 441028 319348 472164 319376
rect 441028 319336 441034 319348
rect 472158 319336 472164 319348
rect 472216 319336 472222 319388
rect 445662 319268 445668 319320
rect 445720 319308 445726 319320
rect 473814 319308 473820 319320
rect 445720 319280 473820 319308
rect 445720 319268 445726 319280
rect 473814 319268 473820 319280
rect 473872 319268 473878 319320
rect 445294 319200 445300 319252
rect 445352 319240 445358 319252
rect 482922 319240 482928 319252
rect 445352 319212 482928 319240
rect 445352 319200 445358 319212
rect 482922 319200 482928 319212
rect 482980 319200 482986 319252
rect 487246 319200 487252 319252
rect 487304 319240 487310 319252
rect 488350 319240 488356 319252
rect 487304 319212 488356 319240
rect 487304 319200 487310 319212
rect 488350 319200 488356 319212
rect 488408 319200 488414 319252
rect 442810 319132 442816 319184
rect 442868 319172 442874 319184
rect 470778 319172 470784 319184
rect 442868 319144 470784 319172
rect 442868 319132 442874 319144
rect 470778 319132 470784 319144
rect 470836 319132 470842 319184
rect 483658 319132 483664 319184
rect 483716 319172 483722 319184
rect 484854 319172 484860 319184
rect 483716 319144 484860 319172
rect 483716 319132 483722 319144
rect 484854 319132 484860 319144
rect 484912 319132 484918 319184
rect 494146 319132 494152 319184
rect 494204 319172 494210 319184
rect 494422 319172 494428 319184
rect 494204 319144 494428 319172
rect 494204 319132 494210 319144
rect 494422 319132 494428 319144
rect 494480 319132 494486 319184
rect 509418 319132 509424 319184
rect 509476 319172 509482 319184
rect 509694 319172 509700 319184
rect 509476 319144 509700 319172
rect 509476 319132 509482 319144
rect 509694 319132 509700 319144
rect 509752 319132 509758 319184
rect 446950 319064 446956 319116
rect 447008 319104 447014 319116
rect 483750 319104 483756 319116
rect 447008 319076 483756 319104
rect 447008 319064 447014 319076
rect 483750 319064 483756 319076
rect 483808 319064 483814 319116
rect 484762 319064 484768 319116
rect 484820 319104 484826 319116
rect 485590 319104 485596 319116
rect 484820 319076 485596 319104
rect 484820 319064 484826 319076
rect 485590 319064 485596 319076
rect 485648 319064 485654 319116
rect 485866 319064 485872 319116
rect 485924 319104 485930 319116
rect 486970 319104 486976 319116
rect 485924 319076 486976 319104
rect 485924 319064 485930 319076
rect 486970 319064 486976 319076
rect 487028 319064 487034 319116
rect 487798 319064 487804 319116
rect 487856 319104 487862 319116
rect 488350 319104 488356 319116
rect 487856 319076 488356 319104
rect 487856 319064 487862 319076
rect 488350 319064 488356 319076
rect 488408 319064 488414 319116
rect 488902 319064 488908 319116
rect 488960 319104 488966 319116
rect 489454 319104 489460 319116
rect 488960 319076 489460 319104
rect 488960 319064 488966 319076
rect 489454 319064 489460 319076
rect 489512 319064 489518 319116
rect 491662 319064 491668 319116
rect 491720 319104 491726 319116
rect 492214 319104 492220 319116
rect 491720 319076 492220 319104
rect 491720 319064 491726 319076
rect 492214 319064 492220 319076
rect 492272 319064 492278 319116
rect 493318 319064 493324 319116
rect 493376 319104 493382 319116
rect 493870 319104 493876 319116
rect 493376 319076 493876 319104
rect 493376 319064 493382 319076
rect 493870 319064 493876 319076
rect 493928 319064 493934 319116
rect 494698 319064 494704 319116
rect 494756 319104 494762 319116
rect 495250 319104 495256 319116
rect 494756 319076 495256 319104
rect 494756 319064 494762 319076
rect 495250 319064 495256 319076
rect 495308 319064 495314 319116
rect 499942 319064 499948 319116
rect 500000 319104 500006 319116
rect 500218 319104 500224 319116
rect 500000 319076 500224 319104
rect 500000 319064 500006 319076
rect 500218 319064 500224 319076
rect 500276 319064 500282 319116
rect 501322 319064 501328 319116
rect 501380 319104 501386 319116
rect 501874 319104 501880 319116
rect 501380 319076 501880 319104
rect 501380 319064 501386 319076
rect 501874 319064 501880 319076
rect 501932 319064 501938 319116
rect 464062 318996 464068 319048
rect 464120 319036 464126 319048
rect 464614 319036 464620 319048
rect 464120 319008 464620 319036
rect 464120 318996 464126 319008
rect 464614 318996 464620 319008
rect 464672 318996 464678 319048
rect 465166 318996 465172 319048
rect 465224 319036 465230 319048
rect 465718 319036 465724 319048
rect 465224 319008 465724 319036
rect 465224 318996 465230 319008
rect 465718 318996 465724 319008
rect 465776 318996 465782 319048
rect 466822 318996 466828 319048
rect 466880 319036 466886 319048
rect 467374 319036 467380 319048
rect 466880 319008 467380 319036
rect 466880 318996 466886 319008
rect 467374 318996 467380 319008
rect 467432 318996 467438 319048
rect 475102 318996 475108 319048
rect 475160 319036 475166 319048
rect 475654 319036 475660 319048
rect 475160 319008 475660 319036
rect 475160 318996 475166 319008
rect 475654 318996 475660 319008
rect 475712 318996 475718 319048
rect 484486 318996 484492 319048
rect 484544 319036 484550 319048
rect 485314 319036 485320 319048
rect 484544 319008 485320 319036
rect 484544 318996 484550 319008
rect 485314 318996 485320 319008
rect 485372 318996 485378 319048
rect 488626 318996 488632 319048
rect 488684 319036 488690 319048
rect 489178 319036 489184 319048
rect 488684 319008 489184 319036
rect 488684 318996 488690 319008
rect 489178 318996 489184 319008
rect 489236 318996 489242 319048
rect 491386 318996 491392 319048
rect 491444 319036 491450 319048
rect 492490 319036 492496 319048
rect 491444 319008 492496 319036
rect 491444 318996 491450 319008
rect 492490 318996 492496 319008
rect 492548 318996 492554 319048
rect 493042 318996 493048 319048
rect 493100 319036 493106 319048
rect 493594 319036 493600 319048
rect 493100 319008 493600 319036
rect 493100 318996 493106 319008
rect 493594 318996 493600 319008
rect 493652 318996 493658 319048
rect 463786 318928 463792 318980
rect 463844 318968 463850 318980
rect 464890 318968 464896 318980
rect 463844 318940 464896 318968
rect 463844 318928 463850 318940
rect 464890 318928 464896 318940
rect 464948 318928 464954 318980
rect 467098 318928 467104 318980
rect 467156 318968 467162 318980
rect 467650 318968 467656 318980
rect 467156 318940 467656 318968
rect 467156 318928 467162 318940
rect 467650 318928 467656 318940
rect 467708 318928 467714 318980
rect 490282 318860 490288 318912
rect 490340 318900 490346 318912
rect 491110 318900 491116 318912
rect 490340 318872 491116 318900
rect 490340 318860 490346 318872
rect 491110 318860 491116 318872
rect 491168 318860 491174 318912
rect 432046 318248 432052 318300
rect 432104 318288 432110 318300
rect 435450 318288 435456 318300
rect 432104 318260 435456 318288
rect 432104 318248 432110 318260
rect 435450 318248 435456 318260
rect 435508 318248 435514 318300
rect 454678 318180 454684 318232
rect 454736 318220 454742 318232
rect 488718 318220 488724 318232
rect 454736 318192 488724 318220
rect 454736 318180 454742 318192
rect 488718 318180 488724 318192
rect 488776 318180 488782 318232
rect 451918 318112 451924 318164
rect 451976 318152 451982 318164
rect 495618 318152 495624 318164
rect 451976 318124 495624 318152
rect 451976 318112 451982 318124
rect 495618 318112 495624 318124
rect 495676 318112 495682 318164
rect 496170 318112 496176 318164
rect 496228 318152 496234 318164
rect 540974 318152 540980 318164
rect 496228 318124 540980 318152
rect 496228 318112 496234 318124
rect 540974 318112 540980 318124
rect 541032 318112 541038 318164
rect 477678 318044 477684 318096
rect 477736 318084 477742 318096
rect 547138 318084 547144 318096
rect 477736 318056 547144 318084
rect 477736 318044 477742 318056
rect 547138 318044 547144 318056
rect 547196 318044 547202 318096
rect 478506 317364 478512 317416
rect 478564 317404 478570 317416
rect 479518 317404 479524 317416
rect 478564 317376 479524 317404
rect 478564 317364 478570 317376
rect 479518 317364 479524 317376
rect 479576 317364 479582 317416
rect 457806 317024 457812 317076
rect 457864 317064 457870 317076
rect 461578 317064 461584 317076
rect 457864 317036 461584 317064
rect 457864 317024 457870 317036
rect 461578 317024 461584 317036
rect 461636 317024 461642 317076
rect 501414 316888 501420 316940
rect 501472 316928 501478 316940
rect 539686 316928 539692 316940
rect 501472 316900 539692 316928
rect 501472 316888 501478 316900
rect 539686 316888 539692 316900
rect 539744 316888 539750 316940
rect 500310 316820 500316 316872
rect 500368 316860 500374 316872
rect 539594 316860 539600 316872
rect 500368 316832 539600 316860
rect 500368 316820 500374 316832
rect 539594 316820 539600 316832
rect 539652 316820 539658 316872
rect 487338 316752 487344 316804
rect 487396 316792 487402 316804
rect 529934 316792 529940 316804
rect 487396 316764 529940 316792
rect 487396 316752 487402 316764
rect 529934 316752 529940 316764
rect 529992 316752 529998 316804
rect 458910 316684 458916 316736
rect 458968 316724 458974 316736
rect 491478 316724 491484 316736
rect 458968 316696 491484 316724
rect 458968 316684 458974 316696
rect 491478 316684 491484 316696
rect 491536 316684 491542 316736
rect 496998 316684 497004 316736
rect 497056 316724 497062 316736
rect 542998 316724 543004 316736
rect 497056 316696 543004 316724
rect 497056 316684 497062 316696
rect 542998 316684 543004 316696
rect 543056 316684 543062 316736
rect 457438 316072 457444 316124
rect 457496 316112 457502 316124
rect 457990 316112 457996 316124
rect 457496 316084 457996 316112
rect 457496 316072 457502 316084
rect 457990 316072 457996 316084
rect 458048 316072 458054 316124
rect 465442 316072 465448 316124
rect 465500 316112 465506 316124
rect 465994 316112 466000 316124
rect 465500 316084 466000 316112
rect 465500 316072 465506 316084
rect 465994 316072 466000 316084
rect 466052 316072 466058 316124
rect 486326 316004 486332 316056
rect 486384 316044 486390 316056
rect 486510 316044 486516 316056
rect 486384 316016 486516 316044
rect 486384 316004 486390 316016
rect 486510 316004 486516 316016
rect 486568 316004 486574 316056
rect 361758 315936 361764 315988
rect 361816 315976 361822 315988
rect 371878 315976 371884 315988
rect 361816 315948 371884 315976
rect 361816 315936 361822 315948
rect 371878 315936 371884 315948
rect 371936 315936 371942 315988
rect 501874 315392 501880 315444
rect 501932 315432 501938 315444
rect 539778 315432 539784 315444
rect 501932 315404 539784 315432
rect 501932 315392 501938 315404
rect 539778 315392 539784 315404
rect 539836 315392 539842 315444
rect 457438 315324 457444 315376
rect 457496 315364 457502 315376
rect 491754 315364 491760 315376
rect 457496 315336 491760 315364
rect 457496 315324 457502 315336
rect 491754 315324 491760 315336
rect 491812 315324 491818 315376
rect 502978 315324 502984 315376
rect 503036 315364 503042 315376
rect 542722 315364 542728 315376
rect 503036 315336 542728 315364
rect 503036 315324 503042 315336
rect 542722 315324 542728 315336
rect 542780 315324 542786 315376
rect 455874 315256 455880 315308
rect 455932 315296 455938 315308
rect 562318 315296 562324 315308
rect 455932 315268 562324 315296
rect 455932 315256 455938 315268
rect 562318 315256 562324 315268
rect 562376 315256 562382 315308
rect 454770 313964 454776 314016
rect 454828 314004 454834 314016
rect 491938 314004 491944 314016
rect 454828 313976 491944 314004
rect 454828 313964 454834 313976
rect 491938 313964 491944 313976
rect 491996 313964 492002 314016
rect 497458 313964 497464 314016
rect 497516 314004 497522 314016
rect 542446 314004 542452 314016
rect 497516 313976 542452 314004
rect 497516 313964 497522 313976
rect 542446 313964 542452 313976
rect 542504 313964 542510 314016
rect 432690 313896 432696 313948
rect 432748 313936 432754 313948
rect 443822 313936 443828 313948
rect 432748 313908 443828 313936
rect 432748 313896 432754 313908
rect 443822 313896 443828 313908
rect 443880 313896 443886 313948
rect 477034 313896 477040 313948
rect 477092 313936 477098 313948
rect 566458 313936 566464 313948
rect 477092 313908 566464 313936
rect 477092 313896 477098 313908
rect 566458 313896 566464 313908
rect 566516 313896 566522 313948
rect 482646 313284 482652 313336
rect 482704 313324 482710 313336
rect 485038 313324 485044 313336
rect 482704 313296 485044 313324
rect 482704 313284 482710 313296
rect 485038 313284 485044 313296
rect 485096 313284 485102 313336
rect 469030 313216 469036 313268
rect 469088 313256 469094 313268
rect 580166 313256 580172 313268
rect 469088 313228 580172 313256
rect 469088 313216 469094 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 467374 312536 467380 312588
rect 467432 312576 467438 312588
rect 551278 312576 551284 312588
rect 467432 312548 551284 312576
rect 467432 312536 467438 312548
rect 551278 312536 551284 312548
rect 551336 312536 551342 312588
rect 459002 311176 459008 311228
rect 459060 311216 459066 311228
rect 493042 311216 493048 311228
rect 459060 311188 493048 311216
rect 459060 311176 459066 311188
rect 493042 311176 493048 311188
rect 493100 311176 493106 311228
rect 503530 311176 503536 311228
rect 503588 311216 503594 311228
rect 538950 311216 538956 311228
rect 503588 311188 538956 311216
rect 503588 311176 503594 311188
rect 538950 311176 538956 311188
rect 539008 311176 539014 311228
rect 462958 311108 462964 311160
rect 463016 311148 463022 311160
rect 464338 311148 464344 311160
rect 463016 311120 464344 311148
rect 463016 311108 463022 311120
rect 464338 311108 464344 311120
rect 464396 311108 464402 311160
rect 478138 311108 478144 311160
rect 478196 311148 478202 311160
rect 548518 311148 548524 311160
rect 478196 311120 548524 311148
rect 478196 311108 478202 311120
rect 548518 311108 548524 311120
rect 548576 311108 548582 311160
rect 482462 310496 482468 310548
rect 482520 310536 482526 310548
rect 483658 310536 483664 310548
rect 482520 310508 483664 310536
rect 482520 310496 482526 310508
rect 483658 310496 483664 310508
rect 483716 310496 483722 310548
rect 461670 310292 461676 310344
rect 461728 310332 461734 310344
rect 464154 310332 464160 310344
rect 461728 310304 464160 310332
rect 461728 310292 461734 310304
rect 464154 310292 464160 310304
rect 464212 310292 464218 310344
rect 454954 309816 454960 309868
rect 455012 309856 455018 309868
rect 494422 309856 494428 309868
rect 455012 309828 494428 309856
rect 455012 309816 455018 309828
rect 494422 309816 494428 309828
rect 494480 309816 494486 309868
rect 497642 309816 497648 309868
rect 497700 309856 497706 309868
rect 542538 309856 542544 309868
rect 497700 309828 542544 309856
rect 497700 309816 497706 309828
rect 542538 309816 542544 309828
rect 542596 309816 542602 309868
rect 447962 309748 447968 309800
rect 448020 309788 448026 309800
rect 533430 309788 533436 309800
rect 448020 309760 533436 309788
rect 448020 309748 448026 309760
rect 533430 309748 533436 309760
rect 533488 309748 533494 309800
rect 452010 308456 452016 308508
rect 452068 308496 452074 308508
rect 494790 308496 494796 308508
rect 452068 308468 494796 308496
rect 452068 308456 452074 308468
rect 494790 308456 494796 308468
rect 494848 308456 494854 308508
rect 498838 308456 498844 308508
rect 498896 308496 498902 308508
rect 542630 308496 542636 308508
rect 498896 308468 542636 308496
rect 498896 308456 498902 308468
rect 542630 308456 542636 308468
rect 542688 308456 542694 308508
rect 457162 308388 457168 308440
rect 457220 308428 457226 308440
rect 536098 308428 536104 308440
rect 457220 308400 536104 308428
rect 457220 308388 457226 308400
rect 536098 308388 536104 308400
rect 536156 308388 536162 308440
rect 473998 307776 474004 307828
rect 474056 307816 474062 307828
rect 482646 307816 482652 307828
rect 474056 307788 482652 307816
rect 474056 307776 474062 307788
rect 482646 307776 482652 307788
rect 482704 307776 482710 307828
rect 3418 307708 3424 307760
rect 3476 307748 3482 307760
rect 4798 307748 4804 307760
rect 3476 307720 4804 307748
rect 3476 307708 3482 307720
rect 4798 307708 4804 307720
rect 4856 307708 4862 307760
rect 481082 307300 481088 307352
rect 481140 307340 481146 307352
rect 482462 307340 482468 307352
rect 481140 307312 482468 307340
rect 481140 307300 481146 307312
rect 482462 307300 482468 307312
rect 482520 307300 482526 307352
rect 454862 307164 454868 307216
rect 454920 307204 454926 307216
rect 490282 307204 490288 307216
rect 454920 307176 490288 307204
rect 454920 307164 454926 307176
rect 490282 307164 490288 307176
rect 490340 307164 490346 307216
rect 477310 307096 477316 307148
rect 477368 307136 477374 307148
rect 544378 307136 544384 307148
rect 477368 307108 544384 307136
rect 477368 307096 477374 307108
rect 544378 307096 544384 307108
rect 544436 307096 544442 307148
rect 380158 307028 380164 307080
rect 380216 307068 380222 307080
rect 506934 307068 506940 307080
rect 380216 307040 506940 307068
rect 380216 307028 380222 307040
rect 506934 307028 506940 307040
rect 506992 307028 506998 307080
rect 383194 306280 383200 306332
rect 383252 306320 383258 306332
rect 465442 306320 465448 306332
rect 383252 306292 465448 306320
rect 383252 306280 383258 306292
rect 465442 306280 465448 306292
rect 465500 306280 465506 306332
rect 381998 306212 382004 306264
rect 382056 306252 382062 306264
rect 465350 306252 465356 306264
rect 382056 306224 465356 306252
rect 382056 306212 382062 306224
rect 465350 306212 465356 306224
rect 465408 306212 465414 306264
rect 378870 306144 378876 306196
rect 378928 306184 378934 306196
rect 463786 306184 463792 306196
rect 378928 306156 463792 306184
rect 378928 306144 378934 306156
rect 463786 306144 463792 306156
rect 463844 306144 463850 306196
rect 384666 306076 384672 306128
rect 384724 306116 384730 306128
rect 475654 306116 475660 306128
rect 384724 306088 475660 306116
rect 384724 306076 384730 306088
rect 475654 306076 475660 306088
rect 475712 306076 475718 306128
rect 381814 306008 381820 306060
rect 381872 306048 381878 306060
rect 475102 306048 475108 306060
rect 381872 306020 475108 306048
rect 381872 306008 381878 306020
rect 475102 306008 475108 306020
rect 475160 306008 475166 306060
rect 378778 305940 378784 305992
rect 378836 305980 378842 305992
rect 475470 305980 475476 305992
rect 378836 305952 475476 305980
rect 378836 305940 378842 305952
rect 475470 305940 475476 305952
rect 475528 305940 475534 305992
rect 477402 305940 477408 305992
rect 477460 305980 477466 305992
rect 569218 305980 569224 305992
rect 477460 305952 569224 305980
rect 477460 305940 477466 305952
rect 569218 305940 569224 305952
rect 569276 305940 569282 305992
rect 384850 305872 384856 305924
rect 384908 305912 384914 305924
rect 486142 305912 486148 305924
rect 384908 305884 486148 305912
rect 384908 305872 384914 305884
rect 486142 305872 486148 305884
rect 486200 305872 486206 305924
rect 384482 305804 384488 305856
rect 384540 305844 384546 305856
rect 486510 305844 486516 305856
rect 384540 305816 486516 305844
rect 384540 305804 384546 305816
rect 486510 305804 486516 305816
rect 486568 305804 486574 305856
rect 381630 305736 381636 305788
rect 381688 305776 381694 305788
rect 486050 305776 486056 305788
rect 381688 305748 486056 305776
rect 381688 305736 381694 305748
rect 486050 305736 486056 305748
rect 486108 305736 486114 305788
rect 500126 305736 500132 305788
rect 500184 305776 500190 305788
rect 541066 305776 541072 305788
rect 500184 305748 541072 305776
rect 500184 305736 500190 305748
rect 541066 305736 541072 305748
rect 541124 305736 541130 305788
rect 365162 305668 365168 305720
rect 365220 305708 365226 305720
rect 516226 305708 516232 305720
rect 365220 305680 516232 305708
rect 365220 305668 365226 305680
rect 516226 305668 516232 305680
rect 516284 305668 516290 305720
rect 360838 305600 360844 305652
rect 360896 305640 360902 305652
rect 512086 305640 512092 305652
rect 360896 305612 512092 305640
rect 360896 305600 360902 305612
rect 512086 305600 512092 305612
rect 512144 305600 512150 305652
rect 384390 305532 384396 305584
rect 384448 305572 384454 305584
rect 465534 305572 465540 305584
rect 384448 305544 465540 305572
rect 384448 305532 384454 305544
rect 465534 305532 465540 305544
rect 465592 305532 465598 305584
rect 384574 305464 384580 305516
rect 384632 305504 384638 305516
rect 465166 305504 465172 305516
rect 384632 305476 465172 305504
rect 384632 305464 384638 305476
rect 465166 305464 465172 305476
rect 465224 305464 465230 305516
rect 458818 305396 458824 305448
rect 458876 305436 458882 305448
rect 488994 305436 489000 305448
rect 458876 305408 489000 305436
rect 458876 305396 458882 305408
rect 488994 305396 489000 305408
rect 489052 305396 489058 305448
rect 361758 304920 361764 304972
rect 361816 304960 361822 304972
rect 431218 304960 431224 304972
rect 361816 304932 431224 304960
rect 361816 304920 361822 304932
rect 431218 304920 431224 304932
rect 431276 304920 431282 304972
rect 488258 304512 488264 304564
rect 488316 304552 488322 304564
rect 531406 304552 531412 304564
rect 488316 304524 531412 304552
rect 488316 304512 488322 304524
rect 531406 304512 531412 304524
rect 531464 304512 531470 304564
rect 385770 304444 385776 304496
rect 385828 304484 385834 304496
rect 507026 304484 507032 304496
rect 385828 304456 507032 304484
rect 385828 304444 385834 304456
rect 507026 304444 507032 304456
rect 507084 304444 507090 304496
rect 383102 304376 383108 304428
rect 383160 304416 383166 304428
rect 520918 304416 520924 304428
rect 383160 304388 520924 304416
rect 383160 304376 383166 304388
rect 520918 304376 520924 304388
rect 520976 304376 520982 304428
rect 361022 304308 361028 304360
rect 361080 304348 361086 304360
rect 512178 304348 512184 304360
rect 361080 304320 512184 304348
rect 361080 304308 361086 304320
rect 512178 304308 512184 304320
rect 512236 304308 512242 304360
rect 360930 304240 360936 304292
rect 360988 304280 360994 304292
rect 512730 304280 512736 304292
rect 360988 304252 512736 304280
rect 360988 304240 360994 304252
rect 512730 304240 512736 304252
rect 512788 304240 512794 304292
rect 459370 304104 459376 304156
rect 459428 304144 459434 304156
rect 461670 304144 461676 304156
rect 459428 304116 461676 304144
rect 459428 304104 459434 304116
rect 461670 304104 461676 304116
rect 461728 304104 461734 304156
rect 378594 303560 378600 303612
rect 378652 303600 378658 303612
rect 484762 303600 484768 303612
rect 378652 303572 484768 303600
rect 378652 303560 378658 303572
rect 484762 303560 484768 303572
rect 484820 303560 484826 303612
rect 375834 303492 375840 303544
rect 375892 303532 375898 303544
rect 484486 303532 484492 303544
rect 375892 303504 484492 303532
rect 375892 303492 375898 303504
rect 484486 303492 484492 303504
rect 484544 303492 484550 303544
rect 371878 303424 371884 303476
rect 371936 303464 371942 303476
rect 485866 303464 485872 303476
rect 371936 303436 485872 303464
rect 371936 303424 371942 303436
rect 485866 303424 485872 303436
rect 485924 303424 485930 303476
rect 456334 303356 456340 303408
rect 456392 303396 456398 303408
rect 574738 303396 574744 303408
rect 456392 303368 574744 303396
rect 456392 303356 456398 303368
rect 574738 303356 574744 303368
rect 574796 303356 574802 303408
rect 376018 303288 376024 303340
rect 376076 303328 376082 303340
rect 509510 303328 509516 303340
rect 376076 303300 509516 303328
rect 376076 303288 376082 303300
rect 509510 303288 509516 303300
rect 509568 303288 509574 303340
rect 376478 303220 376484 303272
rect 376536 303260 376542 303272
rect 510798 303260 510804 303272
rect 376536 303232 510804 303260
rect 376536 303220 376542 303232
rect 510798 303220 510804 303232
rect 510856 303220 510862 303272
rect 379422 303152 379428 303204
rect 379480 303192 379486 303204
rect 515214 303192 515220 303204
rect 379480 303164 515220 303192
rect 379480 303152 379486 303164
rect 515214 303152 515220 303164
rect 515272 303152 515278 303204
rect 379238 303084 379244 303136
rect 379296 303124 379302 303136
rect 515306 303124 515312 303136
rect 379296 303096 515312 303124
rect 379296 303084 379302 303096
rect 515306 303084 515312 303096
rect 515364 303084 515370 303136
rect 376386 303016 376392 303068
rect 376444 303056 376450 303068
rect 513742 303056 513748 303068
rect 376444 303028 513748 303056
rect 376444 303016 376450 303028
rect 513742 303016 513748 303028
rect 513800 303016 513806 303068
rect 376570 302948 376576 303000
rect 376628 302988 376634 303000
rect 515122 302988 515128 303000
rect 376628 302960 515128 302988
rect 376628 302948 376634 302960
rect 515122 302948 515128 302960
rect 515180 302948 515186 303000
rect 367738 302880 367744 302932
rect 367796 302920 367802 302932
rect 512362 302920 512368 302932
rect 367796 302892 512368 302920
rect 367796 302880 367802 302892
rect 512362 302880 512368 302892
rect 512420 302880 512426 302932
rect 373718 302812 373724 302864
rect 373776 302852 373782 302864
rect 475378 302852 475384 302864
rect 373776 302824 475384 302852
rect 373776 302812 373782 302824
rect 475378 302812 475384 302824
rect 475436 302812 475442 302864
rect 376662 302744 376668 302796
rect 376720 302784 376726 302796
rect 474826 302784 474832 302796
rect 376720 302756 474832 302784
rect 376720 302744 376726 302756
rect 474826 302744 474832 302756
rect 474884 302744 474890 302796
rect 375926 302676 375932 302728
rect 375984 302716 375990 302728
rect 464062 302716 464068 302728
rect 375984 302688 464068 302716
rect 375984 302676 375990 302688
rect 464062 302676 464068 302688
rect 464120 302676 464126 302728
rect 478874 301656 478880 301708
rect 478932 301696 478938 301708
rect 481082 301696 481088 301708
rect 478932 301668 481088 301696
rect 478932 301656 478938 301668
rect 481082 301656 481088 301668
rect 481140 301656 481146 301708
rect 456610 301588 456616 301640
rect 456668 301628 456674 301640
rect 571978 301628 571984 301640
rect 456668 301600 571984 301628
rect 456668 301588 456674 301600
rect 571978 301588 571984 301600
rect 572036 301588 572042 301640
rect 367830 301520 367836 301572
rect 367888 301560 367894 301572
rect 512454 301560 512460 301572
rect 367888 301532 512460 301560
rect 367888 301520 367894 301532
rect 512454 301520 512460 301532
rect 512512 301520 512518 301572
rect 364978 301452 364984 301504
rect 365036 301492 365042 301504
rect 512546 301492 512552 301504
rect 365036 301464 512552 301492
rect 365036 301452 365042 301464
rect 512546 301452 512552 301464
rect 512604 301452 512610 301504
rect 373350 300772 373356 300824
rect 373408 300812 373414 300824
rect 510614 300812 510620 300824
rect 373408 300784 510620 300812
rect 373408 300772 373414 300784
rect 510614 300772 510620 300784
rect 510672 300772 510678 300824
rect 370866 300704 370872 300756
rect 370924 300744 370930 300756
rect 509326 300744 509332 300756
rect 370924 300716 509332 300744
rect 370924 300704 370930 300716
rect 509326 300704 509332 300716
rect 509384 300704 509390 300756
rect 373534 300636 373540 300688
rect 373592 300676 373598 300688
rect 513650 300676 513656 300688
rect 373592 300648 513656 300676
rect 373592 300636 373598 300648
rect 513650 300636 513656 300648
rect 513708 300636 513714 300688
rect 373442 300568 373448 300620
rect 373500 300608 373506 300620
rect 515030 300608 515036 300620
rect 373500 300580 515036 300608
rect 373500 300568 373506 300580
rect 515030 300568 515036 300580
rect 515088 300568 515094 300620
rect 370958 300500 370964 300552
rect 371016 300540 371022 300552
rect 513558 300540 513564 300552
rect 371016 300512 513564 300540
rect 371016 300500 371022 300512
rect 513558 300500 513564 300512
rect 513616 300500 513622 300552
rect 370774 300432 370780 300484
rect 370832 300472 370838 300484
rect 516410 300472 516416 300484
rect 370832 300444 516416 300472
rect 370832 300432 370838 300444
rect 516410 300432 516416 300444
rect 516468 300432 516474 300484
rect 367922 300364 367928 300416
rect 367980 300404 367986 300416
rect 514846 300404 514852 300416
rect 367980 300376 514852 300404
rect 367980 300364 367986 300376
rect 514846 300364 514852 300376
rect 514904 300364 514910 300416
rect 368198 300296 368204 300348
rect 368256 300336 368262 300348
rect 516318 300336 516324 300348
rect 368256 300308 516324 300336
rect 368256 300296 368262 300308
rect 516318 300296 516324 300308
rect 516376 300296 516382 300348
rect 363598 300228 363604 300280
rect 363656 300268 363662 300280
rect 512638 300268 512644 300280
rect 363656 300240 512644 300268
rect 363656 300228 363662 300240
rect 512638 300228 512644 300240
rect 512696 300228 512702 300280
rect 368014 300160 368020 300212
rect 368072 300200 368078 300212
rect 517606 300200 517612 300212
rect 368072 300172 517612 300200
rect 368072 300160 368078 300172
rect 517606 300160 517612 300172
rect 517664 300160 517670 300212
rect 361114 300092 361120 300144
rect 361172 300132 361178 300144
rect 512270 300132 512276 300144
rect 361172 300104 512276 300132
rect 361172 300092 361178 300104
rect 512270 300092 512276 300104
rect 512328 300092 512334 300144
rect 376202 300024 376208 300076
rect 376260 300064 376266 300076
rect 510154 300064 510160 300076
rect 376260 300036 510160 300064
rect 376260 300024 376266 300036
rect 510154 300024 510160 300036
rect 510212 300024 510218 300076
rect 467742 299956 467748 300008
rect 467800 299996 467806 300008
rect 580258 299996 580264 300008
rect 467800 299968 580264 299996
rect 467800 299956 467806 299968
rect 580258 299956 580264 299968
rect 580316 299956 580322 300008
rect 457530 299888 457536 299940
rect 457588 299928 457594 299940
rect 495802 299928 495808 299940
rect 457588 299900 495808 299928
rect 457588 299888 457594 299900
rect 495802 299888 495808 299900
rect 495860 299888 495866 299940
rect 461578 299412 461584 299464
rect 461636 299452 461642 299464
rect 580166 299452 580172 299464
rect 461636 299424 580172 299452
rect 461636 299412 461642 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 478138 298936 478144 298988
rect 478196 298976 478202 298988
rect 478874 298976 478880 298988
rect 478196 298948 478880 298976
rect 478196 298936 478202 298948
rect 478874 298936 478880 298948
rect 478932 298936 478938 298988
rect 456702 297984 456708 298036
rect 456760 298024 456766 298036
rect 573358 298024 573364 298036
rect 456760 297996 573364 298024
rect 456760 297984 456766 297996
rect 573358 297984 573364 297996
rect 573416 297984 573422 298036
rect 383010 297916 383016 297968
rect 383068 297956 383074 297968
rect 518250 297956 518256 297968
rect 383068 297928 518256 297956
rect 383068 297916 383074 297928
rect 518250 297916 518256 297928
rect 518308 297916 518314 297968
rect 363966 297848 363972 297900
rect 364024 297888 364030 297900
rect 507670 297888 507676 297900
rect 364024 297860 507676 297888
rect 364024 297848 364030 297860
rect 507670 297848 507676 297860
rect 507728 297848 507734 297900
rect 362494 297780 362500 297832
rect 362552 297820 362558 297832
rect 507762 297820 507768 297832
rect 362552 297792 507768 297820
rect 362552 297780 362558 297792
rect 507762 297780 507768 297792
rect 507820 297780 507826 297832
rect 368106 297712 368112 297764
rect 368164 297752 368170 297764
rect 518066 297752 518072 297764
rect 368164 297724 518072 297752
rect 368164 297712 368170 297724
rect 518066 297712 518072 297724
rect 518124 297712 518130 297764
rect 366542 297644 366548 297696
rect 366600 297684 366606 297696
rect 516686 297684 516692 297696
rect 366600 297656 516692 297684
rect 366600 297644 366606 297656
rect 516686 297644 516692 297656
rect 516744 297644 516750 297696
rect 362310 297576 362316 297628
rect 362368 297616 362374 297628
rect 513926 297616 513932 297628
rect 362368 297588 513932 297616
rect 362368 297576 362374 297588
rect 513926 297576 513932 297588
rect 513984 297576 513990 297628
rect 363782 297508 363788 297560
rect 363840 297548 363846 297560
rect 515582 297548 515588 297560
rect 363840 297520 515588 297548
rect 363840 297508 363846 297520
rect 515582 297508 515588 297520
rect 515640 297508 515646 297560
rect 365438 297440 365444 297492
rect 365496 297480 365502 297492
rect 518342 297480 518348 297492
rect 365496 297452 518348 297480
rect 365496 297440 365502 297452
rect 518342 297440 518348 297452
rect 518400 297440 518406 297492
rect 363874 297372 363880 297424
rect 363932 297412 363938 297424
rect 516778 297412 516784 297424
rect 363932 297384 516784 297412
rect 363932 297372 363938 297384
rect 516778 297372 516784 297384
rect 516836 297372 516842 297424
rect 460382 296692 460388 296744
rect 460440 296732 460446 296744
rect 462958 296732 462964 296744
rect 460440 296704 462964 296732
rect 460440 296692 460446 296704
rect 462958 296692 462964 296704
rect 463016 296692 463022 296744
rect 457990 295944 457996 295996
rect 458048 295984 458054 295996
rect 576118 295984 576124 295996
rect 458048 295956 576124 295984
rect 458048 295944 458054 295956
rect 576118 295944 576124 295956
rect 576176 295944 576182 295996
rect 476850 295332 476856 295384
rect 476908 295372 476914 295384
rect 478138 295372 478144 295384
rect 476908 295344 478144 295372
rect 476908 295332 476914 295344
rect 478138 295332 478144 295344
rect 478196 295332 478202 295384
rect 374914 295264 374920 295316
rect 374972 295304 374978 295316
rect 514202 295304 514208 295316
rect 374972 295276 514208 295304
rect 374972 295264 374978 295276
rect 514202 295264 514208 295276
rect 514260 295264 514266 295316
rect 381446 295196 381452 295248
rect 381504 295236 381510 295248
rect 520550 295236 520556 295248
rect 381504 295208 520556 295236
rect 381504 295196 381510 295208
rect 520550 295196 520556 295208
rect 520608 295196 520614 295248
rect 369302 295128 369308 295180
rect 369360 295168 369366 295180
rect 510706 295168 510712 295180
rect 369360 295140 510712 295168
rect 369360 295128 369366 295140
rect 510706 295128 510712 295140
rect 510764 295128 510770 295180
rect 374822 295060 374828 295112
rect 374880 295100 374886 295112
rect 517698 295100 517704 295112
rect 374880 295072 517704 295100
rect 374880 295060 374886 295072
rect 517698 295060 517704 295072
rect 517756 295060 517762 295112
rect 374730 294992 374736 295044
rect 374788 295032 374794 295044
rect 517882 295032 517888 295044
rect 374788 295004 517888 295032
rect 374788 294992 374794 295004
rect 517882 294992 517888 295004
rect 517940 294992 517946 295044
rect 376294 294924 376300 294976
rect 376352 294964 376358 294976
rect 520458 294964 520464 294976
rect 376352 294936 520464 294964
rect 376352 294924 376358 294936
rect 520458 294924 520464 294936
rect 520516 294924 520522 294976
rect 373626 294856 373632 294908
rect 373684 294896 373690 294908
rect 519078 294896 519084 294908
rect 373684 294868 519084 294896
rect 373684 294856 373690 294868
rect 519078 294856 519084 294868
rect 519136 294856 519142 294908
rect 372246 294788 372252 294840
rect 372304 294828 372310 294840
rect 519170 294828 519176 294840
rect 372304 294800 519176 294828
rect 372304 294788 372310 294800
rect 519170 294788 519176 294800
rect 519228 294788 519234 294840
rect 370682 294720 370688 294772
rect 370740 294760 370746 294772
rect 519354 294760 519360 294772
rect 370740 294732 519360 294760
rect 370740 294720 370746 294732
rect 519354 294720 519360 294732
rect 519412 294720 519418 294772
rect 366634 294652 366640 294704
rect 366692 294692 366698 294704
rect 516502 294692 516508 294704
rect 366692 294664 516508 294692
rect 366692 294652 366698 294664
rect 516502 294652 516508 294664
rect 516560 294652 516566 294704
rect 369394 294584 369400 294636
rect 369452 294624 369458 294636
rect 519446 294624 519452 294636
rect 369452 294596 519452 294624
rect 369452 294584 369458 294596
rect 519446 294584 519452 294596
rect 519504 294584 519510 294636
rect 372154 294516 372160 294568
rect 372212 294556 372218 294568
rect 509418 294556 509424 294568
rect 372212 294528 509424 294556
rect 372212 294516 372218 294528
rect 509418 294516 509424 294528
rect 509476 294516 509482 294568
rect 457714 294448 457720 294500
rect 457772 294488 457778 294500
rect 570690 294488 570696 294500
rect 457772 294460 570696 294488
rect 457772 294448 457778 294460
rect 570690 294448 570696 294460
rect 570748 294448 570754 294500
rect 361758 293904 361764 293956
rect 361816 293944 361822 293956
rect 435358 293944 435364 293956
rect 361816 293916 435364 293944
rect 361816 293904 361822 293916
rect 435358 293904 435364 293916
rect 435416 293904 435422 293956
rect 488350 293292 488356 293344
rect 488408 293332 488414 293344
rect 530026 293332 530032 293344
rect 488408 293304 530032 293332
rect 488408 293292 488414 293304
rect 530026 293292 530032 293304
rect 530084 293292 530090 293344
rect 467558 293224 467564 293276
rect 467616 293264 467622 293276
rect 559558 293264 559564 293276
rect 467616 293236 559564 293264
rect 467616 293224 467622 293236
rect 559558 293224 559564 293236
rect 559616 293224 559622 293276
rect 3326 292544 3332 292596
rect 3384 292584 3390 292596
rect 19978 292584 19984 292596
rect 3384 292556 19984 292584
rect 3384 292544 3390 292556
rect 19978 292544 19984 292556
rect 20036 292544 20042 292596
rect 384298 292476 384304 292528
rect 384356 292516 384362 292528
rect 507394 292516 507400 292528
rect 384356 292488 507400 292516
rect 384356 292476 384362 292488
rect 507394 292476 507400 292488
rect 507452 292476 507458 292528
rect 386046 292408 386052 292460
rect 386104 292448 386110 292460
rect 520826 292448 520832 292460
rect 386104 292420 520832 292448
rect 386104 292408 386110 292420
rect 520826 292408 520832 292420
rect 520884 292408 520890 292460
rect 383470 292340 383476 292392
rect 383528 292380 383534 292392
rect 518894 292380 518900 292392
rect 383528 292352 518900 292380
rect 383528 292340 383534 292352
rect 518894 292340 518900 292352
rect 518952 292340 518958 292392
rect 377674 292272 377680 292324
rect 377732 292312 377738 292324
rect 514754 292312 514760 292324
rect 377732 292284 514760 292312
rect 377732 292272 377738 292284
rect 514754 292272 514760 292284
rect 514812 292272 514818 292324
rect 379054 292204 379060 292256
rect 379112 292244 379118 292256
rect 516870 292244 516876 292256
rect 379112 292216 516876 292244
rect 379112 292204 379118 292216
rect 516870 292204 516876 292216
rect 516928 292204 516934 292256
rect 375098 292136 375104 292188
rect 375156 292176 375162 292188
rect 514110 292176 514116 292188
rect 375156 292148 514116 292176
rect 375156 292136 375162 292148
rect 514110 292136 514116 292148
rect 514168 292136 514174 292188
rect 369210 292068 369216 292120
rect 369268 292108 369274 292120
rect 507486 292108 507492 292120
rect 369268 292080 507492 292108
rect 369268 292068 369274 292080
rect 507486 292068 507492 292080
rect 507544 292068 507550 292120
rect 380526 292000 380532 292052
rect 380584 292040 380590 292052
rect 520274 292040 520280 292052
rect 380584 292012 520280 292040
rect 380584 292000 380590 292012
rect 520274 292000 520280 292012
rect 520332 292000 520338 292052
rect 377766 291932 377772 291984
rect 377824 291972 377830 291984
rect 520366 291972 520372 291984
rect 377824 291944 520372 291972
rect 377824 291932 377830 291944
rect 520366 291932 520372 291944
rect 520424 291932 520430 291984
rect 366358 291864 366364 291916
rect 366416 291904 366422 291916
rect 516594 291904 516600 291916
rect 366416 291876 516600 291904
rect 366416 291864 366422 291876
rect 516594 291864 516600 291876
rect 516652 291864 516658 291916
rect 363690 291796 363696 291848
rect 363748 291836 363754 291848
rect 519722 291836 519728 291848
rect 363748 291808 519728 291836
rect 363748 291796 363754 291808
rect 519722 291796 519728 291808
rect 519780 291796 519786 291848
rect 385954 291728 385960 291780
rect 386012 291768 386018 291780
rect 507578 291768 507584 291780
rect 386012 291740 507584 291768
rect 386012 291728 386018 291740
rect 507578 291728 507584 291740
rect 507636 291728 507642 291780
rect 471238 291660 471244 291712
rect 471296 291700 471302 291712
rect 473998 291700 474004 291712
rect 471296 291672 474004 291700
rect 471296 291660 471302 291672
rect 473998 291660 474004 291672
rect 474056 291660 474062 291712
rect 478414 291660 478420 291712
rect 478472 291700 478478 291712
rect 559650 291700 559656 291712
rect 478472 291672 559656 291700
rect 478472 291660 478478 291672
rect 559650 291660 559656 291672
rect 559708 291660 559714 291712
rect 467650 290436 467656 290488
rect 467708 290476 467714 290488
rect 558178 290476 558184 290488
rect 467708 290448 558184 290476
rect 467708 290436 467714 290448
rect 558178 290436 558184 290448
rect 558236 290436 558242 290488
rect 375006 289756 375012 289808
rect 375064 289796 375070 289808
rect 507302 289796 507308 289808
rect 375064 289768 507308 289796
rect 375064 289756 375070 289768
rect 507302 289756 507308 289768
rect 507360 289756 507366 289808
rect 384758 289688 384764 289740
rect 384816 289728 384822 289740
rect 518986 289728 518992 289740
rect 384816 289700 518992 289728
rect 384816 289688 384822 289700
rect 518986 289688 518992 289700
rect 519044 289688 519050 289740
rect 380250 289620 380256 289672
rect 380308 289660 380314 289672
rect 517790 289660 517796 289672
rect 380308 289632 517796 289660
rect 380308 289620 380314 289632
rect 517790 289620 517796 289632
rect 517848 289620 517854 289672
rect 382182 289552 382188 289604
rect 382240 289592 382246 289604
rect 521838 289592 521844 289604
rect 382240 289564 521844 289592
rect 382240 289552 382246 289564
rect 521838 289552 521844 289564
rect 521896 289552 521902 289604
rect 383286 289484 383292 289536
rect 383344 289524 383350 289536
rect 523218 289524 523224 289536
rect 383344 289496 523224 289524
rect 383344 289484 383350 289496
rect 523218 289484 523224 289496
rect 523276 289484 523282 289536
rect 377582 289416 377588 289468
rect 377640 289456 377646 289468
rect 519262 289456 519268 289468
rect 377640 289428 519268 289456
rect 377640 289416 377646 289428
rect 519262 289416 519268 289428
rect 519320 289416 519326 289468
rect 380342 289348 380348 289400
rect 380400 289388 380406 289400
rect 523310 289388 523316 289400
rect 380400 289360 523316 289388
rect 380400 289348 380406 289360
rect 523310 289348 523316 289360
rect 523368 289348 523374 289400
rect 378962 289280 378968 289332
rect 379020 289320 379026 289332
rect 523126 289320 523132 289332
rect 379020 289292 523132 289320
rect 379020 289280 379026 289292
rect 523126 289280 523132 289292
rect 523184 289280 523190 289332
rect 377490 289212 377496 289264
rect 377548 289252 377554 289264
rect 521930 289252 521936 289264
rect 377548 289224 521936 289252
rect 377548 289212 377554 289224
rect 521930 289212 521936 289224
rect 521988 289212 521994 289264
rect 376110 289144 376116 289196
rect 376168 289184 376174 289196
rect 521746 289184 521752 289196
rect 376168 289156 521752 289184
rect 376168 289144 376174 289156
rect 521746 289144 521752 289156
rect 521804 289144 521810 289196
rect 372338 289076 372344 289128
rect 372396 289116 372402 289128
rect 520642 289116 520648 289128
rect 372396 289088 520648 289116
rect 372396 289076 372402 289088
rect 520642 289076 520648 289088
rect 520700 289076 520706 289128
rect 383378 289008 383384 289060
rect 383436 289048 383442 289060
rect 514938 289048 514944 289060
rect 383436 289020 514944 289048
rect 383436 289008 383442 289020
rect 514938 289008 514944 289020
rect 514996 289008 515002 289060
rect 385862 288940 385868 288992
rect 385920 288980 385926 288992
rect 507210 288980 507216 288992
rect 385920 288952 507216 288980
rect 385920 288940 385926 288952
rect 507210 288940 507216 288952
rect 507268 288940 507274 288992
rect 467282 288872 467288 288924
rect 467340 288912 467346 288924
rect 555418 288912 555424 288924
rect 467340 288884 555424 288912
rect 467340 288872 467346 288884
rect 555418 288872 555424 288884
rect 555476 288872 555482 288924
rect 475378 287784 475384 287836
rect 475436 287824 475442 287836
rect 476850 287824 476856 287836
rect 475436 287796 476856 287824
rect 475436 287784 475442 287796
rect 476850 287784 476856 287796
rect 476908 287784 476914 287836
rect 461394 286696 461400 286748
rect 461452 286736 461458 286748
rect 471238 286736 471244 286748
rect 461452 286708 471244 286736
rect 461452 286696 461458 286708
rect 471238 286696 471244 286708
rect 471296 286696 471302 286748
rect 452102 286628 452108 286680
rect 452160 286668 452166 286680
rect 490834 286668 490840 286680
rect 452160 286640 490840 286668
rect 452160 286628 452166 286640
rect 490834 286628 490840 286640
rect 490892 286628 490898 286680
rect 370498 286560 370504 286612
rect 370556 286600 370562 286612
rect 476482 286600 476488 286612
rect 370556 286572 476488 286600
rect 370556 286560 370562 286572
rect 476482 286560 476488 286572
rect 476540 286560 476546 286612
rect 488074 286560 488080 286612
rect 488132 286600 488138 286612
rect 531314 286600 531320 286612
rect 488132 286572 531320 286600
rect 488132 286560 488138 286572
rect 531314 286560 531320 286572
rect 531372 286560 531378 286612
rect 372062 286492 372068 286544
rect 372120 286532 372126 286544
rect 507118 286532 507124 286544
rect 372120 286504 507124 286532
rect 372120 286492 372126 286504
rect 507118 286492 507124 286504
rect 507176 286492 507182 286544
rect 377398 286424 377404 286476
rect 377456 286464 377462 286476
rect 520734 286464 520740 286476
rect 377456 286436 520740 286464
rect 377456 286424 377462 286436
rect 520734 286424 520740 286436
rect 520792 286424 520798 286476
rect 366450 286356 366456 286408
rect 366508 286396 366514 286408
rect 521654 286396 521660 286408
rect 366508 286368 521660 286396
rect 366508 286356 366514 286368
rect 521654 286356 521660 286368
rect 521712 286356 521718 286408
rect 365254 286288 365260 286340
rect 365312 286328 365318 286340
rect 523034 286328 523040 286340
rect 365312 286300 523040 286328
rect 365312 286288 365318 286300
rect 523034 286288 523040 286300
rect 523092 286288 523098 286340
rect 453298 284928 453304 284980
rect 453356 284968 453362 284980
rect 489178 284968 489184 284980
rect 453356 284940 489184 284968
rect 453356 284928 453362 284940
rect 489178 284928 489184 284940
rect 489236 284928 489242 284980
rect 498010 284928 498016 284980
rect 498068 284968 498074 284980
rect 539870 284968 539876 284980
rect 498068 284940 539876 284968
rect 498068 284928 498074 284940
rect 539870 284928 539876 284940
rect 539928 284928 539934 284980
rect 452378 283568 452384 283620
rect 452436 283608 452442 283620
rect 494974 283608 494980 283620
rect 452436 283580 494980 283608
rect 452436 283568 452442 283580
rect 494974 283568 494980 283580
rect 495032 283568 495038 283620
rect 459462 282888 459468 282940
rect 459520 282928 459526 282940
rect 460382 282928 460388 282940
rect 459520 282900 460388 282928
rect 459520 282888 459526 282900
rect 460382 282888 460388 282900
rect 460440 282888 460446 282940
rect 361758 282820 361764 282872
rect 361816 282860 361822 282872
rect 436830 282860 436836 282872
rect 361816 282832 436836 282860
rect 361816 282820 361822 282832
rect 436830 282820 436836 282832
rect 436888 282820 436894 282872
rect 459278 282140 459284 282192
rect 459336 282180 459342 282192
rect 494146 282180 494152 282192
rect 459336 282152 494152 282180
rect 459336 282140 459342 282152
rect 494146 282140 494152 282152
rect 494204 282140 494210 282192
rect 455046 280780 455052 280832
rect 455104 280820 455110 280832
rect 493410 280820 493416 280832
rect 455104 280792 493416 280820
rect 455104 280780 455110 280792
rect 493410 280780 493416 280792
rect 493468 280780 493474 280832
rect 453666 279488 453672 279540
rect 453724 279528 453730 279540
rect 461394 279528 461400 279540
rect 453724 279500 461400 279528
rect 453724 279488 453730 279500
rect 461394 279488 461400 279500
rect 461452 279488 461458 279540
rect 453390 279420 453396 279472
rect 453448 279460 453454 279472
rect 490650 279460 490656 279472
rect 453448 279432 490656 279460
rect 453448 279420 453454 279432
rect 490650 279420 490656 279432
rect 490708 279420 490714 279472
rect 503622 279420 503628 279472
rect 503680 279460 503686 279472
rect 539042 279460 539048 279472
rect 503680 279432 539048 279460
rect 503680 279420 503686 279432
rect 539042 279420 539048 279432
rect 539100 279420 539106 279472
rect 453482 278060 453488 278112
rect 453540 278100 453546 278112
rect 490006 278100 490012 278112
rect 453540 278072 490012 278100
rect 453540 278060 453546 278072
rect 490006 278060 490012 278072
rect 490064 278060 490070 278112
rect 381354 277992 381360 278044
rect 381412 278032 381418 278044
rect 486418 278032 486424 278044
rect 381412 278004 486424 278032
rect 381412 277992 381418 278004
rect 486418 277992 486424 278004
rect 486476 277992 486482 278044
rect 501782 277992 501788 278044
rect 501840 278032 501846 278044
rect 540238 278032 540244 278044
rect 501840 278004 540244 278032
rect 501840 277992 501846 278004
rect 540238 277992 540244 278004
rect 540296 277992 540302 278044
rect 455230 276632 455236 276684
rect 455288 276672 455294 276684
rect 494698 276672 494704 276684
rect 455288 276644 494704 276672
rect 455288 276632 455294 276644
rect 494698 276632 494704 276644
rect 494756 276632 494762 276684
rect 500218 276632 500224 276684
rect 500276 276672 500282 276684
rect 539962 276672 539968 276684
rect 500276 276644 539968 276672
rect 500276 276632 500282 276644
rect 539962 276632 539968 276644
rect 540020 276632 540026 276684
rect 459186 275272 459192 275324
rect 459244 275312 459250 275324
rect 493134 275312 493140 275324
rect 459244 275284 493140 275312
rect 459244 275272 459250 275284
rect 493134 275272 493140 275284
rect 493192 275272 493198 275324
rect 499022 275272 499028 275324
rect 499080 275312 499086 275324
rect 541250 275312 541256 275324
rect 499080 275284 541256 275312
rect 499080 275272 499086 275284
rect 541250 275272 541256 275284
rect 541308 275272 541314 275324
rect 473354 274660 473360 274712
rect 473412 274700 473418 274712
rect 475378 274700 475384 274712
rect 473412 274672 475384 274700
rect 473412 274660 473418 274672
rect 475378 274660 475384 274672
rect 475436 274660 475442 274712
rect 457622 273980 457628 274032
rect 457680 274020 457686 274032
rect 491386 274020 491392 274032
rect 457680 273992 491392 274020
rect 457680 273980 457686 273992
rect 491386 273980 491392 273992
rect 491444 273980 491450 274032
rect 499390 273980 499396 274032
rect 499448 274020 499454 274032
rect 541342 274020 541348 274032
rect 499448 273992 541348 274020
rect 499448 273980 499454 273992
rect 541342 273980 541348 273992
rect 541400 273980 541406 274032
rect 452194 273912 452200 273964
rect 452252 273952 452258 273964
rect 488626 273952 488632 273964
rect 452252 273924 488632 273952
rect 452252 273912 452258 273924
rect 488626 273912 488632 273924
rect 488684 273912 488690 273964
rect 497734 273912 497740 273964
rect 497792 273952 497798 273964
rect 542814 273952 542820 273964
rect 497792 273924 542820 273952
rect 497792 273912 497798 273924
rect 542814 273912 542820 273924
rect 542872 273912 542878 273964
rect 479518 273164 479524 273216
rect 479576 273204 479582 273216
rect 579890 273204 579896 273216
rect 479576 273176 579896 273204
rect 479576 273164 479582 273176
rect 579890 273164 579896 273176
rect 579948 273164 579954 273216
rect 453574 272552 453580 272604
rect 453632 272592 453638 272604
rect 488902 272592 488908 272604
rect 453632 272564 488908 272592
rect 453632 272552 453638 272564
rect 488902 272552 488908 272564
rect 488960 272552 488966 272604
rect 455138 272484 455144 272536
rect 455196 272524 455202 272536
rect 492766 272524 492772 272536
rect 455196 272496 492772 272524
rect 455196 272484 455202 272496
rect 492766 272484 492772 272496
rect 492824 272484 492830 272536
rect 500770 272484 500776 272536
rect 500828 272524 500834 272536
rect 541434 272524 541440 272536
rect 500828 272496 541440 272524
rect 500828 272484 500834 272496
rect 541434 272484 541440 272496
rect 541492 272484 541498 272536
rect 361758 271804 361764 271856
rect 361816 271844 361822 271856
rect 439682 271844 439688 271856
rect 361816 271816 439688 271844
rect 361816 271804 361822 271816
rect 439682 271804 439688 271816
rect 439740 271804 439746 271856
rect 459094 271192 459100 271244
rect 459152 271232 459158 271244
rect 491662 271232 491668 271244
rect 459152 271204 491668 271232
rect 459152 271192 459158 271204
rect 491662 271192 491668 271204
rect 491720 271192 491726 271244
rect 500494 271192 500500 271244
rect 500552 271232 500558 271244
rect 540146 271232 540152 271244
rect 500552 271204 540152 271232
rect 500552 271192 500558 271204
rect 540146 271192 540152 271204
rect 540204 271192 540210 271244
rect 457714 271124 457720 271176
rect 457772 271164 457778 271176
rect 493318 271164 493324 271176
rect 457772 271136 493324 271164
rect 457772 271124 457778 271136
rect 493318 271124 493324 271136
rect 493376 271124 493382 271176
rect 499114 271124 499120 271176
rect 499172 271164 499178 271176
rect 540054 271164 540060 271176
rect 499172 271136 540060 271164
rect 499172 271124 499178 271136
rect 540054 271124 540060 271136
rect 540112 271124 540118 271176
rect 456242 271056 456248 271108
rect 456300 271096 456306 271108
rect 459462 271096 459468 271108
rect 456300 271068 459468 271096
rect 456300 271056 456306 271068
rect 459462 271056 459468 271068
rect 459520 271056 459526 271108
rect 456702 269900 456708 269952
rect 456760 269940 456766 269952
rect 473722 269940 473728 269952
rect 456760 269912 473728 269940
rect 456760 269900 456766 269912
rect 473722 269900 473728 269912
rect 473780 269900 473786 269952
rect 505002 269900 505008 269952
rect 505060 269940 505066 269952
rect 543734 269940 543740 269952
rect 505060 269912 543740 269940
rect 505060 269900 505066 269912
rect 543734 269900 543740 269912
rect 543792 269900 543798 269952
rect 456150 269832 456156 269884
rect 456208 269872 456214 269884
rect 487246 269872 487252 269884
rect 456208 269844 487252 269872
rect 456208 269832 456214 269844
rect 487246 269832 487252 269844
rect 487304 269832 487310 269884
rect 496722 269832 496728 269884
rect 496780 269872 496786 269884
rect 541158 269872 541164 269884
rect 496780 269844 541164 269872
rect 496780 269832 496786 269844
rect 541158 269832 541164 269844
rect 541216 269832 541222 269884
rect 468754 269764 468760 269816
rect 468812 269804 468818 269816
rect 580350 269804 580356 269816
rect 468812 269776 580356 269804
rect 468812 269764 468818 269776
rect 580350 269764 580356 269776
rect 580408 269764 580414 269816
rect 459554 268540 459560 268592
rect 459612 268580 459618 268592
rect 473354 268580 473360 268592
rect 459612 268552 473360 268580
rect 459612 268540 459618 268552
rect 473354 268540 473360 268552
rect 473412 268540 473418 268592
rect 452286 268472 452292 268524
rect 452344 268512 452350 268524
rect 490558 268512 490564 268524
rect 452344 268484 490564 268512
rect 452344 268472 452350 268484
rect 490558 268472 490564 268484
rect 490616 268472 490622 268524
rect 466362 268404 466368 268456
rect 466420 268444 466426 268456
rect 570598 268444 570604 268456
rect 466420 268416 570604 268444
rect 466420 268404 466426 268416
rect 570598 268404 570604 268416
rect 570656 268404 570662 268456
rect 361206 268336 361212 268388
rect 361264 268376 361270 268388
rect 511994 268376 512000 268388
rect 361264 268348 512000 268376
rect 361264 268336 361270 268348
rect 511994 268336 512000 268348
rect 512052 268336 512058 268388
rect 3602 266364 3608 266416
rect 3660 266404 3666 266416
rect 4890 266404 4896 266416
rect 3660 266376 4896 266404
rect 3660 266364 3666 266376
rect 4890 266364 4896 266376
rect 4948 266364 4954 266416
rect 456886 266364 456892 266416
rect 456944 266404 456950 266416
rect 459554 266404 459560 266416
rect 456944 266376 459560 266404
rect 456944 266364 456950 266376
rect 459554 266364 459560 266376
rect 459612 266364 459618 266416
rect 453942 263576 453948 263628
rect 454000 263616 454006 263628
rect 456886 263616 456892 263628
rect 454000 263588 456892 263616
rect 454000 263576 454006 263588
rect 456886 263576 456892 263588
rect 456944 263576 456950 263628
rect 449802 263508 449808 263560
rect 449860 263548 449866 263560
rect 456794 263548 456800 263560
rect 449860 263520 456800 263548
rect 449860 263508 449866 263520
rect 456794 263508 456800 263520
rect 456852 263508 456858 263560
rect 448514 262896 448520 262948
rect 448572 262936 448578 262948
rect 456702 262936 456708 262948
rect 448572 262908 456708 262936
rect 448572 262896 448578 262908
rect 456702 262896 456708 262908
rect 456760 262896 456766 262948
rect 420178 262828 420184 262880
rect 420236 262868 420242 262880
rect 453666 262868 453672 262880
rect 420236 262840 453672 262868
rect 420236 262828 420242 262840
rect 453666 262828 453672 262840
rect 453724 262828 453730 262880
rect 361758 260788 361764 260840
rect 361816 260828 361822 260840
rect 440878 260828 440884 260840
rect 361816 260800 440884 260828
rect 361816 260788 361822 260800
rect 440878 260788 440884 260800
rect 440936 260788 440942 260840
rect 437750 258680 437756 258732
rect 437808 258720 437814 258732
rect 448514 258720 448520 258732
rect 437808 258692 448520 258720
rect 437808 258680 437814 258692
rect 448514 258680 448520 258692
rect 448572 258680 448578 258732
rect 449158 258068 449164 258120
rect 449216 258108 449222 258120
rect 453942 258108 453948 258120
rect 449216 258080 453948 258108
rect 449216 258068 449222 258080
rect 453942 258068 453948 258080
rect 454000 258068 454006 258120
rect 414658 256708 414664 256760
rect 414716 256748 414722 256760
rect 420178 256748 420184 256760
rect 414716 256720 420184 256748
rect 414716 256708 414722 256720
rect 420178 256708 420184 256720
rect 420236 256708 420242 256760
rect 429838 253172 429844 253224
rect 429896 253212 429902 253224
rect 437750 253212 437756 253224
rect 429896 253184 437756 253212
rect 429896 253172 429902 253184
rect 437750 253172 437756 253184
rect 437808 253172 437814 253224
rect 456886 250928 456892 250980
rect 456944 250968 456950 250980
rect 459370 250968 459376 250980
rect 456944 250940 459376 250968
rect 456944 250928 456950 250940
rect 459370 250928 459376 250940
rect 459428 250928 459434 250980
rect 361758 249704 361764 249756
rect 361816 249744 361822 249756
rect 399478 249744 399484 249756
rect 361816 249716 399484 249744
rect 361816 249704 361822 249716
rect 399478 249704 399484 249716
rect 399536 249704 399542 249756
rect 447134 249704 447140 249756
rect 447192 249744 447198 249756
rect 456794 249744 456800 249756
rect 447192 249716 456800 249744
rect 447192 249704 447198 249716
rect 456794 249704 456800 249716
rect 456852 249704 456858 249756
rect 446398 248888 446404 248940
rect 446456 248928 446462 248940
rect 447134 248928 447140 248940
rect 446456 248900 447140 248928
rect 446456 248888 446462 248900
rect 447134 248888 447140 248900
rect 447192 248888 447198 248940
rect 447226 247664 447232 247716
rect 447284 247704 447290 247716
rect 456886 247704 456892 247716
rect 447284 247676 456892 247704
rect 447284 247664 447290 247676
rect 456886 247664 456892 247676
rect 456944 247664 456950 247716
rect 449158 247092 449164 247104
rect 447152 247064 449164 247092
rect 445754 246984 445760 247036
rect 445812 247024 445818 247036
rect 447152 247024 447180 247064
rect 449158 247052 449164 247064
rect 449216 247052 449222 247104
rect 445812 246996 447180 247024
rect 445812 246984 445818 246996
rect 447226 245664 447232 245676
rect 445772 245636 447232 245664
rect 445662 245556 445668 245608
rect 445720 245596 445726 245608
rect 445772 245596 445800 245636
rect 447226 245624 447232 245636
rect 447284 245624 447290 245676
rect 445720 245568 445800 245596
rect 445720 245556 445726 245568
rect 570690 245556 570696 245608
rect 570748 245596 570754 245608
rect 580166 245596 580172 245608
rect 570748 245568 580172 245596
rect 570748 245556 570754 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 449158 243516 449164 243568
rect 449216 243556 449222 243568
rect 456242 243556 456248 243568
rect 449216 243528 456248 243556
rect 449216 243516 449222 243528
rect 456242 243516 456248 243528
rect 456300 243516 456306 243568
rect 3970 241408 3976 241460
rect 4028 241448 4034 241460
rect 5074 241448 5080 241460
rect 4028 241420 5080 241448
rect 4028 241408 4034 241420
rect 5074 241408 5080 241420
rect 5132 241408 5138 241460
rect 427078 241408 427084 241460
rect 427136 241448 427142 241460
rect 429838 241448 429844 241460
rect 427136 241420 429844 241448
rect 427136 241408 427142 241420
rect 429838 241408 429844 241420
rect 429896 241408 429902 241460
rect 443178 241136 443184 241188
rect 443236 241176 443242 241188
rect 445662 241176 445668 241188
rect 443236 241148 445668 241176
rect 443236 241136 443242 241148
rect 445662 241136 445668 241148
rect 445720 241136 445726 241188
rect 445202 239776 445208 239828
rect 445260 239816 445266 239828
rect 445754 239816 445760 239828
rect 445260 239788 445760 239816
rect 445260 239776 445266 239788
rect 445754 239776 445760 239788
rect 445812 239776 445818 239828
rect 361758 238688 361764 238740
rect 361816 238728 361822 238740
rect 443730 238728 443736 238740
rect 361816 238700 443736 238728
rect 361816 238688 361822 238700
rect 443730 238688 443736 238700
rect 443788 238688 443794 238740
rect 442258 237396 442264 237448
rect 442316 237436 442322 237448
rect 443178 237436 443184 237448
rect 442316 237408 443184 237436
rect 442316 237396 442322 237408
rect 443178 237396 443184 237408
rect 443236 237396 443242 237448
rect 443914 237396 443920 237448
rect 443972 237436 443978 237448
rect 445202 237436 445208 237448
rect 443972 237408 445208 237436
rect 443972 237396 443978 237408
rect 445202 237396 445208 237408
rect 445260 237396 445266 237448
rect 450722 235220 450728 235272
rect 450780 235260 450786 235272
rect 456794 235260 456800 235272
rect 450780 235232 456800 235260
rect 450780 235220 450786 235232
rect 456794 235220 456800 235232
rect 456852 235220 456858 235272
rect 3786 233180 3792 233232
rect 3844 233220 3850 233232
rect 4982 233220 4988 233232
rect 3844 233192 4988 233220
rect 3844 233180 3850 233192
rect 4982 233180 4988 233192
rect 5040 233180 5046 233232
rect 559650 233180 559656 233232
rect 559708 233220 559714 233232
rect 580166 233220 580172 233232
rect 559708 233192 580172 233220
rect 559708 233180 559714 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 442442 229984 442448 230036
rect 442500 230024 442506 230036
rect 443914 230024 443920 230036
rect 442500 229996 443920 230024
rect 442500 229984 442506 229996
rect 443914 229984 443920 229996
rect 443972 229984 443978 230036
rect 421558 229712 421564 229764
rect 421616 229752 421622 229764
rect 427078 229752 427084 229764
rect 421616 229724 427084 229752
rect 421616 229712 421622 229724
rect 427078 229712 427084 229724
rect 427136 229712 427142 229764
rect 361758 227672 361764 227724
rect 361816 227712 361822 227724
rect 443638 227712 443644 227724
rect 361816 227684 443644 227712
rect 361816 227672 361822 227684
rect 443638 227672 443644 227684
rect 443696 227672 443702 227724
rect 440878 226584 440884 226636
rect 440936 226624 440942 226636
rect 442442 226624 442448 226636
rect 440936 226596 442448 226624
rect 440936 226584 440942 226596
rect 442442 226584 442448 226596
rect 442500 226584 442506 226636
rect 450538 221416 450544 221468
rect 450596 221456 450602 221468
rect 457898 221456 457904 221468
rect 450596 221428 457904 221456
rect 450596 221416 450602 221428
rect 457898 221416 457904 221428
rect 457956 221416 457962 221468
rect 361666 216316 361672 216368
rect 361724 216356 361730 216368
rect 364058 216356 364064 216368
rect 361724 216328 364064 216356
rect 361724 216316 361730 216328
rect 364058 216316 364064 216328
rect 364116 216316 364122 216368
rect 439682 213868 439688 213920
rect 439740 213908 439746 213920
rect 440878 213908 440884 213920
rect 439740 213880 440884 213908
rect 439740 213868 439746 213880
rect 440878 213868 440884 213880
rect 440936 213868 440942 213920
rect 437474 208360 437480 208412
rect 437532 208400 437538 208412
rect 439682 208400 439688 208412
rect 437532 208372 439688 208400
rect 437532 208360 437538 208372
rect 439682 208360 439688 208372
rect 439740 208360 439746 208412
rect 450630 207612 450636 207664
rect 450688 207652 450694 207664
rect 459554 207652 459560 207664
rect 450688 207624 459560 207652
rect 450688 207612 450694 207624
rect 459554 207612 459560 207624
rect 459612 207652 459618 207664
rect 460014 207652 460020 207664
rect 459612 207624 460020 207652
rect 459612 207612 459618 207624
rect 460014 207612 460020 207624
rect 460072 207612 460078 207664
rect 576118 206932 576124 206984
rect 576176 206972 576182 206984
rect 579798 206972 579804 206984
rect 576176 206944 579804 206972
rect 576176 206932 576182 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 361758 205572 361764 205624
rect 361816 205612 361822 205624
rect 439590 205612 439596 205624
rect 361816 205584 439596 205612
rect 361816 205572 361822 205584
rect 439590 205572 439596 205584
rect 439648 205572 439654 205624
rect 3878 205096 3884 205148
rect 3936 205136 3942 205148
rect 5166 205136 5172 205148
rect 3936 205108 5172 205136
rect 3936 205096 3942 205108
rect 5166 205096 5172 205108
rect 5224 205096 5230 205148
rect 440878 204212 440884 204264
rect 440936 204252 440942 204264
rect 442258 204252 442264 204264
rect 440936 204224 442264 204252
rect 440936 204212 440942 204224
rect 442258 204212 442264 204224
rect 442316 204212 442322 204264
rect 410518 203396 410524 203448
rect 410576 203436 410582 203448
rect 414658 203436 414664 203448
rect 410576 203408 414664 203436
rect 410576 203396 410582 203408
rect 414658 203396 414664 203408
rect 414716 203396 414722 203448
rect 437474 202892 437480 202904
rect 436112 202864 437480 202892
rect 433334 202784 433340 202836
rect 433392 202824 433398 202836
rect 436112 202824 436140 202864
rect 437474 202852 437480 202864
rect 437532 202852 437538 202904
rect 433392 202796 436140 202824
rect 433392 202784 433398 202796
rect 447778 201288 447784 201340
rect 447836 201328 447842 201340
rect 449158 201328 449164 201340
rect 447836 201300 449164 201328
rect 447836 201288 447842 201300
rect 449158 201288 449164 201300
rect 449216 201288 449222 201340
rect 460658 200676 460664 200728
rect 460716 200716 460722 200728
rect 462314 200716 462320 200728
rect 460716 200688 462320 200716
rect 460716 200676 460722 200688
rect 462314 200676 462320 200688
rect 462372 200676 462378 200728
rect 447318 199384 447324 199436
rect 447376 199424 447382 199436
rect 461578 199424 461584 199436
rect 447376 199396 461584 199424
rect 447376 199384 447382 199396
rect 461578 199384 461584 199396
rect 461636 199384 461642 199436
rect 361758 194488 361764 194540
rect 361816 194528 361822 194540
rect 436738 194528 436744 194540
rect 361816 194500 436744 194528
rect 361816 194488 361822 194500
rect 436738 194488 436744 194500
rect 436796 194488 436802 194540
rect 418522 193128 418528 193180
rect 418580 193168 418586 193180
rect 421558 193168 421564 193180
rect 418580 193140 421564 193168
rect 418580 193128 418586 193140
rect 421558 193128 421564 193140
rect 421616 193128 421622 193180
rect 548518 193128 548524 193180
rect 548576 193168 548582 193180
rect 580166 193168 580172 193180
rect 548576 193140 580172 193168
rect 548576 193128 548582 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 439590 191768 439596 191820
rect 439648 191808 439654 191820
rect 440878 191808 440884 191820
rect 439648 191780 440884 191808
rect 439648 191768 439654 191780
rect 440878 191768 440884 191780
rect 440936 191768 440942 191820
rect 431218 190476 431224 190528
rect 431276 190516 431282 190528
rect 433242 190516 433248 190528
rect 431276 190488 433248 190516
rect 431276 190476 431282 190488
rect 433242 190476 433248 190488
rect 433300 190476 433306 190528
rect 407022 186940 407028 186992
rect 407080 186980 407086 186992
rect 418522 186980 418528 186992
rect 407080 186952 418528 186980
rect 407080 186940 407086 186952
rect 418522 186940 418528 186952
rect 418580 186940 418586 186992
rect 395338 184152 395344 184204
rect 395396 184192 395402 184204
rect 407022 184192 407028 184204
rect 395396 184164 407028 184192
rect 395396 184152 395402 184164
rect 407022 184152 407028 184164
rect 407080 184152 407086 184204
rect 361758 183472 361764 183524
rect 361816 183512 361822 183524
rect 447226 183512 447232 183524
rect 361816 183484 447232 183512
rect 361816 183472 361822 183484
rect 447226 183472 447232 183484
rect 447284 183472 447290 183524
rect 447226 182792 447232 182844
rect 447284 182832 447290 182844
rect 448146 182832 448152 182844
rect 447284 182804 448152 182832
rect 447284 182792 447290 182804
rect 448146 182792 448152 182804
rect 448204 182832 448210 182844
rect 528554 182832 528560 182844
rect 448204 182804 528560 182832
rect 448204 182792 448210 182804
rect 528554 182792 528560 182804
rect 528612 182792 528618 182844
rect 559558 179324 559564 179376
rect 559616 179364 559622 179376
rect 580166 179364 580172 179376
rect 559616 179336 580172 179364
rect 559616 179324 559622 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 419534 175924 419540 175976
rect 419592 175964 419598 175976
rect 431218 175964 431224 175976
rect 419592 175936 431224 175964
rect 419592 175924 419598 175936
rect 431218 175924 431224 175936
rect 431276 175924 431282 175976
rect 439590 175284 439596 175296
rect 437492 175256 439596 175284
rect 436738 175176 436744 175228
rect 436796 175216 436802 175228
rect 437492 175216 437520 175256
rect 439590 175244 439596 175256
rect 439648 175244 439654 175296
rect 436796 175188 437520 175216
rect 436796 175176 436802 175188
rect 389818 174564 389824 174616
rect 389876 174604 389882 174616
rect 395338 174604 395344 174616
rect 389876 174576 395344 174604
rect 389876 174564 389882 174576
rect 395338 174564 395344 174576
rect 395396 174564 395402 174616
rect 414658 173884 414664 173936
rect 414716 173924 414722 173936
rect 419534 173924 419540 173936
rect 414716 173896 419540 173924
rect 414716 173884 414722 173896
rect 419534 173884 419540 173896
rect 419592 173884 419598 173936
rect 361758 172456 361764 172508
rect 361816 172496 361822 172508
rect 447226 172496 447232 172508
rect 361816 172468 447232 172496
rect 361816 172456 361822 172468
rect 447226 172456 447232 172468
rect 447284 172456 447290 172508
rect 447226 171776 447232 171828
rect 447284 171816 447290 171828
rect 448330 171816 448336 171828
rect 447284 171788 448336 171816
rect 447284 171776 447290 171788
rect 448330 171776 448336 171788
rect 448388 171816 448394 171828
rect 524414 171816 524420 171828
rect 448388 171788 524420 171816
rect 448388 171776 448394 171788
rect 524414 171776 524420 171788
rect 524472 171776 524478 171828
rect 414658 169776 414664 169788
rect 412606 169748 414664 169776
rect 411254 169668 411260 169720
rect 411312 169708 411318 169720
rect 412606 169708 412634 169748
rect 414658 169736 414664 169748
rect 414716 169736 414722 169788
rect 432230 169736 432236 169788
rect 432288 169776 432294 169788
rect 436738 169776 436744 169788
rect 432288 169748 436744 169776
rect 432288 169736 432294 169748
rect 436738 169736 436744 169748
rect 436796 169736 436802 169788
rect 444006 169736 444012 169788
rect 444064 169776 444070 169788
rect 447778 169776 447784 169788
rect 444064 169748 447784 169776
rect 444064 169736 444070 169748
rect 447778 169736 447784 169748
rect 447836 169736 447842 169788
rect 411312 169680 412634 169708
rect 411312 169668 411318 169680
rect 432230 168416 432236 168428
rect 431926 168388 432236 168416
rect 429838 168308 429844 168360
rect 429896 168348 429902 168360
rect 431926 168348 431954 168388
rect 432230 168376 432236 168388
rect 432288 168376 432294 168428
rect 429896 168320 431954 168348
rect 429896 168308 429902 168320
rect 536098 166948 536104 167000
rect 536156 166988 536162 167000
rect 580166 166988 580172 167000
rect 536156 166960 580172 166988
rect 536156 166948 536162 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 369026 166268 369032 166320
rect 369084 166308 369090 166320
rect 389818 166308 389824 166320
rect 369084 166280 389824 166308
rect 369084 166268 369090 166280
rect 389818 166268 389824 166280
rect 389876 166268 389882 166320
rect 440234 165928 440240 165980
rect 440292 165968 440298 165980
rect 444006 165968 444012 165980
rect 440292 165940 444012 165968
rect 440292 165928 440298 165940
rect 444006 165928 444012 165940
rect 444064 165928 444070 165980
rect 411254 164268 411260 164280
rect 409892 164240 411260 164268
rect 408494 164160 408500 164212
rect 408552 164200 408558 164212
rect 409892 164200 409920 164240
rect 411254 164228 411260 164240
rect 411312 164228 411318 164280
rect 408552 164172 409920 164200
rect 408552 164160 408558 164172
rect 448422 164160 448428 164212
rect 448480 164200 448486 164212
rect 449342 164200 449348 164212
rect 448480 164172 449348 164200
rect 448480 164160 448486 164172
rect 449342 164160 449348 164172
rect 449400 164160 449406 164212
rect 438578 163616 438584 163668
rect 438636 163656 438642 163668
rect 439498 163656 439504 163668
rect 438636 163628 439504 163656
rect 438636 163616 438642 163628
rect 439498 163616 439504 163628
rect 439556 163616 439562 163668
rect 445202 163616 445208 163668
rect 445260 163656 445266 163668
rect 446398 163656 446404 163668
rect 445260 163628 446404 163656
rect 445260 163616 445266 163628
rect 446398 163616 446404 163628
rect 446456 163616 446462 163668
rect 361574 163480 361580 163532
rect 361632 163520 361638 163532
rect 369026 163520 369032 163532
rect 361632 163492 369032 163520
rect 361632 163480 361638 163492
rect 369026 163480 369032 163492
rect 369084 163480 369090 163532
rect 437566 162256 437572 162308
rect 437624 162296 437630 162308
rect 440234 162296 440240 162308
rect 437624 162268 440240 162296
rect 437624 162256 437630 162268
rect 440234 162256 440240 162268
rect 440292 162256 440298 162308
rect 418706 162188 418712 162240
rect 418764 162228 418770 162240
rect 457806 162228 457812 162240
rect 418764 162200 457812 162228
rect 418764 162188 418770 162200
rect 457806 162188 457812 162200
rect 457864 162228 457870 162240
rect 489914 162228 489920 162240
rect 457864 162200 489920 162228
rect 457864 162188 457870 162200
rect 489914 162188 489920 162200
rect 489972 162188 489978 162240
rect 415118 162120 415124 162172
rect 415176 162160 415182 162172
rect 457898 162160 457904 162172
rect 415176 162132 457904 162160
rect 415176 162120 415182 162132
rect 457898 162120 457904 162132
rect 457956 162160 457962 162172
rect 485774 162160 485780 162172
rect 457956 162132 485780 162160
rect 457956 162120 457962 162132
rect 485774 162120 485780 162132
rect 485832 162120 485838 162172
rect 445202 161576 445208 161628
rect 445260 161616 445266 161628
rect 450538 161616 450544 161628
rect 445260 161588 450544 161616
rect 445260 161576 445266 161588
rect 450538 161576 450544 161588
rect 450596 161576 450602 161628
rect 375190 161508 375196 161560
rect 375248 161548 375254 161560
rect 418706 161548 418712 161560
rect 375248 161520 418712 161548
rect 375248 161508 375254 161520
rect 418706 161508 418712 161520
rect 418764 161508 418770 161560
rect 431862 161508 431868 161560
rect 431920 161548 431926 161560
rect 450630 161548 450636 161560
rect 431920 161520 450636 161548
rect 431920 161508 431926 161520
rect 450630 161508 450636 161520
rect 450688 161508 450694 161560
rect 412082 161440 412088 161492
rect 412140 161480 412146 161492
rect 459554 161480 459560 161492
rect 412140 161452 459560 161480
rect 412140 161440 412146 161452
rect 459554 161440 459560 161452
rect 459612 161480 459618 161492
rect 460382 161480 460388 161492
rect 459612 161452 460388 161480
rect 459612 161440 459618 161452
rect 460382 161440 460388 161452
rect 460440 161440 460446 161492
rect 361758 161372 361764 161424
rect 361816 161412 361822 161424
rect 448330 161412 448336 161424
rect 361816 161384 448336 161412
rect 361816 161372 361822 161384
rect 448330 161372 448336 161384
rect 448388 161372 448394 161424
rect 448330 160692 448336 160744
rect 448388 160732 448394 160744
rect 521654 160732 521660 160744
rect 448388 160704 521660 160732
rect 448388 160692 448394 160704
rect 521654 160692 521660 160704
rect 521712 160692 521718 160744
rect 425330 160420 425336 160472
rect 425388 160460 425394 160472
rect 425882 160460 425888 160472
rect 425388 160432 425888 160460
rect 425388 160420 425394 160432
rect 425882 160420 425888 160432
rect 425940 160460 425946 160472
rect 496814 160460 496820 160472
rect 425940 160432 496820 160460
rect 425940 160420 425946 160432
rect 496814 160420 496820 160432
rect 496872 160420 496878 160472
rect 428642 160352 428648 160404
rect 428700 160392 428706 160404
rect 500954 160392 500960 160404
rect 428700 160364 500960 160392
rect 428700 160352 428706 160364
rect 500954 160352 500960 160364
rect 501012 160352 501018 160404
rect 421834 160284 421840 160336
rect 421892 160324 421898 160336
rect 494054 160324 494060 160336
rect 421892 160296 494060 160324
rect 421892 160284 421898 160296
rect 494054 160284 494060 160296
rect 494112 160284 494118 160336
rect 435266 160216 435272 160268
rect 435324 160256 435330 160268
rect 436002 160256 436008 160268
rect 435324 160228 436008 160256
rect 435324 160216 435330 160228
rect 436002 160216 436008 160228
rect 436060 160256 436066 160268
rect 509234 160256 509240 160268
rect 436060 160228 509240 160256
rect 436060 160216 436066 160228
rect 509234 160216 509240 160228
rect 509292 160216 509298 160268
rect 386138 160148 386144 160200
rect 386196 160188 386202 160200
rect 415118 160188 415124 160200
rect 386196 160160 415124 160188
rect 386196 160148 386202 160160
rect 415118 160148 415124 160160
rect 415176 160148 415182 160200
rect 427814 160148 427820 160200
rect 427872 160188 427878 160200
rect 429838 160188 429844 160200
rect 427872 160160 429844 160188
rect 427872 160148 427878 160160
rect 429838 160148 429844 160160
rect 429896 160148 429902 160200
rect 438578 160148 438584 160200
rect 438636 160188 438642 160200
rect 513374 160188 513380 160200
rect 438636 160160 513380 160188
rect 438636 160148 438642 160160
rect 513374 160148 513380 160160
rect 513432 160148 513438 160200
rect 409506 160080 409512 160132
rect 409564 160120 409570 160132
rect 441568 160120 441574 160132
rect 409564 160092 441574 160120
rect 409564 160080 409570 160092
rect 441568 160080 441574 160092
rect 441626 160120 441632 160132
rect 442902 160120 442908 160132
rect 441626 160092 442908 160120
rect 441626 160080 441632 160092
rect 442902 160080 442908 160092
rect 442960 160120 442966 160132
rect 517514 160120 517520 160132
rect 442960 160092 517520 160120
rect 442960 160080 442966 160092
rect 517514 160080 517520 160092
rect 517572 160080 517578 160132
rect 401594 159808 401600 159860
rect 401652 159848 401658 159860
rect 408494 159848 408500 159860
rect 401652 159820 408500 159848
rect 401652 159808 401658 159820
rect 408494 159808 408500 159820
rect 408552 159808 408558 159860
rect 409414 159740 409420 159792
rect 409472 159780 409478 159792
rect 427814 159780 427820 159792
rect 409472 159752 427820 159780
rect 409472 159740 409478 159752
rect 427814 159740 427820 159752
rect 427872 159740 427878 159792
rect 409138 159672 409144 159724
rect 409196 159712 409202 159724
rect 427998 159712 428004 159724
rect 409196 159684 428004 159712
rect 409196 159672 409202 159684
rect 427998 159672 428004 159684
rect 428056 159672 428062 159724
rect 409230 159604 409236 159656
rect 409288 159644 409294 159656
rect 434806 159644 434812 159656
rect 409288 159616 434812 159644
rect 409288 159604 409294 159616
rect 434806 159604 434812 159616
rect 434864 159604 434870 159656
rect 409322 159536 409328 159588
rect 409380 159576 409386 159588
rect 437934 159576 437940 159588
rect 409380 159548 437940 159576
rect 409380 159536 409386 159548
rect 437934 159536 437940 159548
rect 437992 159536 437998 159588
rect 406102 159468 406108 159520
rect 406160 159508 406166 159520
rect 437566 159508 437572 159520
rect 406160 159480 437572 159508
rect 406160 159468 406166 159480
rect 437566 159468 437572 159480
rect 437624 159468 437630 159520
rect 384206 159400 384212 159452
rect 384264 159440 384270 159452
rect 421374 159440 421380 159452
rect 384264 159412 421380 159440
rect 384264 159400 384270 159412
rect 421374 159400 421380 159412
rect 421432 159400 421438 159452
rect 386230 159332 386236 159384
rect 386288 159372 386294 159384
rect 425146 159372 425152 159384
rect 386288 159344 425152 159372
rect 386288 159332 386294 159344
rect 425146 159332 425152 159344
rect 425204 159332 425210 159384
rect 451734 158244 451740 158296
rect 451792 158284 451798 158296
rect 456150 158284 456156 158296
rect 451792 158256 456156 158284
rect 451792 158244 451798 158256
rect 456150 158244 456156 158256
rect 456208 158244 456214 158296
rect 404262 157496 404268 157548
rect 404320 157536 404326 157548
rect 406102 157536 406108 157548
rect 404320 157508 406108 157536
rect 404320 157496 404326 157508
rect 406102 157496 406108 157508
rect 406160 157496 406166 157548
rect 451734 157292 451740 157344
rect 451792 157332 451798 157344
rect 457530 157332 457536 157344
rect 451792 157304 457536 157332
rect 451792 157292 451798 157304
rect 457530 157292 457536 157304
rect 457588 157292 457594 157344
rect 400858 156612 400864 156664
rect 400916 156652 400922 156664
rect 410518 156652 410524 156664
rect 400916 156624 410524 156652
rect 400916 156612 400922 156624
rect 410518 156612 410524 156624
rect 410576 156612 410582 156664
rect 396718 156136 396724 156188
rect 396776 156176 396782 156188
rect 404262 156176 404268 156188
rect 396776 156148 404268 156176
rect 396776 156136 396782 156148
rect 404262 156136 404268 156148
rect 404320 156136 404326 156188
rect 359458 155320 359464 155372
rect 359516 155360 359522 155372
rect 361574 155360 361580 155372
rect 359516 155332 361580 155360
rect 359516 155320 359522 155332
rect 361574 155320 361580 155332
rect 361632 155320 361638 155372
rect 451918 154164 451924 154216
rect 451976 154204 451982 154216
rect 455230 154204 455236 154216
rect 451976 154176 455236 154204
rect 451976 154164 451982 154176
rect 455230 154164 455236 154176
rect 455288 154164 455294 154216
rect 401594 153252 401600 153264
rect 398852 153224 401600 153252
rect 396902 153144 396908 153196
rect 396960 153184 396966 153196
rect 398852 153184 398880 153224
rect 401594 153212 401600 153224
rect 401652 153212 401658 153264
rect 396960 153156 398880 153184
rect 396960 153144 396966 153156
rect 547138 153144 547144 153196
rect 547196 153184 547202 153196
rect 580166 153184 580172 153196
rect 547196 153156 580172 153184
rect 547196 153144 547202 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 395154 150424 395160 150476
rect 395212 150464 395218 150476
rect 396902 150464 396908 150476
rect 395212 150436 396908 150464
rect 395212 150424 395218 150436
rect 396902 150424 396908 150436
rect 396960 150424 396966 150476
rect 361758 150356 361764 150408
rect 361816 150396 361822 150408
rect 409506 150396 409512 150408
rect 361816 150368 409512 150396
rect 361816 150356 361822 150368
rect 409506 150356 409512 150368
rect 409564 150356 409570 150408
rect 452470 150220 452476 150272
rect 452528 150260 452534 150272
rect 459278 150260 459284 150272
rect 452528 150232 459284 150260
rect 452528 150220 452534 150232
rect 459278 150220 459284 150232
rect 459336 150220 459342 150272
rect 452562 148724 452568 148776
rect 452620 148764 452626 148776
rect 454954 148764 454960 148776
rect 452620 148736 454960 148764
rect 452620 148724 452626 148736
rect 454954 148724 454960 148736
rect 455012 148724 455018 148776
rect 391198 147636 391204 147688
rect 391256 147676 391262 147688
rect 395154 147676 395160 147688
rect 391256 147648 395160 147676
rect 391256 147636 391262 147648
rect 395154 147636 395160 147648
rect 395212 147636 395218 147688
rect 407114 147636 407120 147688
rect 407172 147676 407178 147688
rect 409414 147676 409420 147688
rect 407172 147648 409420 147676
rect 407172 147636 407178 147648
rect 409414 147636 409420 147648
rect 409472 147636 409478 147688
rect 451734 147364 451740 147416
rect 451792 147404 451798 147416
rect 457714 147404 457720 147416
rect 451792 147376 457720 147404
rect 451792 147364 451798 147376
rect 457714 147364 457720 147376
rect 457772 147364 457778 147416
rect 452562 146004 452568 146056
rect 452620 146044 452626 146056
rect 459002 146044 459008 146056
rect 452620 146016 459008 146044
rect 452620 146004 452626 146016
rect 459002 146004 459008 146016
rect 459060 146004 459066 146056
rect 396810 145120 396816 145172
rect 396868 145160 396874 145172
rect 400858 145160 400864 145172
rect 396868 145132 400864 145160
rect 396868 145120 396874 145132
rect 400858 145120 400864 145132
rect 400916 145120 400922 145172
rect 404814 145120 404820 145172
rect 404872 145160 404878 145172
rect 407114 145160 407120 145172
rect 404872 145132 407120 145160
rect 404872 145120 404878 145132
rect 407114 145120 407120 145132
rect 407172 145120 407178 145172
rect 451458 144780 451464 144832
rect 451516 144820 451522 144832
rect 455046 144820 455052 144832
rect 451516 144792 455052 144820
rect 451516 144780 451522 144792
rect 455046 144780 455052 144792
rect 455104 144780 455110 144832
rect 460382 143488 460388 143540
rect 460440 143528 460446 143540
rect 460842 143528 460848 143540
rect 460440 143500 460848 143528
rect 460440 143488 460446 143500
rect 460842 143488 460848 143500
rect 460900 143488 460906 143540
rect 533430 143488 533436 143540
rect 533488 143528 533494 143540
rect 537294 143528 537300 143540
rect 533488 143500 537300 143528
rect 533488 143488 533494 143500
rect 537294 143488 537300 143500
rect 537352 143488 537358 143540
rect 452562 143284 452568 143336
rect 452620 143324 452626 143336
rect 459186 143324 459192 143336
rect 452620 143296 459192 143324
rect 452620 143284 452626 143296
rect 459186 143284 459192 143296
rect 459244 143284 459250 143336
rect 460842 142264 460848 142316
rect 460900 142304 460906 142316
rect 481910 142304 481916 142316
rect 460900 142276 481916 142304
rect 460900 142264 460906 142276
rect 481910 142264 481916 142276
rect 481968 142264 481974 142316
rect 450630 142196 450636 142248
rect 450688 142236 450694 142248
rect 505646 142236 505652 142248
rect 450688 142208 505652 142236
rect 450688 142196 450694 142208
rect 505646 142196 505652 142208
rect 505704 142196 505710 142248
rect 540330 142236 540336 142248
rect 538186 142208 540336 142236
rect 401594 142128 401600 142180
rect 401652 142168 401658 142180
rect 404814 142168 404820 142180
rect 401652 142140 404820 142168
rect 401652 142128 401658 142140
rect 404814 142128 404820 142140
rect 404872 142128 404878 142180
rect 450538 142128 450544 142180
rect 450596 142168 450602 142180
rect 533982 142168 533988 142180
rect 450596 142140 533988 142168
rect 450596 142128 450602 142140
rect 533982 142128 533988 142140
rect 534040 142168 534046 142180
rect 538186 142168 538214 142208
rect 540330 142196 540336 142208
rect 540388 142196 540394 142248
rect 534040 142140 538214 142168
rect 534040 142128 534046 142140
rect 452562 141924 452568 141976
rect 452620 141964 452626 141976
rect 455138 141964 455144 141976
rect 452620 141936 455144 141964
rect 452620 141924 452626 141936
rect 455138 141924 455144 141936
rect 455196 141924 455202 141976
rect 452562 140564 452568 140616
rect 452620 140604 452626 140616
rect 457622 140604 457628 140616
rect 452620 140576 457628 140604
rect 452620 140564 452626 140576
rect 457622 140564 457628 140576
rect 457680 140564 457686 140616
rect 534718 140088 534724 140140
rect 534776 140128 534782 140140
rect 542906 140128 542912 140140
rect 534776 140100 542912 140128
rect 534776 140088 534782 140100
rect 542906 140088 542912 140100
rect 542964 140088 542970 140140
rect 533338 140020 533344 140072
rect 533396 140060 533402 140072
rect 543182 140060 543188 140072
rect 533396 140032 543188 140060
rect 533396 140020 533402 140032
rect 543182 140020 543188 140032
rect 543240 140020 543246 140072
rect 361758 139340 361764 139392
rect 361816 139380 361822 139392
rect 409322 139380 409328 139392
rect 361816 139352 409328 139380
rect 361816 139340 361822 139352
rect 409322 139340 409328 139352
rect 409380 139340 409386 139392
rect 555418 139340 555424 139392
rect 555476 139380 555482 139392
rect 580166 139380 580172 139392
rect 555476 139352 580172 139380
rect 555476 139340 555482 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 452562 139204 452568 139256
rect 452620 139244 452626 139256
rect 459094 139244 459100 139256
rect 452620 139216 459100 139244
rect 452620 139204 452626 139216
rect 459094 139204 459100 139216
rect 459152 139204 459158 139256
rect 538858 138592 538864 138644
rect 538916 138632 538922 138644
rect 543090 138632 543096 138644
rect 538916 138604 543096 138632
rect 538916 138592 538922 138604
rect 543090 138592 543096 138604
rect 543148 138592 543154 138644
rect 452562 137844 452568 137896
rect 452620 137884 452626 137896
rect 454770 137884 454776 137896
rect 452620 137856 454776 137884
rect 452620 137844 452626 137856
rect 454770 137844 454776 137856
rect 454828 137844 454834 137896
rect 389450 137300 389456 137352
rect 389508 137340 389514 137352
rect 391198 137340 391204 137352
rect 389508 137312 391204 137340
rect 389508 137300 389514 137312
rect 391198 137300 391204 137312
rect 391256 137300 391262 137352
rect 388438 137232 388444 137284
rect 388496 137272 388502 137284
rect 396810 137272 396816 137284
rect 388496 137244 396816 137272
rect 388496 137232 388502 137244
rect 396810 137232 396816 137244
rect 396868 137232 396874 137284
rect 394694 136620 394700 136672
rect 394752 136660 394758 136672
rect 396718 136660 396724 136672
rect 394752 136632 396724 136660
rect 394752 136620 394758 136632
rect 396718 136620 396724 136632
rect 396776 136620 396782 136672
rect 538950 136552 538956 136604
rect 539008 136592 539014 136604
rect 539502 136592 539508 136604
rect 539008 136564 539508 136592
rect 539008 136552 539014 136564
rect 539502 136552 539508 136564
rect 539560 136552 539566 136604
rect 452562 136484 452568 136536
rect 452620 136524 452626 136536
rect 457438 136524 457444 136536
rect 452620 136496 457444 136524
rect 452620 136484 452626 136496
rect 457438 136484 457444 136496
rect 457496 136484 457502 136536
rect 391198 135872 391204 135924
rect 391256 135912 391262 135924
rect 401502 135912 401508 135924
rect 391256 135884 401508 135912
rect 391256 135872 391262 135884
rect 401502 135872 401508 135884
rect 401560 135872 401566 135924
rect 387794 135192 387800 135244
rect 387852 135232 387858 135244
rect 389450 135232 389456 135244
rect 387852 135204 389456 135232
rect 387852 135192 387858 135204
rect 389450 135192 389456 135204
rect 389508 135192 389514 135244
rect 452562 135124 452568 135176
rect 452620 135164 452626 135176
rect 458910 135164 458916 135176
rect 452620 135136 458916 135164
rect 452620 135124 452626 135136
rect 458910 135124 458916 135136
rect 458968 135124 458974 135176
rect 452562 133764 452568 133816
rect 452620 133804 452626 133816
rect 454862 133804 454868 133816
rect 452620 133776 454868 133804
rect 452620 133764 452626 133776
rect 454862 133764 454868 133776
rect 454920 133764 454926 133816
rect 394694 132512 394700 132524
rect 393332 132484 394700 132512
rect 391934 132404 391940 132456
rect 391992 132444 391998 132456
rect 393332 132444 393360 132484
rect 394694 132472 394700 132484
rect 394752 132472 394758 132524
rect 391992 132416 393360 132444
rect 391992 132404 391998 132416
rect 452286 131044 452292 131096
rect 452344 131084 452350 131096
rect 453390 131084 453396 131096
rect 452344 131056 453396 131084
rect 452344 131044 452350 131056
rect 453390 131044 453396 131056
rect 453448 131044 453454 131096
rect 389174 129820 389180 129872
rect 389232 129860 389238 129872
rect 391198 129860 391204 129872
rect 389232 129832 391204 129860
rect 389232 129820 389238 129832
rect 391198 129820 391204 129832
rect 391256 129820 391262 129872
rect 387058 129752 387064 129804
rect 387116 129792 387122 129804
rect 391934 129792 391940 129804
rect 387116 129764 391940 129792
rect 387116 129752 387122 129764
rect 391934 129752 391940 129764
rect 391992 129752 391998 129804
rect 452378 129684 452384 129736
rect 452436 129724 452442 129736
rect 453482 129724 453488 129736
rect 452436 129696 453488 129724
rect 452436 129684 452442 129696
rect 453482 129684 453488 129696
rect 453540 129684 453546 129736
rect 359550 129004 359556 129056
rect 359608 129044 359614 129056
rect 388438 129044 388444 129056
rect 359608 129016 388444 129044
rect 359608 129004 359614 129016
rect 388438 129004 388444 129016
rect 388496 129004 388502 129056
rect 361758 128256 361764 128308
rect 361816 128296 361822 128308
rect 409230 128296 409236 128308
rect 361816 128268 409236 128296
rect 361816 128256 361822 128268
rect 409230 128256 409236 128268
rect 409288 128256 409294 128308
rect 452286 126896 452292 126948
rect 452344 126936 452350 126948
rect 453298 126936 453304 126948
rect 452344 126908 453304 126936
rect 452344 126896 452350 126908
rect 453298 126896 453304 126908
rect 453356 126896 453362 126948
rect 573358 126896 573364 126948
rect 573416 126936 573422 126948
rect 580166 126936 580172 126948
rect 573416 126908 580172 126936
rect 573416 126896 573422 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 451734 126352 451740 126404
rect 451792 126392 451798 126404
rect 453574 126392 453580 126404
rect 451792 126364 453580 126392
rect 451792 126352 451798 126364
rect 453574 126352 453580 126364
rect 453632 126352 453638 126404
rect 368290 126216 368296 126268
rect 368348 126256 368354 126268
rect 387702 126256 387708 126268
rect 368348 126228 387708 126256
rect 368348 126216 368354 126228
rect 387702 126216 387708 126228
rect 387760 126216 387766 126268
rect 362954 124856 362960 124908
rect 363012 124896 363018 124908
rect 389082 124896 389088 124908
rect 363012 124868 389088 124896
rect 363012 124856 363018 124868
rect 389082 124856 389088 124868
rect 389140 124856 389146 124908
rect 451826 124108 451832 124160
rect 451884 124148 451890 124160
rect 458818 124148 458824 124160
rect 451884 124120 458824 124148
rect 451884 124108 451890 124120
rect 458818 124108 458824 124120
rect 458876 124108 458882 124160
rect 451734 122204 451740 122256
rect 451792 122244 451798 122256
rect 454678 122244 454684 122256
rect 451792 122216 454684 122244
rect 451792 122204 451798 122216
rect 454678 122204 454684 122216
rect 454736 122204 454742 122256
rect 371234 122068 371240 122120
rect 371292 122108 371298 122120
rect 387058 122108 387064 122120
rect 371292 122080 387064 122108
rect 371292 122068 371298 122080
rect 387058 122068 387064 122080
rect 387116 122068 387122 122120
rect 384942 119348 384948 119400
rect 385000 119388 385006 119400
rect 456058 119388 456064 119400
rect 385000 119360 456064 119388
rect 385000 119348 385006 119360
rect 456058 119348 456064 119360
rect 456116 119348 456122 119400
rect 361298 118668 361304 118720
rect 361356 118708 361362 118720
rect 362862 118708 362868 118720
rect 361356 118680 362868 118708
rect 361356 118668 361362 118680
rect 362862 118668 362868 118680
rect 362920 118668 362926 118720
rect 371234 118708 371240 118720
rect 369872 118680 371240 118708
rect 366910 118600 366916 118652
rect 366968 118640 366974 118652
rect 369872 118640 369900 118680
rect 371234 118668 371240 118680
rect 371292 118668 371298 118720
rect 366968 118612 369900 118640
rect 366968 118600 366974 118612
rect 362586 117920 362592 117972
rect 362644 117960 362650 117972
rect 368290 117960 368296 117972
rect 362644 117932 368296 117960
rect 362644 117920 362650 117932
rect 368290 117920 368296 117932
rect 368348 117920 368354 117972
rect 361758 117240 361764 117292
rect 361816 117280 361822 117292
rect 450630 117280 450636 117292
rect 361816 117252 450636 117280
rect 361816 117240 361822 117252
rect 450630 117240 450636 117252
rect 450688 117240 450694 117292
rect 364058 116832 364064 116884
rect 364116 116872 364122 116884
rect 366910 116872 366916 116884
rect 364116 116844 366916 116872
rect 364116 116832 364122 116844
rect 366910 116832 366916 116844
rect 366968 116832 366974 116884
rect 569218 113092 569224 113144
rect 569276 113132 569282 113144
rect 579798 113132 579804 113144
rect 569276 113104 579804 113132
rect 569276 113092 569282 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 361390 111800 361396 111852
rect 361448 111840 361454 111852
rect 364058 111840 364064 111852
rect 361448 111812 364064 111840
rect 361448 111800 361454 111812
rect 364058 111800 364064 111812
rect 364116 111800 364122 111852
rect 389818 106904 389824 106956
rect 389876 106944 389882 106956
rect 450538 106944 450544 106956
rect 389876 106916 450544 106944
rect 389876 106904 389882 106916
rect 450538 106904 450544 106916
rect 450596 106904 450602 106956
rect 361758 106224 361764 106276
rect 361816 106264 361822 106276
rect 409138 106264 409144 106276
rect 361816 106236 409144 106264
rect 361816 106224 361822 106236
rect 409138 106224 409144 106236
rect 409196 106224 409202 106276
rect 558178 100648 558184 100700
rect 558236 100688 558242 100700
rect 580166 100688 580172 100700
rect 558236 100660 580172 100688
rect 558236 100648 558242 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 361758 95140 361764 95192
rect 361816 95180 361822 95192
rect 386230 95180 386236 95192
rect 361816 95152 386236 95180
rect 361816 95140 361822 95152
rect 386230 95140 386236 95152
rect 386288 95140 386294 95192
rect 571978 86912 571984 86964
rect 572036 86952 572042 86964
rect 580166 86952 580172 86964
rect 572036 86924 580172 86952
rect 572036 86912 572042 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3142 84192 3148 84244
rect 3200 84232 3206 84244
rect 20898 84232 20904 84244
rect 3200 84204 20904 84232
rect 3200 84192 3206 84204
rect 20898 84192 20904 84204
rect 20956 84192 20962 84244
rect 361758 84124 361764 84176
rect 361816 84164 361822 84176
rect 384206 84164 384212 84176
rect 361816 84136 384212 84164
rect 361816 84124 361822 84136
rect 384206 84124 384212 84136
rect 384264 84124 384270 84176
rect 5074 80044 5080 80096
rect 5132 80084 5138 80096
rect 5132 80056 6914 80084
rect 5132 80044 5138 80056
rect 6886 80016 6914 80056
rect 8570 80016 8576 80028
rect 6886 79988 8576 80016
rect 8570 79976 8576 79988
rect 8628 79976 8634 80028
rect 8570 78480 8576 78532
rect 8628 78520 8634 78532
rect 10318 78520 10324 78532
rect 8628 78492 10324 78520
rect 8628 78480 8634 78492
rect 10318 78480 10324 78492
rect 10376 78480 10382 78532
rect 361758 73108 361764 73160
rect 361816 73148 361822 73160
rect 375190 73148 375196 73160
rect 361816 73120 375196 73148
rect 361816 73108 361822 73120
rect 375190 73108 375196 73120
rect 375248 73108 375254 73160
rect 544378 73108 544384 73160
rect 544436 73148 544442 73160
rect 580166 73148 580172 73160
rect 544436 73120 580172 73148
rect 544436 73108 544442 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3142 70388 3148 70440
rect 3200 70428 3206 70440
rect 20070 70428 20076 70440
rect 3200 70400 20076 70428
rect 3200 70388 3206 70400
rect 20070 70388 20076 70400
rect 20128 70388 20134 70440
rect 5166 68960 5172 69012
rect 5224 69000 5230 69012
rect 7558 69000 7564 69012
rect 5224 68972 7564 69000
rect 5224 68960 5230 68972
rect 7558 68960 7564 68972
rect 7616 68960 7622 69012
rect 4890 68892 4896 68944
rect 4948 68932 4954 68944
rect 5534 68932 5540 68944
rect 4948 68904 5540 68932
rect 4948 68892 4954 68904
rect 5534 68892 5540 68904
rect 5592 68892 5598 68944
rect 5534 66240 5540 66292
rect 5592 66280 5598 66292
rect 5592 66252 6914 66280
rect 5592 66240 5598 66252
rect 6886 66212 6914 66252
rect 8294 66212 8300 66224
rect 6886 66184 8300 66212
rect 8294 66172 8300 66184
rect 8352 66172 8358 66224
rect 10318 63860 10324 63912
rect 10376 63900 10382 63912
rect 12066 63900 12072 63912
rect 10376 63872 12072 63900
rect 10376 63860 10382 63872
rect 12066 63860 12072 63872
rect 12124 63860 12130 63912
rect 8294 62636 8300 62688
rect 8352 62676 8358 62688
rect 10410 62676 10416 62688
rect 8352 62648 10416 62676
rect 8352 62636 8358 62648
rect 10410 62636 10416 62648
rect 10468 62636 10474 62688
rect 361758 62024 361764 62076
rect 361816 62064 361822 62076
rect 386138 62064 386144 62076
rect 361816 62036 386144 62064
rect 361816 62024 361822 62036
rect 386138 62024 386144 62036
rect 386196 62024 386202 62076
rect 7558 60664 7564 60716
rect 7616 60704 7622 60716
rect 9582 60704 9588 60716
rect 7616 60676 9588 60704
rect 7616 60664 7622 60676
rect 9582 60664 9588 60676
rect 9640 60664 9646 60716
rect 551278 60664 551284 60716
rect 551336 60704 551342 60716
rect 580166 60704 580172 60716
rect 551336 60676 580172 60704
rect 551336 60664 551342 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3418 59984 3424 60036
rect 3476 60024 3482 60036
rect 20898 60024 20904 60036
rect 3476 59996 20904 60024
rect 3476 59984 3482 59996
rect 20898 59984 20904 59996
rect 20956 59984 20962 60036
rect 4798 59304 4804 59356
rect 4856 59344 4862 59356
rect 7558 59344 7564 59356
rect 4856 59316 7564 59344
rect 4856 59304 4862 59316
rect 7558 59304 7564 59316
rect 7616 59304 7622 59356
rect 4982 57876 4988 57928
rect 5040 57916 5046 57928
rect 5534 57916 5540 57928
rect 5040 57888 5540 57916
rect 5040 57876 5046 57888
rect 5534 57876 5540 57888
rect 5592 57876 5598 57928
rect 7558 56584 7564 56636
rect 7616 56624 7622 56636
rect 7616 56596 8340 56624
rect 7616 56584 7622 56596
rect 8312 56556 8340 56596
rect 10778 56556 10784 56568
rect 8312 56528 10784 56556
rect 10778 56516 10784 56528
rect 10836 56516 10842 56568
rect 12066 56516 12072 56568
rect 12124 56556 12130 56568
rect 13722 56556 13728 56568
rect 12124 56528 13728 56556
rect 12124 56516 12130 56528
rect 13722 56516 13728 56528
rect 13780 56516 13786 56568
rect 17954 56556 17960 56568
rect 16546 56528 17960 56556
rect 10410 56448 10416 56500
rect 10468 56488 10474 56500
rect 12434 56488 12440 56500
rect 10468 56460 12440 56488
rect 10468 56448 10474 56460
rect 12434 56448 12440 56460
rect 12492 56448 12498 56500
rect 9674 56380 9680 56432
rect 9732 56420 9738 56432
rect 16546 56420 16574 56528
rect 17954 56516 17960 56528
rect 18012 56516 18018 56568
rect 9732 56392 16574 56420
rect 9732 56380 9738 56392
rect 10778 54612 10784 54664
rect 10836 54652 10842 54664
rect 13630 54652 13636 54664
rect 10836 54624 13636 54652
rect 10836 54612 10842 54624
rect 13630 54612 13636 54624
rect 13688 54612 13694 54664
rect 5534 54476 5540 54528
rect 5592 54516 5598 54528
rect 11698 54516 11704 54528
rect 5592 54488 11704 54516
rect 5592 54476 5598 54488
rect 11698 54476 11704 54488
rect 11756 54476 11762 54528
rect 17954 54068 17960 54120
rect 18012 54108 18018 54120
rect 20622 54108 20628 54120
rect 18012 54080 20628 54108
rect 18012 54068 18018 54080
rect 20622 54068 20628 54080
rect 20680 54068 20686 54120
rect 13722 52980 13728 53032
rect 13780 53020 13786 53032
rect 15194 53020 15200 53032
rect 13780 52992 15200 53020
rect 13780 52980 13786 52992
rect 15194 52980 15200 52992
rect 15252 52980 15258 53032
rect 12434 52708 12440 52760
rect 12492 52748 12498 52760
rect 14550 52748 14556 52760
rect 12492 52720 14556 52748
rect 12492 52708 12498 52720
rect 14550 52708 14556 52720
rect 14608 52708 14614 52760
rect 13630 52436 13636 52488
rect 13688 52476 13694 52488
rect 13688 52448 13860 52476
rect 13688 52436 13694 52448
rect 13832 52408 13860 52448
rect 19242 52408 19248 52420
rect 13832 52380 19248 52408
rect 19242 52368 19248 52380
rect 19300 52368 19306 52420
rect 11698 51076 11704 51128
rect 11756 51116 11762 51128
rect 11756 51088 12480 51116
rect 11756 51076 11762 51088
rect 12452 51048 12480 51088
rect 361758 51076 361764 51128
rect 361816 51116 361822 51128
rect 386138 51116 386144 51128
rect 361816 51088 386144 51116
rect 361816 51076 361822 51088
rect 386138 51076 386144 51088
rect 386196 51076 386202 51128
rect 540606 51076 540612 51128
rect 540664 51116 540670 51128
rect 543734 51116 543740 51128
rect 540664 51088 543740 51116
rect 540664 51076 540670 51088
rect 543734 51076 543740 51088
rect 543792 51076 543798 51128
rect 15286 51048 15292 51060
rect 12452 51020 15292 51048
rect 15286 51008 15292 51020
rect 15344 51008 15350 51060
rect 15194 49648 15200 49700
rect 15252 49688 15258 49700
rect 16850 49688 16856 49700
rect 15252 49660 16856 49688
rect 15252 49648 15258 49660
rect 16850 49648 16856 49660
rect 16908 49648 16914 49700
rect 16850 48152 16856 48204
rect 16908 48192 16914 48204
rect 20806 48192 20812 48204
rect 16908 48164 20812 48192
rect 16908 48152 16914 48164
rect 20806 48152 20812 48164
rect 20864 48152 20870 48204
rect 15286 47268 15292 47320
rect 15344 47308 15350 47320
rect 19242 47308 19248 47320
rect 15344 47280 19248 47308
rect 15344 47268 15350 47280
rect 19242 47268 19248 47280
rect 19300 47268 19306 47320
rect 3234 46996 3240 47048
rect 3292 47036 3298 47048
rect 384850 47036 384856 47048
rect 3292 47008 384856 47036
rect 3292 46996 3298 47008
rect 384850 46996 384856 47008
rect 384908 46996 384914 47048
rect 3326 46860 3332 46912
rect 3384 46900 3390 46912
rect 381814 46900 381820 46912
rect 3384 46872 381820 46900
rect 3384 46860 3390 46872
rect 381814 46860 381820 46872
rect 381872 46860 381878 46912
rect 574738 46860 574744 46912
rect 574796 46900 574802 46912
rect 580166 46900 580172 46912
rect 574796 46872 580172 46900
rect 574796 46860 574802 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 4062 46792 4068 46844
rect 4120 46832 4126 46844
rect 381998 46832 382004 46844
rect 4120 46804 382004 46832
rect 4120 46792 4126 46804
rect 381998 46792 382004 46804
rect 382056 46792 382062 46844
rect 3786 46724 3792 46776
rect 3844 46764 3850 46776
rect 378870 46764 378876 46776
rect 3844 46736 378876 46764
rect 3844 46724 3850 46736
rect 378870 46724 378876 46736
rect 378928 46724 378934 46776
rect 3694 46656 3700 46708
rect 3752 46696 3758 46708
rect 378594 46696 378600 46708
rect 3752 46668 378600 46696
rect 3752 46656 3758 46668
rect 378594 46656 378600 46668
rect 378652 46656 378658 46708
rect 3602 46588 3608 46640
rect 3660 46628 3666 46640
rect 376662 46628 376668 46640
rect 3660 46600 376668 46628
rect 3660 46588 3666 46600
rect 376662 46588 376668 46600
rect 376720 46588 376726 46640
rect 3510 46520 3516 46572
rect 3568 46560 3574 46572
rect 375926 46560 375932 46572
rect 3568 46532 375932 46560
rect 3568 46520 3574 46532
rect 375926 46520 375932 46532
rect 375984 46520 375990 46572
rect 20070 46452 20076 46504
rect 20128 46492 20134 46504
rect 384574 46492 384580 46504
rect 20128 46464 384580 46492
rect 20128 46452 20134 46464
rect 384574 46452 384580 46464
rect 384632 46452 384638 46504
rect 21358 46384 21364 46436
rect 21416 46424 21422 46436
rect 384482 46424 384488 46436
rect 21416 46396 384488 46424
rect 21416 46384 21422 46396
rect 384482 46384 384488 46396
rect 384540 46384 384546 46436
rect 19978 46316 19984 46368
rect 20036 46356 20042 46368
rect 375834 46356 375840 46368
rect 20036 46328 375840 46356
rect 20036 46316 20042 46328
rect 375834 46316 375840 46328
rect 375892 46316 375898 46368
rect 14550 46248 14556 46300
rect 14608 46288 14614 46300
rect 359550 46288 359556 46300
rect 14608 46260 359556 46288
rect 14608 46248 14614 46260
rect 359550 46248 359556 46260
rect 359608 46248 359614 46300
rect 19242 46180 19248 46232
rect 19300 46220 19306 46232
rect 362586 46220 362592 46232
rect 19300 46192 362592 46220
rect 19300 46180 19306 46192
rect 362586 46180 362592 46192
rect 362644 46180 362650 46232
rect 20806 46112 20812 46164
rect 20864 46152 20870 46164
rect 361390 46152 361396 46164
rect 20864 46124 361396 46152
rect 20864 46112 20870 46124
rect 361390 46112 361396 46124
rect 361448 46112 361454 46164
rect 20714 46044 20720 46096
rect 20772 46084 20778 46096
rect 361298 46084 361304 46096
rect 20772 46056 361304 46084
rect 20772 46044 20778 46056
rect 361298 46044 361304 46056
rect 361356 46044 361362 46096
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 381354 45540 381360 45552
rect 3568 45512 381360 45540
rect 3568 45500 3574 45512
rect 381354 45500 381360 45512
rect 381412 45500 381418 45552
rect 3970 45432 3976 45484
rect 4028 45472 4034 45484
rect 381630 45472 381636 45484
rect 4028 45444 381636 45472
rect 4028 45432 4034 45444
rect 381630 45432 381636 45444
rect 381688 45432 381694 45484
rect 3878 45364 3884 45416
rect 3936 45404 3942 45416
rect 378778 45404 378784 45416
rect 3936 45376 378784 45404
rect 3936 45364 3942 45376
rect 378778 45364 378784 45376
rect 378836 45364 378842 45416
rect 21450 45296 21456 45348
rect 21508 45336 21514 45348
rect 373718 45336 373724 45348
rect 21508 45308 373724 45336
rect 21508 45296 21514 45308
rect 373718 45296 373724 45308
rect 373776 45296 373782 45348
rect 65518 45228 65524 45280
rect 65576 45268 65582 45280
rect 379422 45268 379428 45280
rect 65576 45240 379428 45268
rect 65576 45228 65582 45240
rect 379422 45228 379428 45240
rect 379480 45228 379486 45280
rect 62022 45160 62028 45212
rect 62080 45200 62086 45212
rect 378686 45200 378692 45212
rect 62080 45172 378692 45200
rect 62080 45160 62086 45172
rect 378686 45160 378692 45172
rect 378744 45160 378750 45212
rect 58434 45092 58440 45144
rect 58492 45132 58498 45144
rect 379238 45132 379244 45144
rect 58492 45104 379244 45132
rect 58492 45092 58498 45104
rect 379238 45092 379244 45104
rect 379296 45092 379302 45144
rect 54938 45024 54944 45076
rect 54996 45064 55002 45076
rect 379330 45064 379336 45076
rect 54996 45036 379336 45064
rect 54996 45024 55002 45036
rect 379330 45024 379336 45036
rect 379388 45024 379394 45076
rect 51350 44956 51356 45008
rect 51408 44996 51414 45008
rect 379146 44996 379152 45008
rect 51408 44968 379152 44996
rect 51408 44956 51414 44968
rect 379146 44956 379152 44968
rect 379204 44956 379210 45008
rect 47854 44888 47860 44940
rect 47912 44928 47918 44940
rect 381906 44928 381912 44940
rect 47912 44900 381912 44928
rect 47912 44888 47918 44900
rect 381906 44888 381912 44900
rect 381964 44888 381970 44940
rect 7650 44820 7656 44872
rect 7708 44860 7714 44872
rect 382090 44860 382096 44872
rect 7708 44832 382096 44860
rect 7708 44820 7714 44832
rect 382090 44820 382096 44832
rect 382148 44820 382154 44872
rect 69106 44752 69112 44804
rect 69164 44792 69170 44804
rect 376570 44792 376576 44804
rect 69164 44764 376576 44792
rect 69164 44752 69170 44764
rect 376570 44752 376576 44764
rect 376628 44752 376634 44804
rect 72602 44684 72608 44736
rect 72660 44724 72666 44736
rect 376386 44724 376392 44736
rect 72660 44696 376392 44724
rect 72660 44684 72666 44696
rect 376386 44684 376392 44696
rect 376444 44684 376450 44736
rect 76190 44616 76196 44668
rect 76248 44656 76254 44668
rect 376478 44656 376484 44668
rect 76248 44628 376484 44656
rect 76248 44616 76254 44628
rect 376478 44616 376484 44628
rect 376536 44616 376542 44668
rect 111610 42712 111616 42764
rect 111668 42752 111674 42764
rect 368198 42752 368204 42764
rect 111668 42724 368204 42752
rect 111668 42712 111674 42724
rect 368198 42712 368204 42724
rect 368256 42712 368262 42764
rect 108114 42644 108120 42696
rect 108172 42684 108178 42696
rect 368014 42684 368020 42696
rect 108172 42656 368020 42684
rect 108172 42644 108178 42656
rect 368014 42644 368020 42656
rect 368072 42644 368078 42696
rect 104526 42576 104532 42628
rect 104584 42616 104590 42628
rect 370774 42616 370780 42628
rect 104584 42588 370780 42616
rect 104584 42576 104590 42588
rect 370774 42576 370780 42588
rect 370832 42576 370838 42628
rect 101030 42508 101036 42560
rect 101088 42548 101094 42560
rect 370590 42548 370596 42560
rect 101088 42520 370596 42548
rect 101088 42508 101094 42520
rect 370590 42508 370596 42520
rect 370648 42508 370654 42560
rect 97442 42440 97448 42492
rect 97500 42480 97506 42492
rect 370866 42480 370872 42492
rect 97500 42452 370872 42480
rect 97500 42440 97506 42452
rect 370866 42440 370872 42452
rect 370924 42440 370930 42492
rect 93946 42372 93952 42424
rect 94004 42412 94010 42424
rect 370958 42412 370964 42424
rect 94004 42384 370964 42412
rect 94004 42372 94010 42384
rect 370958 42372 370964 42384
rect 371016 42372 371022 42424
rect 90358 42304 90364 42356
rect 90416 42344 90422 42356
rect 373534 42344 373540 42356
rect 90416 42316 373540 42344
rect 90416 42304 90422 42316
rect 373534 42304 373540 42316
rect 373592 42304 373598 42356
rect 86862 42236 86868 42288
rect 86920 42276 86926 42288
rect 373442 42276 373448 42288
rect 86920 42248 373448 42276
rect 86920 42236 86926 42248
rect 373442 42236 373448 42248
rect 373500 42236 373506 42288
rect 83274 42168 83280 42220
rect 83332 42208 83338 42220
rect 373350 42208 373356 42220
rect 83332 42180 373356 42208
rect 83332 42168 83338 42180
rect 373350 42168 373356 42180
rect 373408 42168 373414 42220
rect 79686 42100 79692 42152
rect 79744 42140 79750 42152
rect 376018 42140 376024 42152
rect 79744 42112 376024 42140
rect 79744 42100 79750 42112
rect 376018 42100 376024 42112
rect 376076 42100 376082 42152
rect 12342 42032 12348 42084
rect 12400 42072 12406 42084
rect 376202 42072 376208 42084
rect 12400 42044 376208 42072
rect 12400 42032 12406 42044
rect 376202 42032 376208 42044
rect 376260 42032 376266 42084
rect 115198 41964 115204 42016
rect 115256 42004 115262 42016
rect 367922 42004 367928 42016
rect 115256 41976 367928 42004
rect 115256 41964 115262 41976
rect 367922 41964 367928 41976
rect 367980 41964 367986 42016
rect 461578 41352 461584 41404
rect 461636 41392 461642 41404
rect 536834 41392 536840 41404
rect 461636 41364 536840 41392
rect 461636 41352 461642 41364
rect 536834 41352 536840 41364
rect 536892 41352 536898 41404
rect 118786 39992 118792 40044
rect 118844 40032 118850 40044
rect 365438 40032 365444 40044
rect 118844 40004 365444 40032
rect 118844 39992 118850 40004
rect 365438 39992 365444 40004
rect 365496 39992 365502 40044
rect 63218 39924 63224 39976
rect 63276 39964 63282 39976
rect 369394 39964 369400 39976
rect 63276 39936 369400 39964
rect 63276 39924 63282 39936
rect 369394 39924 369400 39936
rect 369452 39924 369458 39976
rect 59630 39856 59636 39908
rect 59688 39896 59694 39908
rect 366634 39896 366640 39908
rect 59688 39868 366640 39896
rect 59688 39856 59694 39868
rect 366634 39856 366640 39868
rect 366692 39856 366698 39908
rect 56042 39788 56048 39840
rect 56100 39828 56106 39840
rect 368106 39828 368112 39840
rect 56100 39800 368112 39828
rect 56100 39788 56106 39800
rect 368106 39788 368112 39800
rect 368164 39788 368170 39840
rect 52546 39720 52552 39772
rect 52604 39760 52610 39772
rect 366542 39760 366548 39772
rect 52604 39732 366548 39760
rect 52604 39720 52610 39732
rect 366542 39720 366548 39732
rect 366600 39720 366606 39772
rect 48958 39652 48964 39704
rect 49016 39692 49022 39704
rect 363874 39692 363880 39704
rect 49016 39664 363880 39692
rect 49016 39652 49022 39664
rect 363874 39652 363880 39664
rect 363932 39652 363938 39704
rect 40678 39584 40684 39636
rect 40736 39624 40742 39636
rect 363782 39624 363788 39636
rect 40736 39596 363788 39624
rect 40736 39584 40742 39596
rect 363782 39584 363788 39596
rect 363840 39584 363846 39636
rect 37182 39516 37188 39568
rect 37240 39556 37246 39568
rect 362494 39556 362500 39568
rect 37240 39528 362500 39556
rect 37240 39516 37246 39528
rect 362494 39516 362500 39528
rect 362552 39516 362558 39568
rect 33594 39448 33600 39500
rect 33652 39488 33658 39500
rect 363966 39488 363972 39500
rect 33652 39460 363972 39488
rect 33652 39448 33658 39460
rect 363966 39448 363972 39460
rect 364024 39448 364030 39500
rect 26510 39380 26516 39432
rect 26568 39420 26574 39432
rect 362402 39420 362408 39432
rect 26568 39392 362408 39420
rect 26568 39380 26574 39392
rect 362402 39380 362408 39392
rect 362460 39380 362466 39432
rect 4062 39312 4068 39364
rect 4120 39352 4126 39364
rect 365346 39352 365352 39364
rect 4120 39324 365352 39352
rect 4120 39312 4126 39324
rect 365346 39312 365352 39324
rect 365404 39312 365410 39364
rect 122282 39244 122288 39296
rect 122340 39284 122346 39296
rect 365162 39284 365168 39296
rect 122340 39256 365168 39284
rect 122340 39244 122346 39256
rect 365162 39244 365168 39256
rect 365220 39244 365226 39296
rect 102226 37204 102232 37256
rect 102284 37244 102290 37256
rect 375098 37244 375104 37256
rect 102284 37216 375104 37244
rect 102284 37204 102290 37216
rect 375098 37204 375104 37216
rect 375156 37204 375162 37256
rect 98638 37136 98644 37188
rect 98696 37176 98702 37188
rect 374914 37176 374920 37188
rect 98696 37148 374920 37176
rect 98696 37136 98702 37148
rect 374914 37136 374920 37148
rect 374972 37136 374978 37188
rect 95142 37068 95148 37120
rect 95200 37108 95206 37120
rect 376294 37108 376300 37120
rect 95200 37080 376300 37108
rect 95200 37068 95206 37080
rect 376294 37068 376300 37080
rect 376352 37068 376358 37120
rect 87966 37000 87972 37052
rect 88024 37040 88030 37052
rect 374822 37040 374828 37052
rect 88024 37012 374828 37040
rect 88024 37000 88030 37012
rect 374822 37000 374828 37012
rect 374880 37000 374886 37052
rect 91554 36932 91560 36984
rect 91612 36972 91618 36984
rect 381446 36972 381452 36984
rect 91612 36944 381452 36972
rect 91612 36932 91618 36944
rect 381446 36932 381452 36944
rect 381504 36932 381510 36984
rect 84470 36864 84476 36916
rect 84528 36904 84534 36916
rect 374730 36904 374736 36916
rect 84528 36876 374736 36904
rect 84528 36864 84534 36876
rect 374730 36864 374736 36876
rect 374788 36864 374794 36916
rect 80882 36796 80888 36848
rect 80940 36836 80946 36848
rect 373626 36836 373632 36848
rect 80940 36808 373632 36836
rect 80940 36796 80946 36808
rect 373626 36796 373632 36808
rect 373684 36796 373690 36848
rect 77386 36728 77392 36780
rect 77444 36768 77450 36780
rect 372154 36768 372160 36780
rect 77444 36740 372160 36768
rect 77444 36728 77450 36740
rect 372154 36728 372160 36740
rect 372212 36728 372218 36780
rect 73798 36660 73804 36712
rect 73856 36700 73862 36712
rect 372246 36700 372252 36712
rect 73856 36672 372252 36700
rect 73856 36660 73862 36672
rect 372246 36660 372252 36672
rect 372304 36660 372310 36712
rect 70302 36592 70308 36644
rect 70360 36632 70366 36644
rect 369302 36632 369308 36644
rect 70360 36604 369308 36632
rect 70360 36592 70366 36604
rect 369302 36592 369308 36604
rect 369360 36592 369366 36644
rect 66714 36524 66720 36576
rect 66772 36564 66778 36576
rect 370682 36564 370688 36576
rect 66772 36536 370688 36564
rect 66772 36524 66778 36536
rect 370682 36524 370688 36536
rect 370740 36524 370746 36576
rect 105722 36456 105728 36508
rect 105780 36496 105786 36508
rect 377766 36496 377772 36508
rect 105780 36468 377772 36496
rect 105780 36456 105786 36468
rect 377766 36456 377772 36468
rect 377824 36456 377830 36508
rect 119890 34416 119896 34468
rect 119948 34456 119954 34468
rect 383470 34456 383476 34468
rect 119948 34428 383476 34456
rect 119948 34416 119954 34428
rect 383470 34416 383476 34428
rect 383528 34416 383534 34468
rect 116394 34348 116400 34400
rect 116452 34388 116458 34400
rect 380526 34388 380532 34400
rect 116452 34360 380532 34388
rect 116452 34348 116458 34360
rect 380526 34348 380532 34360
rect 380584 34348 380590 34400
rect 112806 34280 112812 34332
rect 112864 34320 112870 34332
rect 377674 34320 377680 34332
rect 112864 34292 377680 34320
rect 112864 34280 112870 34292
rect 377674 34280 377680 34292
rect 377732 34280 377738 34332
rect 109310 34212 109316 34264
rect 109368 34252 109374 34264
rect 379054 34252 379060 34264
rect 109368 34224 379060 34252
rect 109368 34212 109374 34224
rect 379054 34212 379060 34224
rect 379112 34212 379118 34264
rect 50154 34144 50160 34196
rect 50212 34184 50218 34196
rect 375006 34184 375012 34196
rect 50212 34156 375012 34184
rect 50212 34144 50218 34156
rect 375006 34144 375012 34156
rect 375064 34144 375070 34196
rect 45462 34076 45468 34128
rect 45520 34116 45526 34128
rect 372338 34116 372344 34128
rect 45520 34088 372344 34116
rect 45520 34076 45526 34088
rect 372338 34076 372344 34088
rect 372396 34076 372402 34128
rect 41874 34008 41880 34060
rect 41932 34048 41938 34060
rect 369210 34048 369216 34060
rect 41932 34020 369216 34048
rect 41932 34008 41938 34020
rect 369210 34008 369216 34020
rect 369268 34008 369274 34060
rect 34790 33940 34796 33992
rect 34848 33980 34854 33992
rect 363690 33980 363696 33992
rect 34848 33952 363696 33980
rect 34848 33940 34854 33952
rect 363690 33940 363696 33952
rect 363748 33940 363754 33992
rect 31294 33872 31300 33924
rect 31352 33912 31358 33924
rect 386046 33912 386052 33924
rect 31352 33884 386052 33912
rect 31352 33872 31358 33884
rect 386046 33872 386052 33884
rect 386104 33872 386110 33924
rect 18230 33804 18236 33856
rect 18288 33844 18294 33856
rect 380434 33844 380440 33856
rect 18288 33816 380440 33844
rect 18288 33804 18294 33816
rect 380434 33804 380440 33816
rect 380492 33804 380498 33856
rect 23014 33736 23020 33788
rect 23072 33776 23078 33788
rect 385954 33776 385960 33788
rect 23072 33748 385960 33776
rect 23072 33736 23078 33748
rect 385954 33736 385960 33748
rect 386012 33736 386018 33788
rect 123478 33668 123484 33720
rect 123536 33708 123542 33720
rect 382918 33708 382924 33720
rect 123536 33680 382924 33708
rect 123536 33668 123542 33680
rect 382918 33668 382924 33680
rect 382976 33668 382982 33720
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 383194 33096 383200 33108
rect 2924 33068 383200 33096
rect 2924 33056 2930 33068
rect 383194 33056 383200 33068
rect 383252 33056 383258 33108
rect 566458 33056 566464 33108
rect 566516 33096 566522 33108
rect 580166 33096 580172 33108
rect 566516 33068 580172 33096
rect 566516 33056 566522 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 3418 31696 3424 31748
rect 3476 31736 3482 31748
rect 460290 31736 460296 31748
rect 3476 31708 460296 31736
rect 3476 31696 3482 31708
rect 460290 31696 460296 31708
rect 460348 31696 460354 31748
rect 96246 31628 96252 31680
rect 96304 31668 96310 31680
rect 378962 31668 378968 31680
rect 96304 31640 378968 31668
rect 96304 31628 96310 31640
rect 378962 31628 378968 31640
rect 379020 31628 379026 31680
rect 386138 31628 386144 31680
rect 386196 31668 386202 31680
rect 460382 31668 460388 31680
rect 386196 31640 460388 31668
rect 386196 31628 386202 31640
rect 460382 31628 460388 31640
rect 460440 31628 460446 31680
rect 92750 31560 92756 31612
rect 92808 31600 92814 31612
rect 382182 31600 382188 31612
rect 92808 31572 382188 31600
rect 92808 31560 92814 31572
rect 382182 31560 382188 31572
rect 382240 31560 382246 31612
rect 85666 31492 85672 31544
rect 85724 31532 85730 31544
rect 384758 31532 384764 31544
rect 85724 31504 384764 31532
rect 85724 31492 85730 31504
rect 384758 31492 384764 31504
rect 384816 31492 384822 31544
rect 78582 31424 78588 31476
rect 78640 31464 78646 31476
rect 383286 31464 383292 31476
rect 78640 31436 383292 31464
rect 78640 31424 78646 31436
rect 383286 31424 383292 31436
rect 383344 31424 383350 31476
rect 71498 31356 71504 31408
rect 71556 31396 71562 31408
rect 380250 31396 380256 31408
rect 71556 31368 380256 31396
rect 71556 31356 71562 31368
rect 380250 31356 380256 31368
rect 380308 31356 380314 31408
rect 67910 31288 67916 31340
rect 67968 31328 67974 31340
rect 377490 31328 377496 31340
rect 67968 31300 377496 31328
rect 67968 31288 67974 31300
rect 377490 31288 377496 31300
rect 377548 31288 377554 31340
rect 64322 31220 64328 31272
rect 64380 31260 64386 31272
rect 383378 31260 383384 31272
rect 64380 31232 383384 31260
rect 64380 31220 64386 31232
rect 383378 31220 383384 31232
rect 383436 31220 383442 31272
rect 60826 31152 60832 31204
rect 60884 31192 60890 31204
rect 380342 31192 380348 31204
rect 60884 31164 380348 31192
rect 60884 31152 60890 31164
rect 380342 31152 380348 31164
rect 380400 31152 380406 31204
rect 57238 31084 57244 31136
rect 57296 31124 57302 31136
rect 377582 31124 377588 31136
rect 57296 31096 377588 31124
rect 57296 31084 57302 31096
rect 377582 31084 377588 31096
rect 377640 31084 377646 31136
rect 14734 31016 14740 31068
rect 14792 31056 14798 31068
rect 385862 31056 385868 31068
rect 14792 31028 385868 31056
rect 14792 31016 14798 31028
rect 385862 31016 385868 31028
rect 385920 31016 385926 31068
rect 99834 30948 99840 31000
rect 99892 30988 99898 31000
rect 376110 30988 376116 31000
rect 99892 30960 376116 30988
rect 99892 30948 99898 30960
rect 376110 30948 376116 30960
rect 376168 30948 376174 31000
rect 117590 28908 117596 28960
rect 117648 28948 117654 28960
rect 369118 28948 369124 28960
rect 117648 28920 369124 28948
rect 117648 28908 117654 28920
rect 369118 28908 369124 28920
rect 369176 28908 369182 28960
rect 121086 28840 121092 28892
rect 121144 28880 121150 28892
rect 373258 28880 373264 28892
rect 121144 28852 373264 28880
rect 121144 28840 121150 28852
rect 373258 28840 373264 28852
rect 373316 28840 373322 28892
rect 114002 28772 114008 28824
rect 114060 28812 114066 28824
rect 366450 28812 366456 28824
rect 114060 28784 366456 28812
rect 114060 28772 114066 28784
rect 366450 28772 366456 28784
rect 366508 28772 366514 28824
rect 106918 28704 106924 28756
rect 106976 28744 106982 28756
rect 365254 28744 365260 28756
rect 106976 28716 365260 28744
rect 106976 28704 106982 28716
rect 365254 28704 365260 28716
rect 365312 28704 365318 28756
rect 35986 28636 35992 28688
rect 36044 28676 36050 28688
rect 383102 28676 383108 28688
rect 36044 28648 383108 28676
rect 36044 28636 36050 28648
rect 383102 28636 383108 28648
rect 383160 28636 383166 28688
rect 32398 28568 32404 28620
rect 32456 28608 32462 28620
rect 380158 28608 380164 28620
rect 32456 28580 380164 28608
rect 32456 28568 32462 28580
rect 380158 28568 380164 28580
rect 380216 28568 380222 28620
rect 28902 28500 28908 28552
rect 28960 28540 28966 28552
rect 377398 28540 377404 28552
rect 28960 28512 377404 28540
rect 28960 28500 28966 28512
rect 377398 28500 377404 28512
rect 377456 28500 377462 28552
rect 109678 28432 109684 28484
rect 109736 28472 109742 28484
rect 460934 28472 460940 28484
rect 109736 28444 460940 28472
rect 109736 28432 109742 28444
rect 460934 28432 460940 28444
rect 460992 28432 460998 28484
rect 19426 28364 19432 28416
rect 19484 28404 19490 28416
rect 372062 28404 372068 28416
rect 19484 28376 372068 28404
rect 19484 28364 19490 28376
rect 372062 28364 372068 28376
rect 372120 28364 372126 28416
rect 5258 28296 5264 28348
rect 5316 28336 5322 28348
rect 384942 28336 384948 28348
rect 5316 28308 384948 28336
rect 5316 28296 5322 28308
rect 384942 28296 384948 28308
rect 385000 28296 385006 28348
rect 43070 28228 43076 28280
rect 43128 28268 43134 28280
rect 462314 28268 462320 28280
rect 43128 28240 462320 28268
rect 43128 28228 43134 28240
rect 462314 28228 462320 28240
rect 462372 28228 462378 28280
rect 124674 28160 124680 28212
rect 124732 28200 124738 28212
rect 374638 28200 374644 28212
rect 124732 28172 374644 28200
rect 124732 28160 124738 28172
rect 374638 28160 374644 28172
rect 374696 28160 374702 28212
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 370498 20652 370504 20664
rect 3476 20624 370504 20652
rect 3476 20612 3482 20624
rect 370498 20612 370504 20624
rect 370556 20612 370562 20664
rect 570598 20612 570604 20664
rect 570656 20652 570662 20664
rect 579982 20652 579988 20664
rect 570656 20624 579988 20652
rect 570656 20612 570662 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 371878 6848 371884 6860
rect 3476 6820 371884 6848
rect 3476 6808 3482 6820
rect 371878 6808 371884 6820
rect 371936 6808 371942 6860
rect 562318 6808 562324 6860
rect 562376 6848 562382 6860
rect 580166 6848 580172 6860
rect 562376 6820 580172 6848
rect 562376 6808 562382 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 82078 4088 82084 4140
rect 82136 4128 82142 4140
rect 367738 4128 367744 4140
rect 82136 4100 367744 4128
rect 82136 4088 82142 4100
rect 367738 4088 367744 4100
rect 367796 4088 367802 4140
rect 74994 4020 75000 4072
rect 75052 4060 75058 4072
rect 367830 4060 367836 4072
rect 75052 4032 367836 4060
rect 75052 4020 75058 4032
rect 367830 4020 367836 4032
rect 367888 4020 367894 4072
rect 53742 3952 53748 4004
rect 53800 3992 53806 4004
rect 364978 3992 364984 4004
rect 53800 3964 364984 3992
rect 53800 3952 53806 3964
rect 364978 3952 364984 3964
rect 365036 3952 365042 4004
rect 46658 3884 46664 3936
rect 46716 3924 46722 3936
rect 363598 3924 363604 3936
rect 46716 3896 363604 3924
rect 46716 3884 46722 3896
rect 363598 3884 363604 3896
rect 363656 3884 363662 3936
rect 39574 3816 39580 3868
rect 39632 3856 39638 3868
rect 361206 3856 361212 3868
rect 39632 3828 361212 3856
rect 39632 3816 39638 3828
rect 361206 3816 361212 3828
rect 361264 3816 361270 3868
rect 38378 3748 38384 3800
rect 38436 3788 38442 3800
rect 366358 3788 366364 3800
rect 38436 3760 366364 3788
rect 38436 3748 38442 3760
rect 366358 3748 366364 3760
rect 366416 3748 366422 3800
rect 30098 3680 30104 3732
rect 30156 3720 30162 3732
rect 360930 3720 360936 3732
rect 30156 3692 360936 3720
rect 30156 3680 30162 3692
rect 360930 3680 360936 3692
rect 360988 3680 360994 3732
rect 44266 3612 44272 3664
rect 44324 3652 44330 3664
rect 383010 3652 383016 3664
rect 44324 3624 383016 3652
rect 44324 3612 44330 3624
rect 383010 3612 383016 3624
rect 383068 3612 383074 3664
rect 21818 3544 21824 3596
rect 21876 3584 21882 3596
rect 362310 3584 362316 3596
rect 21876 3556 362316 3584
rect 21876 3544 21882 3556
rect 362310 3544 362316 3556
rect 362368 3544 362374 3596
rect 27706 3476 27712 3528
rect 27764 3516 27770 3528
rect 384298 3516 384304 3528
rect 27764 3488 384304 3516
rect 27764 3476 27770 3488
rect 384298 3476 384304 3488
rect 384356 3476 384362 3528
rect 24210 3408 24216 3460
rect 24268 3448 24274 3460
rect 385678 3448 385684 3460
rect 24268 3420 385684 3448
rect 24268 3408 24274 3420
rect 385678 3408 385684 3420
rect 385736 3408 385742 3460
rect 89162 3340 89168 3392
rect 89220 3380 89226 3392
rect 361114 3380 361120 3392
rect 89220 3352 361120 3380
rect 89220 3340 89226 3352
rect 361114 3340 361120 3352
rect 361172 3340 361178 3392
rect 103330 3272 103336 3324
rect 103388 3312 103394 3324
rect 361022 3312 361028 3324
rect 103388 3284 361028 3312
rect 103388 3272 103394 3284
rect 361022 3272 361028 3284
rect 361080 3272 361086 3324
rect 6454 3204 6460 3256
rect 6512 3244 6518 3256
rect 109678 3244 109684 3256
rect 6512 3216 109684 3244
rect 6512 3204 6518 3216
rect 109678 3204 109684 3216
rect 109736 3204 109742 3256
rect 110506 3204 110512 3256
rect 110564 3244 110570 3256
rect 360838 3244 360844 3256
rect 110564 3216 360844 3244
rect 110564 3204 110570 3216
rect 360838 3204 360844 3216
rect 360896 3204 360902 3256
<< via1 >>
rect 397460 700816 397512 700868
rect 445024 700816 445076 700868
rect 364984 700748 365036 700800
rect 446496 700748 446548 700800
rect 332508 700680 332560 700732
rect 444104 700680 444156 700732
rect 218980 700612 219032 700664
rect 418804 700612 418856 700664
rect 235172 700544 235224 700596
rect 446404 700544 446456 700596
rect 202788 700476 202840 700528
rect 446588 700476 446640 700528
rect 154120 700408 154172 700460
rect 418896 700408 418948 700460
rect 447876 700408 447928 700460
rect 478512 700408 478564 700460
rect 170312 700340 170364 700392
rect 449164 700340 449216 700392
rect 40500 700272 40552 700324
rect 446680 700272 446732 700324
rect 447968 700272 448020 700324
rect 494796 700272 494848 700324
rect 576124 696940 576176 696992
rect 580172 696940 580224 696992
rect 300124 690616 300176 690668
rect 449256 690616 449308 690668
rect 348792 687896 348844 687948
rect 445116 687896 445168 687948
rect 8116 686468 8168 686520
rect 445208 686468 445260 686520
rect 267648 685244 267700 685296
rect 418988 685244 419040 685296
rect 89168 685176 89220 685228
rect 416044 685176 416096 685228
rect 72976 685108 73028 685160
rect 445300 685108 445352 685160
rect 3792 684632 3844 684684
rect 420276 684632 420328 684684
rect 3424 684564 3476 684616
rect 420184 684564 420236 684616
rect 3976 684496 4028 684548
rect 446864 684496 446916 684548
rect 24124 683680 24176 683732
rect 359464 683680 359516 683732
rect 21456 683612 21508 683664
rect 420828 683612 420880 683664
rect 3884 683544 3936 683596
rect 420368 683544 420420 683596
rect 3608 683476 3660 683528
rect 420644 683476 420696 683528
rect 3700 683408 3752 683460
rect 420736 683408 420788 683460
rect 3332 683340 3384 683392
rect 420552 683340 420604 683392
rect 21364 683272 21416 683324
rect 445484 683272 445536 683324
rect 3516 683204 3568 683256
rect 445392 683204 445444 683256
rect 4068 683136 4120 683188
rect 447048 683136 447100 683188
rect 11060 682728 11112 682780
rect 24124 682728 24176 682780
rect 3240 682660 3292 682712
rect 446312 682660 446364 682712
rect 6920 675792 6972 675844
rect 10968 675792 11020 675844
rect 359464 672052 359516 672104
rect 360844 672052 360896 672104
rect 447784 669944 447836 669996
rect 462320 669944 462372 669996
rect 4804 667904 4856 667956
rect 6828 667904 6880 667956
rect 361764 667904 361816 667956
rect 378784 667904 378836 667956
rect 361764 656888 361816 656940
rect 376024 656888 376076 656940
rect 3516 656140 3568 656192
rect 20904 656140 20956 656192
rect 361764 645872 361816 645924
rect 374736 645872 374788 645924
rect 571984 643084 572036 643136
rect 580172 643084 580224 643136
rect 361580 634788 361632 634840
rect 400864 634788 400916 634840
rect 3148 633360 3200 633412
rect 20904 633360 20956 633412
rect 574744 630640 574796 630692
rect 580172 630640 580224 630692
rect 361580 623772 361632 623824
rect 371884 623772 371936 623824
rect 570604 616836 570656 616888
rect 580172 616836 580224 616888
rect 361580 612824 361632 612876
rect 363604 612824 363656 612876
rect 458640 603984 458692 604036
rect 458916 603984 458968 604036
rect 459008 603712 459060 603764
rect 459468 603712 459520 603764
rect 360844 602284 360896 602336
rect 362960 602284 363012 602336
rect 459836 602080 459888 602132
rect 460112 602080 460164 602132
rect 361764 601672 361816 601724
rect 370504 601672 370556 601724
rect 460112 600244 460164 600296
rect 462320 600244 462372 600296
rect 457812 600176 457864 600228
rect 461584 600176 461636 600228
rect 458732 599768 458784 599820
rect 465080 599768 465132 599820
rect 459008 599700 459060 599752
rect 466460 599700 466512 599752
rect 457352 599632 457404 599684
rect 467104 599632 467156 599684
rect 457260 599564 457312 599616
rect 468484 599564 468536 599616
rect 457444 598748 457496 598800
rect 461676 598748 461728 598800
rect 459468 598408 459520 598460
rect 463700 598408 463752 598460
rect 362960 598340 363012 598392
rect 365444 598340 365496 598392
rect 488632 598272 488684 598324
rect 494336 598272 494388 598324
rect 460204 598204 460256 598256
rect 467932 598204 467984 598256
rect 493324 598204 493376 598256
rect 526720 598204 526772 598256
rect 457536 597524 457588 597576
rect 462964 597524 463016 597576
rect 459836 596980 459888 597032
rect 466552 596980 466604 597032
rect 457628 596912 457680 596964
rect 464344 596912 464396 596964
rect 458640 596844 458692 596896
rect 469404 596844 469456 596896
rect 450544 596776 450596 596828
rect 494980 596776 495032 596828
rect 457720 595416 457772 595468
rect 468576 595416 468628 595468
rect 459928 594056 459980 594108
rect 463792 594056 463844 594108
rect 460020 592628 460072 592680
rect 465172 592628 465224 592680
rect 361580 590792 361632 590844
rect 363696 590792 363748 590844
rect 519544 590656 519596 590708
rect 579620 590656 579672 590708
rect 365444 590588 365496 590640
rect 367744 590588 367796 590640
rect 459192 587120 459244 587172
rect 470600 587120 470652 587172
rect 459284 584400 459336 584452
rect 470692 584400 470744 584452
rect 367744 582836 367796 582888
rect 371240 582836 371292 582888
rect 361764 579640 361816 579692
rect 367744 579640 367796 579692
rect 371240 578892 371292 578944
rect 374000 578892 374052 578944
rect 511264 576852 511316 576904
rect 579620 576852 579672 576904
rect 374000 575492 374052 575544
rect 378140 575424 378192 575476
rect 378140 569848 378192 569900
rect 380348 569848 380400 569900
rect 361580 568760 361632 568812
rect 363788 568760 363840 568812
rect 515404 563048 515456 563100
rect 579896 563048 579948 563100
rect 380348 562980 380400 563032
rect 382280 562980 382332 563032
rect 382280 559716 382332 559768
rect 385040 559716 385092 559768
rect 361672 557540 361724 557592
rect 403624 557540 403676 557592
rect 385040 555568 385092 555620
rect 387064 555568 387116 555620
rect 387064 553392 387116 553444
rect 389824 553324 389876 553376
rect 457904 551284 457956 551336
rect 467196 551284 467248 551336
rect 361764 546456 361816 546508
rect 419080 546456 419132 546508
rect 389824 540948 389876 541000
rect 392308 540880 392360 540932
rect 392308 536800 392360 536852
rect 394700 536732 394752 536784
rect 361764 535440 361816 535492
rect 406384 535440 406436 535492
rect 394700 529864 394752 529916
rect 396724 529864 396776 529916
rect 361764 524424 361816 524476
rect 407764 524424 407816 524476
rect 457996 523676 458048 523728
rect 465724 523676 465776 523728
rect 482928 520888 482980 520940
rect 520280 520888 520332 520940
rect 461768 520276 461820 520328
rect 488632 520276 488684 520328
rect 459376 519528 459428 519580
rect 469312 519528 469364 519580
rect 458088 518236 458140 518288
rect 464436 518236 464488 518288
rect 449808 518168 449860 518220
rect 469864 518168 469916 518220
rect 494244 518168 494296 518220
rect 476028 517556 476080 517608
rect 494152 517556 494204 517608
rect 450360 517488 450412 517540
rect 494336 517488 494388 517540
rect 482284 517420 482336 517472
rect 450636 516808 450688 516860
rect 476028 516808 476080 516860
rect 449992 516740 450044 516792
rect 492128 516740 492180 516792
rect 3976 514768 4028 514820
rect 4804 514768 4856 514820
rect 502248 514020 502300 514072
rect 545120 514020 545172 514072
rect 361764 513340 361816 513392
rect 410524 513340 410576 513392
rect 492128 512592 492180 512644
rect 535460 512592 535512 512644
rect 396724 511912 396776 511964
rect 400956 511912 401008 511964
rect 519636 510620 519688 510672
rect 579620 510620 579672 510672
rect 494336 509872 494388 509924
rect 538220 509872 538272 509924
rect 494152 508512 494204 508564
rect 532700 508512 532752 508564
rect 495072 505724 495124 505776
rect 529940 505724 529992 505776
rect 361764 502324 361816 502376
rect 411904 502324 411956 502376
rect 461860 497700 461912 497752
rect 482652 497700 482704 497752
rect 457628 497632 457680 497684
rect 480260 497632 480312 497684
rect 457444 497564 457496 497616
rect 483848 497564 483900 497616
rect 458824 497496 458876 497548
rect 485044 497496 485096 497548
rect 453304 497428 453356 497480
rect 481640 497428 481692 497480
rect 455328 497020 455380 497072
rect 459560 497020 459612 497072
rect 456524 496952 456576 497004
rect 461032 496952 461084 497004
rect 455144 496884 455196 496936
rect 458088 496884 458140 496936
rect 452568 496816 452620 496868
rect 453672 496816 453724 496868
rect 453948 496816 454000 496868
rect 456616 496816 456668 496868
rect 400956 495456 401008 495508
rect 402244 495456 402296 495508
rect 361764 491308 361816 491360
rect 381544 491308 381596 491360
rect 518164 484372 518216 484424
rect 580172 484372 580224 484424
rect 361764 480224 361816 480276
rect 419172 480224 419224 480276
rect 515496 470568 515548 470620
rect 579988 470568 580040 470620
rect 361764 469208 361816 469260
rect 396724 469208 396776 469260
rect 494704 462408 494756 462460
rect 527640 462408 527692 462460
rect 402244 462340 402296 462392
rect 405004 462340 405056 462392
rect 450544 462340 450596 462392
rect 542360 462340 542412 462392
rect 448980 461048 449032 461100
rect 524696 461048 524748 461100
rect 468668 460980 468720 461032
rect 553860 460980 553912 461032
rect 458916 460912 458968 460964
rect 550916 460912 550968 460964
rect 361764 458192 361816 458244
rect 414664 458192 414716 458244
rect 449624 457444 449676 457496
rect 489920 457444 489972 457496
rect 569224 456764 569276 456816
rect 580172 456764 580224 456816
rect 488264 456016 488316 456068
rect 494704 456016 494756 456068
rect 452016 455472 452068 455524
rect 480996 455472 481048 455524
rect 454684 455404 454736 455456
rect 488264 455404 488316 455456
rect 449716 454724 449768 454776
rect 485780 454724 485832 454776
rect 449532 454656 449584 454708
rect 487160 454656 487212 454708
rect 459008 454044 459060 454096
rect 473728 454044 473780 454096
rect 405004 453976 405056 454028
rect 408408 453976 408460 454028
rect 408408 448536 408460 448588
rect 410432 448468 410484 448520
rect 447324 447924 447376 447976
rect 448428 447924 448480 447976
rect 459008 447924 459060 447976
rect 447232 447856 447284 447908
rect 448060 447856 448112 447908
rect 458916 447856 458968 447908
rect 447140 447788 447192 447840
rect 447692 447788 447744 447840
rect 468668 447788 468720 447840
rect 422484 447380 422536 447432
rect 447324 447380 447376 447432
rect 437388 447312 437440 447364
rect 447140 447312 447192 447364
rect 432420 447244 432472 447296
rect 447232 447244 447284 447296
rect 427452 447176 427504 447228
rect 445668 447176 445720 447228
rect 361764 447108 361816 447160
rect 399484 447108 399536 447160
rect 410432 445680 410484 445732
rect 413284 445680 413336 445732
rect 429844 445000 429896 445052
rect 447140 445000 447192 445052
rect 442632 444320 442684 444372
rect 446220 444320 446272 444372
rect 361764 436092 361816 436144
rect 416136 436092 416188 436144
rect 413284 433236 413336 433288
rect 414756 433236 414808 433288
rect 573364 430584 573416 430636
rect 579620 430584 579672 430636
rect 458088 429972 458140 430024
rect 474280 429972 474332 430024
rect 459376 429904 459428 429956
rect 476948 429904 477000 429956
rect 459468 429836 459520 429888
rect 479616 429836 479668 429888
rect 480904 429156 480956 429208
rect 482284 429156 482336 429208
rect 483664 429156 483716 429208
rect 484952 429156 485004 429208
rect 457536 428408 457588 428460
rect 471612 428408 471664 428460
rect 361764 425076 361816 425128
rect 417424 425076 417476 425128
rect 529204 423580 529256 423632
rect 530216 423580 530268 423632
rect 530584 423580 530636 423632
rect 532792 423580 532844 423632
rect 511356 423512 511408 423564
rect 523776 423512 523828 423564
rect 522304 423444 522356 423496
rect 549536 423444 549588 423496
rect 502984 423376 503036 423428
rect 522488 423376 522540 423428
rect 523684 423376 523736 423428
rect 552112 423376 552164 423428
rect 487068 423308 487120 423360
rect 526352 423308 526404 423360
rect 526444 423308 526496 423360
rect 554688 423308 554740 423360
rect 488264 423240 488316 423292
rect 528928 423240 528980 423292
rect 489644 423172 489696 423224
rect 531504 423172 531556 423224
rect 498108 423104 498160 423156
rect 545672 423104 545724 423156
rect 499304 423036 499356 423088
rect 548248 423036 548300 423088
rect 500684 422968 500736 423020
rect 550824 422968 550876 423020
rect 444288 422900 444340 422952
rect 447968 422900 448020 422952
rect 502248 422900 502300 422952
rect 553400 422900 553452 422952
rect 484308 421540 484360 421592
rect 521200 421540 521252 421592
rect 414756 420928 414808 420980
rect 420920 420860 420972 420912
rect 495348 420180 495400 420232
rect 541808 420180 541860 420232
rect 442816 419500 442868 419552
rect 447876 419500 447928 419552
rect 424692 417732 424744 417784
rect 506480 417732 506532 417784
rect 421472 417664 421524 417716
rect 503720 417664 503772 417716
rect 425980 417596 426032 417648
rect 507860 417596 507912 417648
rect 420920 417528 420972 417580
rect 425060 417528 425112 417580
rect 425336 417528 425388 417580
rect 507952 417528 508004 417580
rect 422116 417460 422168 417512
rect 503996 417460 504048 417512
rect 424048 417392 424100 417444
rect 506572 417392 506624 417444
rect 423128 416304 423180 416356
rect 423588 416304 423640 416356
rect 486976 416032 487028 416084
rect 527640 416032 527692 416084
rect 361580 413992 361632 414044
rect 443644 413992 443696 414044
rect 425060 413924 425112 413976
rect 427084 413924 427136 413976
rect 361580 402976 361632 403028
rect 439504 402976 439556 403028
rect 503444 402228 503496 402280
rect 557540 402228 557592 402280
rect 497924 400868 497976 400920
rect 546500 400868 546552 400920
rect 494612 399440 494664 399492
rect 539600 399440 539652 399492
rect 493968 398080 494020 398132
rect 538220 398080 538272 398132
rect 427084 397400 427136 397452
rect 428464 397400 428516 397452
rect 493140 396720 493192 396772
rect 536840 396720 536892 396772
rect 460756 395292 460808 395344
rect 483664 395292 483716 395344
rect 492404 395292 492456 395344
rect 535460 395292 535512 395344
rect 496728 394000 496780 394052
rect 543740 394000 543792 394052
rect 423496 393932 423548 393984
rect 505560 393932 505612 393984
rect 463608 392572 463660 392624
rect 487160 392572 487212 392624
rect 491576 392572 491628 392624
rect 534172 392572 534224 392624
rect 361580 391960 361632 392012
rect 443736 391960 443788 392012
rect 495716 391280 495768 391332
rect 542360 391280 542412 391332
rect 423588 391212 423640 391264
rect 505284 391212 505336 391264
rect 459652 389852 459704 389904
rect 480904 389852 480956 389904
rect 464896 389784 464948 389836
rect 489920 389784 489972 389836
rect 490564 389784 490616 389836
rect 534080 389784 534132 389836
rect 465080 389240 465132 389292
rect 465908 389240 465960 389292
rect 466460 389240 466512 389292
rect 467380 389240 467432 389292
rect 470600 389240 470652 389292
rect 471060 389240 471112 389292
rect 486424 389240 486476 389292
rect 487068 389240 487120 389292
rect 497464 389240 497516 389292
rect 498108 389240 498160 389292
rect 506480 389240 506532 389292
rect 507124 389240 507176 389292
rect 507860 389240 507912 389292
rect 508596 389240 508648 389292
rect 453028 389104 453080 389156
rect 454040 389104 454092 389156
rect 456708 389104 456760 389156
rect 457536 389104 457588 389156
rect 468484 389036 468536 389088
rect 474372 389036 474424 389088
rect 467104 388968 467156 389020
rect 475108 388968 475160 389020
rect 461124 388900 461176 388952
rect 463608 388900 463660 388952
rect 468576 388900 468628 388952
rect 478788 388900 478840 388952
rect 502340 388900 502392 388952
rect 467196 388832 467248 388884
rect 480260 388832 480312 388884
rect 483940 388832 483992 388884
rect 502984 388832 503036 388884
rect 526444 388832 526496 388884
rect 461676 388764 461728 388816
rect 475844 388764 475896 388816
rect 499396 388764 499448 388816
rect 522304 388764 522356 388816
rect 464344 388696 464396 388748
rect 478052 388696 478104 388748
rect 500868 388696 500920 388748
rect 523684 388696 523736 388748
rect 462964 388628 463016 388680
rect 476580 388628 476632 388680
rect 484676 388628 484728 388680
rect 511356 388628 511408 388680
rect 465724 388560 465776 388612
rect 480996 388560 481048 388612
rect 485412 388560 485464 388612
rect 524420 388560 524472 388612
rect 447876 388492 447928 388544
rect 458824 388492 458876 388544
rect 464528 388492 464580 388544
rect 481732 388492 481784 388544
rect 489828 388492 489880 388544
rect 530584 388492 530636 388544
rect 448336 388424 448388 388476
rect 461768 388424 461820 388476
rect 463056 388424 463108 388476
rect 482468 388424 482520 388476
rect 488356 388424 488408 388476
rect 529204 388424 529256 388476
rect 461584 388016 461636 388068
rect 462596 388016 462648 388068
rect 462136 387812 462188 387864
rect 464896 387812 464948 387864
rect 428464 387744 428516 387796
rect 431224 387744 431276 387796
rect 442724 387744 442776 387796
rect 447140 387744 447192 387796
rect 450728 387336 450780 387388
rect 454684 387336 454736 387388
rect 447416 387268 447468 387320
rect 457444 387268 457496 387320
rect 447600 387200 447652 387252
rect 461860 387200 461912 387252
rect 449808 387132 449860 387184
rect 491300 387132 491352 387184
rect 441528 387064 441580 387116
rect 447784 387064 447836 387116
rect 449440 387064 449492 387116
rect 513380 387064 513432 387116
rect 448428 386588 448480 386640
rect 553952 386588 554004 386640
rect 382924 386520 382976 386572
rect 512092 386520 512144 386572
rect 374644 386452 374696 386504
rect 512276 386452 512328 386504
rect 369124 386384 369176 386436
rect 512000 386384 512052 386436
rect 448152 385976 448204 386028
rect 453304 385976 453356 386028
rect 447968 385636 448020 385688
rect 457352 385636 457404 385688
rect 448244 385364 448296 385416
rect 452016 385364 452068 385416
rect 449348 385092 449400 385144
rect 563428 385092 563480 385144
rect 373264 385024 373316 385076
rect 512184 385024 512236 385076
rect 513288 383732 513340 383784
rect 530584 383732 530636 383784
rect 512460 383664 512512 383716
rect 548524 383664 548576 383716
rect 362224 383596 362276 383648
rect 447140 383596 447192 383648
rect 378784 383528 378836 383580
rect 447232 383528 447284 383580
rect 512644 382984 512696 383036
rect 519728 382984 519780 383036
rect 513288 382576 513340 382628
rect 518256 382576 518308 382628
rect 512460 382440 512512 382492
rect 515588 382440 515640 382492
rect 374736 382168 374788 382220
rect 447232 382168 447284 382220
rect 376024 382100 376076 382152
rect 447140 382100 447192 382152
rect 361580 380876 361632 380928
rect 443828 380876 443880 380928
rect 512460 380876 512512 380928
rect 547144 380876 547196 380928
rect 363604 380808 363656 380860
rect 447508 380808 447560 380860
rect 371884 380740 371936 380792
rect 447140 380740 447192 380792
rect 400864 380672 400916 380724
rect 447232 380672 447284 380724
rect 512552 379720 512604 379772
rect 515680 379720 515732 379772
rect 513288 379516 513340 379568
rect 549904 379516 549956 379568
rect 363696 379448 363748 379500
rect 447324 379448 447376 379500
rect 370504 379380 370556 379432
rect 447140 379380 447192 379432
rect 513288 378292 513340 378344
rect 522304 378292 522356 378344
rect 512828 378224 512880 378276
rect 547236 378224 547288 378276
rect 514024 378156 514076 378208
rect 580172 378156 580224 378208
rect 363788 378088 363840 378140
rect 447232 378088 447284 378140
rect 367744 378020 367796 378072
rect 447140 378020 447192 378072
rect 513196 377408 513248 377460
rect 548616 377408 548668 377460
rect 512828 376728 512880 376780
rect 516232 376728 516284 376780
rect 403624 376660 403676 376712
rect 447140 376660 447192 376712
rect 419080 376592 419132 376644
rect 447232 376592 447284 376644
rect 513104 375980 513156 376032
rect 544384 375980 544436 376032
rect 513288 375912 513340 375964
rect 518900 375912 518952 375964
rect 513288 375368 513340 375420
rect 518348 375368 518400 375420
rect 406384 375300 406436 375352
rect 447140 375300 447192 375352
rect 407764 375232 407816 375284
rect 447232 375232 447284 375284
rect 512092 374008 512144 374060
rect 520280 374008 520332 374060
rect 410524 373940 410576 373992
rect 447140 373940 447192 373992
rect 411904 373872 411956 373924
rect 447232 373872 447284 373924
rect 512460 372716 512512 372768
rect 521660 372716 521712 372768
rect 512092 372648 512144 372700
rect 514760 372648 514812 372700
rect 512000 372580 512052 372632
rect 514852 372580 514904 372632
rect 381544 372512 381596 372564
rect 447140 372512 447192 372564
rect 419172 372444 419224 372496
rect 447232 372444 447284 372496
rect 512460 371900 512512 371952
rect 516324 371900 516376 371952
rect 396724 371152 396776 371204
rect 447140 371152 447192 371204
rect 414664 371084 414716 371136
rect 447232 371084 447284 371136
rect 512460 370336 512512 370388
rect 517612 370336 517664 370388
rect 512828 369928 512880 369980
rect 516876 369928 516928 369980
rect 361580 369860 361632 369912
rect 409880 369860 409932 369912
rect 513288 369860 513340 369912
rect 523040 369860 523092 369912
rect 399484 369792 399536 369844
rect 447140 369792 447192 369844
rect 416136 369724 416188 369776
rect 447232 369724 447284 369776
rect 431224 369656 431276 369708
rect 432880 369656 432932 369708
rect 512828 368568 512880 368620
rect 516416 368568 516468 368620
rect 513288 368500 513340 368552
rect 520372 368500 520424 368552
rect 417424 368432 417476 368484
rect 447140 368432 447192 368484
rect 443644 368364 443696 368416
rect 447232 368364 447284 368416
rect 513288 367208 513340 367260
rect 517980 367208 518032 367260
rect 512000 367072 512052 367124
rect 514116 367072 514168 367124
rect 439504 367004 439556 367056
rect 447140 367004 447192 367056
rect 443736 366936 443788 366988
rect 447232 366936 447284 366988
rect 512000 365848 512052 365900
rect 514208 365848 514260 365900
rect 513288 365712 513340 365764
rect 521752 365712 521804 365764
rect 409880 365644 409932 365696
rect 447140 365644 447192 365696
rect 443828 365576 443880 365628
rect 447232 365576 447284 365628
rect 512644 365168 512696 365220
rect 520464 365168 520516 365220
rect 513288 364352 513340 364404
rect 523132 364352 523184 364404
rect 576216 364352 576268 364404
rect 580172 364352 580224 364404
rect 432696 362992 432748 363044
rect 447140 362992 447192 363044
rect 512460 362992 512512 363044
rect 521844 362992 521896 363044
rect 432788 362924 432840 362976
rect 447232 362924 447284 362976
rect 512000 362312 512052 362364
rect 513656 362312 513708 362364
rect 442264 361632 442316 361684
rect 447232 361632 447284 361684
rect 432604 361564 432656 361616
rect 447140 361564 447192 361616
rect 513012 361564 513064 361616
rect 520556 361564 520608 361616
rect 512920 360952 512972 361004
rect 518992 360952 519044 361004
rect 512368 360680 512420 360732
rect 515036 360680 515088 360732
rect 513196 360544 513248 360596
rect 517704 360544 517756 360596
rect 439780 360272 439832 360324
rect 447232 360272 447284 360324
rect 436928 360204 436980 360256
rect 447140 360204 447192 360256
rect 547236 360136 547288 360188
rect 552020 360136 552072 360188
rect 530584 360068 530636 360120
rect 566740 360068 566792 360120
rect 522304 360000 522356 360052
rect 550640 360000 550692 360052
rect 549904 359932 549956 359984
rect 554964 359932 555016 359984
rect 547144 359864 547196 359916
rect 558184 359864 558236 359916
rect 515680 359796 515732 359848
rect 553768 359796 553820 359848
rect 548524 359728 548576 359780
rect 565268 359932 565320 359984
rect 443828 358844 443880 358896
rect 447232 358844 447284 358896
rect 435456 358776 435508 358828
rect 447140 358776 447192 358828
rect 512736 358776 512788 358828
rect 517888 358776 517940 358828
rect 548616 358708 548668 358760
rect 556712 358708 556764 358760
rect 518256 358640 518308 358692
rect 562600 358640 562652 358692
rect 519728 358572 519780 358624
rect 564072 358572 564124 358624
rect 544384 358504 544436 358556
rect 559656 358504 559708 358556
rect 515588 358436 515640 358488
rect 561128 358436 561180 358488
rect 513288 357824 513340 357876
rect 519084 357824 519136 357876
rect 513288 356056 513340 356108
rect 523224 356056 523276 356108
rect 513288 354968 513340 355020
rect 519176 354968 519228 355020
rect 512000 353948 512052 354000
rect 513748 353948 513800 354000
rect 513288 353472 513340 353524
rect 517796 353472 517848 353524
rect 445668 353268 445720 353320
rect 447876 353268 447928 353320
rect 446220 353064 446272 353116
rect 447784 353064 447836 353116
rect 512000 352384 512052 352436
rect 515128 352384 515180 352436
rect 513288 351908 513340 351960
rect 521936 351908 521988 351960
rect 512644 350888 512696 350940
rect 519360 350888 519412 350940
rect 512552 350616 512604 350668
rect 515220 350616 515272 350668
rect 407028 350548 407080 350600
rect 447140 350548 447192 350600
rect 513288 349528 513340 349580
rect 519452 349528 519504 349580
rect 512000 349392 512052 349444
rect 514944 349392 514996 349444
rect 512000 349256 512052 349308
rect 513840 349256 513892 349308
rect 432880 349052 432932 349104
rect 437020 349052 437072 349104
rect 512920 348032 512972 348084
rect 516508 348032 516560 348084
rect 361764 347760 361816 347812
rect 402244 347760 402296 347812
rect 513288 347760 513340 347812
rect 523316 347760 523368 347812
rect 362224 347692 362276 347744
rect 447140 347692 447192 347744
rect 513288 346944 513340 346996
rect 519268 346944 519320 346996
rect 512552 346536 512604 346588
rect 515312 346536 515364 346588
rect 513288 346468 513340 346520
rect 518072 346468 518124 346520
rect 513012 343816 513064 343868
rect 516692 343816 516744 343868
rect 512828 343748 512880 343800
rect 517520 343748 517572 343800
rect 513012 342320 513064 342372
rect 516784 342320 516836 342372
rect 513288 341368 513340 341420
rect 520648 341368 520700 341420
rect 513288 341096 513340 341148
rect 518256 341096 518308 341148
rect 444196 340960 444248 341012
rect 447232 340960 447284 341012
rect 361764 340892 361816 340944
rect 447140 340892 447192 340944
rect 512644 339736 512696 339788
rect 516140 339736 516192 339788
rect 431224 339532 431276 339584
rect 447140 339532 447192 339584
rect 371884 339464 371936 339516
rect 447232 339464 447284 339516
rect 512644 339464 512696 339516
rect 515588 339464 515640 339516
rect 513012 338376 513064 338428
rect 516600 338376 516652 338428
rect 436836 338172 436888 338224
rect 447140 338172 447192 338224
rect 435364 338104 435416 338156
rect 447232 338104 447284 338156
rect 450084 337968 450136 338020
rect 450360 337968 450412 338020
rect 402244 337356 402296 337408
rect 447876 337356 447928 337408
rect 448428 337356 448480 337408
rect 513196 337288 513248 337340
rect 519728 337288 519780 337340
rect 513288 337152 513340 337204
rect 520924 337152 520976 337204
rect 440884 336948 440936 337000
rect 447140 336948 447192 337000
rect 416780 336880 416832 336932
rect 450360 336880 450412 336932
rect 413100 336812 413152 336864
rect 450176 336812 450228 336864
rect 409420 336744 409472 336796
rect 450728 336744 450780 336796
rect 418896 336336 418948 336388
rect 440976 336336 441028 336388
rect 418988 336268 419040 336320
rect 441252 336268 441304 336320
rect 418804 336200 418856 336252
rect 441160 336200 441212 336252
rect 416044 336132 416096 336184
rect 441068 336132 441120 336184
rect 413652 336064 413704 336116
rect 449440 336064 449492 336116
rect 362224 335996 362276 336048
rect 444196 335996 444248 336048
rect 443736 335656 443788 335708
rect 447232 335656 447284 335708
rect 399484 335316 399536 335368
rect 447140 335316 447192 335368
rect 439688 335044 439740 335096
rect 447508 335044 447560 335096
rect 420552 334976 420604 335028
rect 439872 334976 439924 335028
rect 420828 334908 420880 334960
rect 442356 334908 442408 334960
rect 420276 334840 420328 334892
rect 442448 334840 442500 334892
rect 513288 334840 513340 334892
rect 520740 334840 520792 334892
rect 420184 334772 420236 334824
rect 444932 334772 444984 334824
rect 420276 334704 420328 334756
rect 445668 334704 445720 334756
rect 513012 334704 513064 334756
rect 520832 334704 520884 334756
rect 420644 334636 420696 334688
rect 449532 334636 449584 334688
rect 420736 334568 420788 334620
rect 449624 334568 449676 334620
rect 443644 334024 443696 334076
rect 447232 334024 447284 334076
rect 364064 333956 364116 334008
rect 447140 333956 447192 334008
rect 439596 332664 439648 332716
rect 447232 332664 447284 332716
rect 436744 332596 436796 332648
rect 447140 332596 447192 332648
rect 512644 331304 512696 331356
rect 513932 331304 513984 331356
rect 447140 330488 447192 330540
rect 447876 330488 447928 330540
rect 450084 330488 450136 330540
rect 450728 330488 450780 330540
rect 439504 330420 439556 330472
rect 447416 330420 447468 330472
rect 448060 330420 448112 330472
rect 442908 330352 442960 330404
rect 447232 330352 447284 330404
rect 432788 330216 432840 330268
rect 439780 330216 439832 330268
rect 512644 328584 512696 328636
rect 516968 328584 517020 328636
rect 436008 328516 436060 328568
rect 449900 328516 449952 328568
rect 431868 328448 431920 328500
rect 450452 328448 450504 328500
rect 446312 327428 446364 327480
rect 449716 327428 449768 327480
rect 509332 326408 509384 326460
rect 509976 326408 510028 326460
rect 509424 326340 509476 326392
rect 509700 326340 509752 326392
rect 437020 324980 437072 325032
rect 439320 324980 439372 325032
rect 432880 324912 432932 324964
rect 442264 324912 442316 324964
rect 510436 324912 510488 324964
rect 580632 324912 580684 324964
rect 511908 323620 511960 323672
rect 580172 323620 580224 323672
rect 510528 323552 510580 323604
rect 580540 323552 580592 323604
rect 432604 322940 432656 322992
rect 436928 322940 436980 322992
rect 445576 322736 445628 322788
rect 459652 322668 459704 322720
rect 570604 322872 570656 322924
rect 569224 322804 569276 322856
rect 461308 322668 461360 322720
rect 473314 322736 473366 322788
rect 571984 322736 572036 322788
rect 459100 322532 459152 322584
rect 473452 322668 473504 322720
rect 480628 322668 480680 322720
rect 462964 322600 463016 322652
rect 478144 322600 478196 322652
rect 480904 322600 480956 322652
rect 519636 322668 519688 322720
rect 469036 322532 469088 322584
rect 445024 322464 445076 322516
rect 480628 322532 480680 322584
rect 515404 322600 515456 322652
rect 515496 322532 515548 322584
rect 446588 322396 446640 322448
rect 507400 322464 507452 322516
rect 509884 322464 509936 322516
rect 439872 322328 439924 322380
rect 473452 322396 473504 322448
rect 442356 322260 442408 322312
rect 463792 322260 463844 322312
rect 482284 322328 482336 322380
rect 473452 322260 473504 322312
rect 478144 322260 478196 322312
rect 480628 322260 480680 322312
rect 506940 322260 506992 322312
rect 511448 322260 511500 322312
rect 439320 322192 439372 322244
rect 474280 322192 474332 322244
rect 475108 322192 475160 322244
rect 475384 322192 475436 322244
rect 490288 322192 490340 322244
rect 490564 322192 490616 322244
rect 442448 322124 442500 322176
rect 459376 322056 459428 322108
rect 462964 322056 463016 322108
rect 484216 322124 484268 322176
rect 509424 321988 509476 322040
rect 509976 321988 510028 322040
rect 507492 321784 507544 321836
rect 511172 321784 511224 321836
rect 458088 321512 458140 321564
rect 580816 321512 580868 321564
rect 458364 321444 458416 321496
rect 580724 321444 580776 321496
rect 446496 321376 446548 321428
rect 460848 321376 460900 321428
rect 468576 321376 468628 321428
rect 576216 321376 576268 321428
rect 449164 321308 449216 321360
rect 461676 321308 461728 321360
rect 469956 321308 470008 321360
rect 574744 321308 574796 321360
rect 479340 321240 479392 321292
rect 573364 321240 573416 321292
rect 444932 321172 444984 321224
rect 484584 321172 484636 321224
rect 507676 321172 507728 321224
rect 509976 321172 510028 321224
rect 447508 321104 447560 321156
rect 463332 321104 463384 321156
rect 479064 321104 479116 321156
rect 514024 321104 514076 321156
rect 447048 321036 447100 321088
rect 484032 321036 484084 321088
rect 507308 321036 507360 321088
rect 517520 321036 517572 321088
rect 460664 320968 460716 321020
rect 516140 320968 516192 321020
rect 441160 320900 441212 320952
rect 471888 320900 471940 320952
rect 502248 320900 502300 320952
rect 580264 320900 580316 320952
rect 446404 320832 446456 320884
rect 451832 320832 451884 320884
rect 444104 320764 444156 320816
rect 459928 320832 459980 320884
rect 580356 320832 580408 320884
rect 481824 320764 481876 320816
rect 507584 320764 507636 320816
rect 451924 320696 451976 320748
rect 461400 320696 461452 320748
rect 507124 320696 507176 320748
rect 512644 320764 512696 320816
rect 512828 320764 512880 320816
rect 441068 320628 441120 320680
rect 446864 320560 446916 320612
rect 447508 320560 447560 320612
rect 472440 320628 472492 320680
rect 513380 320696 513432 320748
rect 513472 320628 513524 320680
rect 449716 320560 449768 320612
rect 463056 320560 463108 320612
rect 441252 320492 441304 320544
rect 482100 320492 482152 320544
rect 441528 320424 441580 320476
rect 481272 320424 481324 320476
rect 507768 320220 507820 320272
rect 511080 320220 511132 320272
rect 479892 320084 479944 320136
rect 580448 320084 580500 320136
rect 442724 320016 442776 320068
rect 460572 320016 460624 320068
rect 480720 320016 480772 320068
rect 576124 320016 576176 320068
rect 444288 319948 444340 320000
rect 460296 319948 460348 320000
rect 469680 319948 469732 320000
rect 511264 319948 511316 320000
rect 449624 319880 449676 319932
rect 463608 319880 463660 319932
rect 468852 319880 468904 319932
rect 510436 319880 510488 319932
rect 449256 319812 449308 319864
rect 461124 319812 461176 319864
rect 469404 319812 469456 319864
rect 510528 319812 510580 319864
rect 449440 319744 449492 319796
rect 471060 319744 471112 319796
rect 480168 319744 480220 319796
rect 519544 319744 519596 319796
rect 445116 319676 445168 319728
rect 471336 319676 471388 319728
rect 479616 319676 479668 319728
rect 518164 319676 518216 319728
rect 449532 319608 449584 319660
rect 474096 319608 474148 319660
rect 478788 319608 478840 319660
rect 511908 319608 511960 319660
rect 445484 319540 445536 319592
rect 462780 319540 462832 319592
rect 470232 319540 470284 319592
rect 502248 319540 502300 319592
rect 502800 319540 502852 319592
rect 533344 319540 533396 319592
rect 445392 319472 445444 319524
rect 483480 319472 483532 319524
rect 498660 319472 498712 319524
rect 534724 319472 534776 319524
rect 460296 319404 460348 319456
rect 476304 319404 476356 319456
rect 502156 319404 502208 319456
rect 538864 319404 538916 319456
rect 440976 319336 441028 319388
rect 472164 319336 472216 319388
rect 445668 319268 445720 319320
rect 473820 319268 473872 319320
rect 445300 319200 445352 319252
rect 482928 319200 482980 319252
rect 487252 319200 487304 319252
rect 488356 319200 488408 319252
rect 442816 319132 442868 319184
rect 470784 319132 470836 319184
rect 483664 319132 483716 319184
rect 484860 319132 484912 319184
rect 494152 319132 494204 319184
rect 494428 319132 494480 319184
rect 509424 319132 509476 319184
rect 509700 319132 509752 319184
rect 446956 319064 447008 319116
rect 483756 319064 483808 319116
rect 484768 319064 484820 319116
rect 485596 319064 485648 319116
rect 485872 319064 485924 319116
rect 486976 319064 487028 319116
rect 487804 319064 487856 319116
rect 488356 319064 488408 319116
rect 488908 319064 488960 319116
rect 489460 319064 489512 319116
rect 491668 319064 491720 319116
rect 492220 319064 492272 319116
rect 493324 319064 493376 319116
rect 493876 319064 493928 319116
rect 494704 319064 494756 319116
rect 495256 319064 495308 319116
rect 499948 319064 500000 319116
rect 500224 319064 500276 319116
rect 501328 319064 501380 319116
rect 501880 319064 501932 319116
rect 464068 318996 464120 319048
rect 464620 318996 464672 319048
rect 465172 318996 465224 319048
rect 465724 318996 465776 319048
rect 466828 318996 466880 319048
rect 467380 318996 467432 319048
rect 475108 318996 475160 319048
rect 475660 318996 475712 319048
rect 484492 318996 484544 319048
rect 485320 318996 485372 319048
rect 488632 318996 488684 319048
rect 489184 318996 489236 319048
rect 491392 318996 491444 319048
rect 492496 318996 492548 319048
rect 493048 318996 493100 319048
rect 493600 318996 493652 319048
rect 463792 318928 463844 318980
rect 464896 318928 464948 318980
rect 467104 318928 467156 318980
rect 467656 318928 467708 318980
rect 490288 318860 490340 318912
rect 491116 318860 491168 318912
rect 432052 318248 432104 318300
rect 435456 318248 435508 318300
rect 454684 318180 454736 318232
rect 488724 318180 488776 318232
rect 451924 318112 451976 318164
rect 495624 318112 495676 318164
rect 496176 318112 496228 318164
rect 540980 318112 541032 318164
rect 477684 318044 477736 318096
rect 547144 318044 547196 318096
rect 478512 317364 478564 317416
rect 479524 317364 479576 317416
rect 457812 317024 457864 317076
rect 461584 317024 461636 317076
rect 501420 316888 501472 316940
rect 539692 316888 539744 316940
rect 500316 316820 500368 316872
rect 539600 316820 539652 316872
rect 487344 316752 487396 316804
rect 529940 316752 529992 316804
rect 458916 316684 458968 316736
rect 491484 316684 491536 316736
rect 497004 316684 497056 316736
rect 543004 316684 543056 316736
rect 457444 316072 457496 316124
rect 457996 316072 458048 316124
rect 465448 316072 465500 316124
rect 466000 316072 466052 316124
rect 486332 316004 486384 316056
rect 486516 316004 486568 316056
rect 361764 315936 361816 315988
rect 371884 315936 371936 315988
rect 501880 315392 501932 315444
rect 539784 315392 539836 315444
rect 457444 315324 457496 315376
rect 491760 315324 491812 315376
rect 502984 315324 503036 315376
rect 542728 315324 542780 315376
rect 455880 315256 455932 315308
rect 562324 315256 562376 315308
rect 454776 313964 454828 314016
rect 491944 313964 491996 314016
rect 497464 313964 497516 314016
rect 542452 313964 542504 314016
rect 432696 313896 432748 313948
rect 443828 313896 443880 313948
rect 477040 313896 477092 313948
rect 566464 313896 566516 313948
rect 482652 313284 482704 313336
rect 485044 313284 485096 313336
rect 469036 313216 469088 313268
rect 580172 313216 580224 313268
rect 467380 312536 467432 312588
rect 551284 312536 551336 312588
rect 459008 311176 459060 311228
rect 493048 311176 493100 311228
rect 503536 311176 503588 311228
rect 538956 311176 539008 311228
rect 462964 311108 463016 311160
rect 464344 311108 464396 311160
rect 478144 311108 478196 311160
rect 548524 311108 548576 311160
rect 482468 310496 482520 310548
rect 483664 310496 483716 310548
rect 461676 310292 461728 310344
rect 464160 310292 464212 310344
rect 454960 309816 455012 309868
rect 494428 309816 494480 309868
rect 497648 309816 497700 309868
rect 542544 309816 542596 309868
rect 447968 309748 448020 309800
rect 533436 309748 533488 309800
rect 452016 308456 452068 308508
rect 494796 308456 494848 308508
rect 498844 308456 498896 308508
rect 542636 308456 542688 308508
rect 457168 308388 457220 308440
rect 536104 308388 536156 308440
rect 474004 307776 474056 307828
rect 482652 307776 482704 307828
rect 3424 307708 3476 307760
rect 4804 307708 4856 307760
rect 481088 307300 481140 307352
rect 482468 307300 482520 307352
rect 454868 307164 454920 307216
rect 490288 307164 490340 307216
rect 477316 307096 477368 307148
rect 544384 307096 544436 307148
rect 380164 307028 380216 307080
rect 506940 307028 506992 307080
rect 383200 306280 383252 306332
rect 465448 306280 465500 306332
rect 382004 306212 382056 306264
rect 465356 306212 465408 306264
rect 378876 306144 378928 306196
rect 463792 306144 463844 306196
rect 384672 306076 384724 306128
rect 475660 306076 475712 306128
rect 381820 306008 381872 306060
rect 475108 306008 475160 306060
rect 378784 305940 378836 305992
rect 475476 305940 475528 305992
rect 477408 305940 477460 305992
rect 569224 305940 569276 305992
rect 384856 305872 384908 305924
rect 486148 305872 486200 305924
rect 384488 305804 384540 305856
rect 486516 305804 486568 305856
rect 381636 305736 381688 305788
rect 486056 305736 486108 305788
rect 500132 305736 500184 305788
rect 541072 305736 541124 305788
rect 365168 305668 365220 305720
rect 516232 305668 516284 305720
rect 360844 305600 360896 305652
rect 512092 305600 512144 305652
rect 384396 305532 384448 305584
rect 465540 305532 465592 305584
rect 384580 305464 384632 305516
rect 465172 305464 465224 305516
rect 458824 305396 458876 305448
rect 489000 305396 489052 305448
rect 361764 304920 361816 304972
rect 431224 304920 431276 304972
rect 488264 304512 488316 304564
rect 531412 304512 531464 304564
rect 385776 304444 385828 304496
rect 507032 304444 507084 304496
rect 383108 304376 383160 304428
rect 520924 304376 520976 304428
rect 361028 304308 361080 304360
rect 512184 304308 512236 304360
rect 360936 304240 360988 304292
rect 512736 304240 512788 304292
rect 459376 304104 459428 304156
rect 461676 304104 461728 304156
rect 378600 303560 378652 303612
rect 484768 303560 484820 303612
rect 375840 303492 375892 303544
rect 484492 303492 484544 303544
rect 371884 303424 371936 303476
rect 485872 303424 485924 303476
rect 456340 303356 456392 303408
rect 574744 303356 574796 303408
rect 376024 303288 376076 303340
rect 509516 303288 509568 303340
rect 376484 303220 376536 303272
rect 510804 303220 510856 303272
rect 379428 303152 379480 303204
rect 515220 303152 515272 303204
rect 379244 303084 379296 303136
rect 515312 303084 515364 303136
rect 376392 303016 376444 303068
rect 513748 303016 513800 303068
rect 376576 302948 376628 303000
rect 515128 302948 515180 303000
rect 367744 302880 367796 302932
rect 512368 302880 512420 302932
rect 373724 302812 373776 302864
rect 475384 302812 475436 302864
rect 376668 302744 376720 302796
rect 474832 302744 474884 302796
rect 375932 302676 375984 302728
rect 464068 302676 464120 302728
rect 478880 301656 478932 301708
rect 481088 301656 481140 301708
rect 456616 301588 456668 301640
rect 571984 301588 572036 301640
rect 367836 301520 367888 301572
rect 512460 301520 512512 301572
rect 364984 301452 365036 301504
rect 512552 301452 512604 301504
rect 373356 300772 373408 300824
rect 510620 300772 510672 300824
rect 370872 300704 370924 300756
rect 509332 300704 509384 300756
rect 373540 300636 373592 300688
rect 513656 300636 513708 300688
rect 373448 300568 373500 300620
rect 515036 300568 515088 300620
rect 370964 300500 371016 300552
rect 513564 300500 513616 300552
rect 370780 300432 370832 300484
rect 516416 300432 516468 300484
rect 367928 300364 367980 300416
rect 514852 300364 514904 300416
rect 368204 300296 368256 300348
rect 516324 300296 516376 300348
rect 363604 300228 363656 300280
rect 512644 300228 512696 300280
rect 368020 300160 368072 300212
rect 517612 300160 517664 300212
rect 361120 300092 361172 300144
rect 512276 300092 512328 300144
rect 376208 300024 376260 300076
rect 510160 300024 510212 300076
rect 467748 299956 467800 300008
rect 580264 299956 580316 300008
rect 457536 299888 457588 299940
rect 495808 299888 495860 299940
rect 461584 299412 461636 299464
rect 580172 299412 580224 299464
rect 478144 298936 478196 298988
rect 478880 298936 478932 298988
rect 456708 297984 456760 298036
rect 573364 297984 573416 298036
rect 383016 297916 383068 297968
rect 518256 297916 518308 297968
rect 363972 297848 364024 297900
rect 507676 297848 507728 297900
rect 362500 297780 362552 297832
rect 507768 297780 507820 297832
rect 368112 297712 368164 297764
rect 518072 297712 518124 297764
rect 366548 297644 366600 297696
rect 516692 297644 516744 297696
rect 362316 297576 362368 297628
rect 513932 297576 513984 297628
rect 363788 297508 363840 297560
rect 515588 297508 515640 297560
rect 365444 297440 365496 297492
rect 518348 297440 518400 297492
rect 363880 297372 363932 297424
rect 516784 297372 516836 297424
rect 460388 296692 460440 296744
rect 462964 296692 463016 296744
rect 457996 295944 458048 295996
rect 576124 295944 576176 295996
rect 476856 295332 476908 295384
rect 478144 295332 478196 295384
rect 374920 295264 374972 295316
rect 514208 295264 514260 295316
rect 381452 295196 381504 295248
rect 520556 295196 520608 295248
rect 369308 295128 369360 295180
rect 510712 295128 510764 295180
rect 374828 295060 374880 295112
rect 517704 295060 517756 295112
rect 374736 294992 374788 295044
rect 517888 294992 517940 295044
rect 376300 294924 376352 294976
rect 520464 294924 520516 294976
rect 373632 294856 373684 294908
rect 519084 294856 519136 294908
rect 372252 294788 372304 294840
rect 519176 294788 519228 294840
rect 370688 294720 370740 294772
rect 519360 294720 519412 294772
rect 366640 294652 366692 294704
rect 516508 294652 516560 294704
rect 369400 294584 369452 294636
rect 519452 294584 519504 294636
rect 372160 294516 372212 294568
rect 509424 294516 509476 294568
rect 457720 294448 457772 294500
rect 570696 294448 570748 294500
rect 361764 293904 361816 293956
rect 435364 293904 435416 293956
rect 488356 293292 488408 293344
rect 530032 293292 530084 293344
rect 467564 293224 467616 293276
rect 559564 293224 559616 293276
rect 3332 292544 3384 292596
rect 19984 292544 20036 292596
rect 384304 292476 384356 292528
rect 507400 292476 507452 292528
rect 386052 292408 386104 292460
rect 520832 292408 520884 292460
rect 383476 292340 383528 292392
rect 518900 292340 518952 292392
rect 377680 292272 377732 292324
rect 514760 292272 514812 292324
rect 379060 292204 379112 292256
rect 516876 292204 516928 292256
rect 375104 292136 375156 292188
rect 514116 292136 514168 292188
rect 369216 292068 369268 292120
rect 507492 292068 507544 292120
rect 380532 292000 380584 292052
rect 520280 292000 520332 292052
rect 377772 291932 377824 291984
rect 520372 291932 520424 291984
rect 366364 291864 366416 291916
rect 516600 291864 516652 291916
rect 363696 291796 363748 291848
rect 519728 291796 519780 291848
rect 385960 291728 386012 291780
rect 507584 291728 507636 291780
rect 471244 291660 471296 291712
rect 474004 291660 474056 291712
rect 478420 291660 478472 291712
rect 559656 291660 559708 291712
rect 467656 290436 467708 290488
rect 558184 290436 558236 290488
rect 375012 289756 375064 289808
rect 507308 289756 507360 289808
rect 384764 289688 384816 289740
rect 518992 289688 519044 289740
rect 380256 289620 380308 289672
rect 517796 289620 517848 289672
rect 382188 289552 382240 289604
rect 521844 289552 521896 289604
rect 383292 289484 383344 289536
rect 523224 289484 523276 289536
rect 377588 289416 377640 289468
rect 519268 289416 519320 289468
rect 380348 289348 380400 289400
rect 523316 289348 523368 289400
rect 378968 289280 379020 289332
rect 523132 289280 523184 289332
rect 377496 289212 377548 289264
rect 521936 289212 521988 289264
rect 376116 289144 376168 289196
rect 521752 289144 521804 289196
rect 372344 289076 372396 289128
rect 520648 289076 520700 289128
rect 383384 289008 383436 289060
rect 514944 289008 514996 289060
rect 385868 288940 385920 288992
rect 507216 288940 507268 288992
rect 467288 288872 467340 288924
rect 555424 288872 555476 288924
rect 475384 287784 475436 287836
rect 476856 287784 476908 287836
rect 461400 286696 461452 286748
rect 471244 286696 471296 286748
rect 452108 286628 452160 286680
rect 490840 286628 490892 286680
rect 370504 286560 370556 286612
rect 476488 286560 476540 286612
rect 488080 286560 488132 286612
rect 531320 286560 531372 286612
rect 372068 286492 372120 286544
rect 507124 286492 507176 286544
rect 377404 286424 377456 286476
rect 520740 286424 520792 286476
rect 366456 286356 366508 286408
rect 521660 286356 521712 286408
rect 365260 286288 365312 286340
rect 523040 286288 523092 286340
rect 453304 284928 453356 284980
rect 489184 284928 489236 284980
rect 498016 284928 498068 284980
rect 539876 284928 539928 284980
rect 452384 283568 452436 283620
rect 494980 283568 495032 283620
rect 459468 282888 459520 282940
rect 460388 282888 460440 282940
rect 361764 282820 361816 282872
rect 436836 282820 436888 282872
rect 459284 282140 459336 282192
rect 494152 282140 494204 282192
rect 455052 280780 455104 280832
rect 493416 280780 493468 280832
rect 453672 279488 453724 279540
rect 461400 279488 461452 279540
rect 453396 279420 453448 279472
rect 490656 279420 490708 279472
rect 503628 279420 503680 279472
rect 539048 279420 539100 279472
rect 453488 278060 453540 278112
rect 490012 278060 490064 278112
rect 381360 277992 381412 278044
rect 486424 277992 486476 278044
rect 501788 277992 501840 278044
rect 540244 277992 540296 278044
rect 455236 276632 455288 276684
rect 494704 276632 494756 276684
rect 500224 276632 500276 276684
rect 539968 276632 540020 276684
rect 459192 275272 459244 275324
rect 493140 275272 493192 275324
rect 499028 275272 499080 275324
rect 541256 275272 541308 275324
rect 473360 274660 473412 274712
rect 475384 274660 475436 274712
rect 457628 273980 457680 274032
rect 491392 273980 491444 274032
rect 499396 273980 499448 274032
rect 541348 273980 541400 274032
rect 452200 273912 452252 273964
rect 488632 273912 488684 273964
rect 497740 273912 497792 273964
rect 542820 273912 542872 273964
rect 479524 273164 479576 273216
rect 579896 273164 579948 273216
rect 453580 272552 453632 272604
rect 488908 272552 488960 272604
rect 455144 272484 455196 272536
rect 492772 272484 492824 272536
rect 500776 272484 500828 272536
rect 541440 272484 541492 272536
rect 361764 271804 361816 271856
rect 439688 271804 439740 271856
rect 459100 271192 459152 271244
rect 491668 271192 491720 271244
rect 500500 271192 500552 271244
rect 540152 271192 540204 271244
rect 457720 271124 457772 271176
rect 493324 271124 493376 271176
rect 499120 271124 499172 271176
rect 540060 271124 540112 271176
rect 456248 271056 456300 271108
rect 459468 271056 459520 271108
rect 456708 269900 456760 269952
rect 473728 269900 473780 269952
rect 505008 269900 505060 269952
rect 543740 269900 543792 269952
rect 456156 269832 456208 269884
rect 487252 269832 487304 269884
rect 496728 269832 496780 269884
rect 541164 269832 541216 269884
rect 468760 269764 468812 269816
rect 580356 269764 580408 269816
rect 459560 268540 459612 268592
rect 473360 268540 473412 268592
rect 452292 268472 452344 268524
rect 490564 268472 490616 268524
rect 466368 268404 466420 268456
rect 570604 268404 570656 268456
rect 361212 268336 361264 268388
rect 512000 268336 512052 268388
rect 3608 266364 3660 266416
rect 4896 266364 4948 266416
rect 456892 266364 456944 266416
rect 459560 266364 459612 266416
rect 453948 263576 454000 263628
rect 456892 263576 456944 263628
rect 449808 263508 449860 263560
rect 456800 263508 456852 263560
rect 448520 262896 448572 262948
rect 456708 262896 456760 262948
rect 420184 262828 420236 262880
rect 453672 262828 453724 262880
rect 361764 260788 361816 260840
rect 440884 260788 440936 260840
rect 437756 258680 437808 258732
rect 448520 258680 448572 258732
rect 449164 258068 449216 258120
rect 453948 258068 454000 258120
rect 414664 256708 414716 256760
rect 420184 256708 420236 256760
rect 429844 253172 429896 253224
rect 437756 253172 437808 253224
rect 456892 250928 456944 250980
rect 459376 250928 459428 250980
rect 361764 249704 361816 249756
rect 399484 249704 399536 249756
rect 447140 249704 447192 249756
rect 456800 249704 456852 249756
rect 446404 248888 446456 248940
rect 447140 248888 447192 248940
rect 447232 247664 447284 247716
rect 456892 247664 456944 247716
rect 445760 246984 445812 247036
rect 449164 247052 449216 247104
rect 445668 245556 445720 245608
rect 447232 245624 447284 245676
rect 570696 245556 570748 245608
rect 580172 245556 580224 245608
rect 449164 243516 449216 243568
rect 456248 243516 456300 243568
rect 3976 241408 4028 241460
rect 5080 241408 5132 241460
rect 427084 241408 427136 241460
rect 429844 241408 429896 241460
rect 443184 241136 443236 241188
rect 445668 241136 445720 241188
rect 445208 239776 445260 239828
rect 445760 239776 445812 239828
rect 361764 238688 361816 238740
rect 443736 238688 443788 238740
rect 442264 237396 442316 237448
rect 443184 237396 443236 237448
rect 443920 237396 443972 237448
rect 445208 237396 445260 237448
rect 450728 235220 450780 235272
rect 456800 235220 456852 235272
rect 3792 233180 3844 233232
rect 4988 233180 5040 233232
rect 559656 233180 559708 233232
rect 580172 233180 580224 233232
rect 442448 229984 442500 230036
rect 443920 229984 443972 230036
rect 421564 229712 421616 229764
rect 427084 229712 427136 229764
rect 361764 227672 361816 227724
rect 443644 227672 443696 227724
rect 440884 226584 440936 226636
rect 442448 226584 442500 226636
rect 450544 221416 450596 221468
rect 457904 221416 457956 221468
rect 361672 216316 361724 216368
rect 364064 216316 364116 216368
rect 439688 213868 439740 213920
rect 440884 213868 440936 213920
rect 437480 208360 437532 208412
rect 439688 208360 439740 208412
rect 450636 207612 450688 207664
rect 459560 207612 459612 207664
rect 460020 207612 460072 207664
rect 576124 206932 576176 206984
rect 579804 206932 579856 206984
rect 361764 205572 361816 205624
rect 439596 205572 439648 205624
rect 3884 205096 3936 205148
rect 5172 205096 5224 205148
rect 440884 204212 440936 204264
rect 442264 204212 442316 204264
rect 410524 203396 410576 203448
rect 414664 203396 414716 203448
rect 433340 202784 433392 202836
rect 437480 202852 437532 202904
rect 447784 201288 447836 201340
rect 449164 201288 449216 201340
rect 460664 200676 460716 200728
rect 462320 200676 462372 200728
rect 447324 199384 447376 199436
rect 461584 199384 461636 199436
rect 361764 194488 361816 194540
rect 436744 194488 436796 194540
rect 418528 193128 418580 193180
rect 421564 193128 421616 193180
rect 548524 193128 548576 193180
rect 580172 193128 580224 193180
rect 439596 191768 439648 191820
rect 440884 191768 440936 191820
rect 431224 190476 431276 190528
rect 433248 190476 433300 190528
rect 407028 186940 407080 186992
rect 418528 186940 418580 186992
rect 395344 184152 395396 184204
rect 407028 184152 407080 184204
rect 361764 183472 361816 183524
rect 447232 183472 447284 183524
rect 447232 182792 447284 182844
rect 448152 182792 448204 182844
rect 528560 182792 528612 182844
rect 559564 179324 559616 179376
rect 580172 179324 580224 179376
rect 419540 175924 419592 175976
rect 431224 175924 431276 175976
rect 436744 175176 436796 175228
rect 439596 175244 439648 175296
rect 389824 174564 389876 174616
rect 395344 174564 395396 174616
rect 414664 173884 414716 173936
rect 419540 173884 419592 173936
rect 361764 172456 361816 172508
rect 447232 172456 447284 172508
rect 447232 171776 447284 171828
rect 448336 171776 448388 171828
rect 524420 171776 524472 171828
rect 411260 169668 411312 169720
rect 414664 169736 414716 169788
rect 432236 169736 432288 169788
rect 436744 169736 436796 169788
rect 444012 169736 444064 169788
rect 447784 169736 447836 169788
rect 429844 168308 429896 168360
rect 432236 168376 432288 168428
rect 536104 166948 536156 167000
rect 580172 166948 580224 167000
rect 369032 166268 369084 166320
rect 389824 166268 389876 166320
rect 440240 165928 440292 165980
rect 444012 165928 444064 165980
rect 408500 164160 408552 164212
rect 411260 164228 411312 164280
rect 448428 164160 448480 164212
rect 449348 164160 449400 164212
rect 438584 163616 438636 163668
rect 439504 163616 439556 163668
rect 445208 163616 445260 163668
rect 446404 163616 446456 163668
rect 361580 163480 361632 163532
rect 369032 163480 369084 163532
rect 437572 162256 437624 162308
rect 440240 162256 440292 162308
rect 418712 162188 418764 162240
rect 457812 162188 457864 162240
rect 489920 162188 489972 162240
rect 415124 162120 415176 162172
rect 457904 162120 457956 162172
rect 485780 162120 485832 162172
rect 445208 161576 445260 161628
rect 450544 161576 450596 161628
rect 375196 161508 375248 161560
rect 418712 161508 418764 161560
rect 431868 161508 431920 161560
rect 450636 161508 450688 161560
rect 412088 161440 412140 161492
rect 459560 161440 459612 161492
rect 460388 161440 460440 161492
rect 361764 161372 361816 161424
rect 448336 161372 448388 161424
rect 448336 160692 448388 160744
rect 521660 160692 521712 160744
rect 425336 160420 425388 160472
rect 425888 160420 425940 160472
rect 496820 160420 496872 160472
rect 428648 160352 428700 160404
rect 500960 160352 501012 160404
rect 421840 160284 421892 160336
rect 494060 160284 494112 160336
rect 435272 160216 435324 160268
rect 436008 160216 436060 160268
rect 509240 160216 509292 160268
rect 386144 160148 386196 160200
rect 415124 160148 415176 160200
rect 427820 160148 427872 160200
rect 429844 160148 429896 160200
rect 438584 160148 438636 160200
rect 513380 160148 513432 160200
rect 409512 160080 409564 160132
rect 441574 160080 441626 160132
rect 442908 160080 442960 160132
rect 517520 160080 517572 160132
rect 401600 159808 401652 159860
rect 408500 159808 408552 159860
rect 409420 159740 409472 159792
rect 427820 159740 427872 159792
rect 409144 159672 409196 159724
rect 428004 159672 428056 159724
rect 409236 159604 409288 159656
rect 434812 159604 434864 159656
rect 409328 159536 409380 159588
rect 437940 159536 437992 159588
rect 406108 159468 406160 159520
rect 437572 159468 437624 159520
rect 384212 159400 384264 159452
rect 421380 159400 421432 159452
rect 386236 159332 386288 159384
rect 425152 159332 425204 159384
rect 451740 158244 451792 158296
rect 456156 158244 456208 158296
rect 404268 157496 404320 157548
rect 406108 157496 406160 157548
rect 451740 157292 451792 157344
rect 457536 157292 457588 157344
rect 400864 156612 400916 156664
rect 410524 156612 410576 156664
rect 396724 156136 396776 156188
rect 404268 156136 404320 156188
rect 359464 155320 359516 155372
rect 361580 155320 361632 155372
rect 451924 154164 451976 154216
rect 455236 154164 455288 154216
rect 396908 153144 396960 153196
rect 401600 153212 401652 153264
rect 547144 153144 547196 153196
rect 580172 153144 580224 153196
rect 395160 150424 395212 150476
rect 396908 150424 396960 150476
rect 361764 150356 361816 150408
rect 409512 150356 409564 150408
rect 452476 150220 452528 150272
rect 459284 150220 459336 150272
rect 452568 148724 452620 148776
rect 454960 148724 455012 148776
rect 391204 147636 391256 147688
rect 395160 147636 395212 147688
rect 407120 147636 407172 147688
rect 409420 147636 409472 147688
rect 451740 147364 451792 147416
rect 457720 147364 457772 147416
rect 452568 146004 452620 146056
rect 459008 146004 459060 146056
rect 396816 145120 396868 145172
rect 400864 145120 400916 145172
rect 404820 145120 404872 145172
rect 407120 145120 407172 145172
rect 451464 144780 451516 144832
rect 455052 144780 455104 144832
rect 460388 143488 460440 143540
rect 460848 143488 460900 143540
rect 533436 143488 533488 143540
rect 537300 143488 537352 143540
rect 452568 143284 452620 143336
rect 459192 143284 459244 143336
rect 460848 142264 460900 142316
rect 481916 142264 481968 142316
rect 450636 142196 450688 142248
rect 505652 142196 505704 142248
rect 401600 142128 401652 142180
rect 404820 142128 404872 142180
rect 450544 142128 450596 142180
rect 533988 142128 534040 142180
rect 540336 142196 540388 142248
rect 452568 141924 452620 141976
rect 455144 141924 455196 141976
rect 452568 140564 452620 140616
rect 457628 140564 457680 140616
rect 534724 140088 534776 140140
rect 542912 140088 542964 140140
rect 533344 140020 533396 140072
rect 543188 140020 543240 140072
rect 361764 139340 361816 139392
rect 409328 139340 409380 139392
rect 555424 139340 555476 139392
rect 580172 139340 580224 139392
rect 452568 139204 452620 139256
rect 459100 139204 459152 139256
rect 538864 138592 538916 138644
rect 543096 138592 543148 138644
rect 452568 137844 452620 137896
rect 454776 137844 454828 137896
rect 389456 137300 389508 137352
rect 391204 137300 391256 137352
rect 388444 137232 388496 137284
rect 396816 137232 396868 137284
rect 394700 136620 394752 136672
rect 396724 136620 396776 136672
rect 538956 136552 539008 136604
rect 539508 136552 539560 136604
rect 452568 136484 452620 136536
rect 457444 136484 457496 136536
rect 391204 135872 391256 135924
rect 401508 135872 401560 135924
rect 387800 135192 387852 135244
rect 389456 135192 389508 135244
rect 452568 135124 452620 135176
rect 458916 135124 458968 135176
rect 452568 133764 452620 133816
rect 454868 133764 454920 133816
rect 391940 132404 391992 132456
rect 394700 132472 394752 132524
rect 452292 131044 452344 131096
rect 453396 131044 453448 131096
rect 389180 129820 389232 129872
rect 391204 129820 391256 129872
rect 387064 129752 387116 129804
rect 391940 129752 391992 129804
rect 452384 129684 452436 129736
rect 453488 129684 453540 129736
rect 359556 129004 359608 129056
rect 388444 129004 388496 129056
rect 361764 128256 361816 128308
rect 409236 128256 409288 128308
rect 452292 126896 452344 126948
rect 453304 126896 453356 126948
rect 573364 126896 573416 126948
rect 580172 126896 580224 126948
rect 451740 126352 451792 126404
rect 453580 126352 453632 126404
rect 368296 126216 368348 126268
rect 387708 126216 387760 126268
rect 362960 124856 363012 124908
rect 389088 124856 389140 124908
rect 451832 124108 451884 124160
rect 458824 124108 458876 124160
rect 451740 122204 451792 122256
rect 454684 122204 454736 122256
rect 371240 122068 371292 122120
rect 387064 122068 387116 122120
rect 384948 119348 385000 119400
rect 456064 119348 456116 119400
rect 361304 118668 361356 118720
rect 362868 118668 362920 118720
rect 366916 118600 366968 118652
rect 371240 118668 371292 118720
rect 362592 117920 362644 117972
rect 368296 117920 368348 117972
rect 361764 117240 361816 117292
rect 450636 117240 450688 117292
rect 364064 116832 364116 116884
rect 366916 116832 366968 116884
rect 569224 113092 569276 113144
rect 579804 113092 579856 113144
rect 361396 111800 361448 111852
rect 364064 111800 364116 111852
rect 389824 106904 389876 106956
rect 450544 106904 450596 106956
rect 361764 106224 361816 106276
rect 409144 106224 409196 106276
rect 558184 100648 558236 100700
rect 580172 100648 580224 100700
rect 361764 95140 361816 95192
rect 386236 95140 386288 95192
rect 571984 86912 572036 86964
rect 580172 86912 580224 86964
rect 3148 84192 3200 84244
rect 20904 84192 20956 84244
rect 361764 84124 361816 84176
rect 384212 84124 384264 84176
rect 5080 80044 5132 80096
rect 8576 79976 8628 80028
rect 8576 78480 8628 78532
rect 10324 78480 10376 78532
rect 361764 73108 361816 73160
rect 375196 73108 375248 73160
rect 544384 73108 544436 73160
rect 580172 73108 580224 73160
rect 3148 70388 3200 70440
rect 20076 70388 20128 70440
rect 5172 68960 5224 69012
rect 7564 68960 7616 69012
rect 4896 68892 4948 68944
rect 5540 68892 5592 68944
rect 5540 66240 5592 66292
rect 8300 66172 8352 66224
rect 10324 63860 10376 63912
rect 12072 63860 12124 63912
rect 8300 62636 8352 62688
rect 10416 62636 10468 62688
rect 361764 62024 361816 62076
rect 386144 62024 386196 62076
rect 7564 60664 7616 60716
rect 9588 60664 9640 60716
rect 551284 60664 551336 60716
rect 580172 60664 580224 60716
rect 3424 59984 3476 60036
rect 20904 59984 20956 60036
rect 4804 59304 4856 59356
rect 7564 59304 7616 59356
rect 4988 57876 5040 57928
rect 5540 57876 5592 57928
rect 7564 56584 7616 56636
rect 10784 56516 10836 56568
rect 12072 56516 12124 56568
rect 13728 56516 13780 56568
rect 10416 56448 10468 56500
rect 12440 56448 12492 56500
rect 9680 56380 9732 56432
rect 17960 56516 18012 56568
rect 10784 54612 10836 54664
rect 13636 54612 13688 54664
rect 5540 54476 5592 54528
rect 11704 54476 11756 54528
rect 17960 54068 18012 54120
rect 20628 54068 20680 54120
rect 13728 52980 13780 53032
rect 15200 52980 15252 53032
rect 12440 52708 12492 52760
rect 14556 52708 14608 52760
rect 13636 52436 13688 52488
rect 19248 52368 19300 52420
rect 11704 51076 11756 51128
rect 361764 51076 361816 51128
rect 386144 51076 386196 51128
rect 540612 51076 540664 51128
rect 543740 51076 543792 51128
rect 15292 51008 15344 51060
rect 15200 49648 15252 49700
rect 16856 49648 16908 49700
rect 16856 48152 16908 48204
rect 20812 48152 20864 48204
rect 15292 47268 15344 47320
rect 19248 47268 19300 47320
rect 3240 46996 3292 47048
rect 384856 46996 384908 47048
rect 3332 46860 3384 46912
rect 381820 46860 381872 46912
rect 574744 46860 574796 46912
rect 580172 46860 580224 46912
rect 4068 46792 4120 46844
rect 382004 46792 382056 46844
rect 3792 46724 3844 46776
rect 378876 46724 378928 46776
rect 3700 46656 3752 46708
rect 378600 46656 378652 46708
rect 3608 46588 3660 46640
rect 376668 46588 376720 46640
rect 3516 46520 3568 46572
rect 375932 46520 375984 46572
rect 20076 46452 20128 46504
rect 384580 46452 384632 46504
rect 21364 46384 21416 46436
rect 384488 46384 384540 46436
rect 19984 46316 20036 46368
rect 375840 46316 375892 46368
rect 14556 46248 14608 46300
rect 359556 46248 359608 46300
rect 19248 46180 19300 46232
rect 362592 46180 362644 46232
rect 20812 46112 20864 46164
rect 361396 46112 361448 46164
rect 20720 46044 20772 46096
rect 361304 46044 361356 46096
rect 3516 45500 3568 45552
rect 381360 45500 381412 45552
rect 3976 45432 4028 45484
rect 381636 45432 381688 45484
rect 3884 45364 3936 45416
rect 378784 45364 378836 45416
rect 21456 45296 21508 45348
rect 373724 45296 373776 45348
rect 65524 45228 65576 45280
rect 379428 45228 379480 45280
rect 62028 45160 62080 45212
rect 378692 45160 378744 45212
rect 58440 45092 58492 45144
rect 379244 45092 379296 45144
rect 54944 45024 54996 45076
rect 379336 45024 379388 45076
rect 51356 44956 51408 45008
rect 379152 44956 379204 45008
rect 47860 44888 47912 44940
rect 381912 44888 381964 44940
rect 7656 44820 7708 44872
rect 382096 44820 382148 44872
rect 69112 44752 69164 44804
rect 376576 44752 376628 44804
rect 72608 44684 72660 44736
rect 376392 44684 376444 44736
rect 76196 44616 76248 44668
rect 376484 44616 376536 44668
rect 111616 42712 111668 42764
rect 368204 42712 368256 42764
rect 108120 42644 108172 42696
rect 368020 42644 368072 42696
rect 104532 42576 104584 42628
rect 370780 42576 370832 42628
rect 101036 42508 101088 42560
rect 370596 42508 370648 42560
rect 97448 42440 97500 42492
rect 370872 42440 370924 42492
rect 93952 42372 94004 42424
rect 370964 42372 371016 42424
rect 90364 42304 90416 42356
rect 373540 42304 373592 42356
rect 86868 42236 86920 42288
rect 373448 42236 373500 42288
rect 83280 42168 83332 42220
rect 373356 42168 373408 42220
rect 79692 42100 79744 42152
rect 376024 42100 376076 42152
rect 12348 42032 12400 42084
rect 376208 42032 376260 42084
rect 115204 41964 115256 42016
rect 367928 41964 367980 42016
rect 461584 41352 461636 41404
rect 536840 41352 536892 41404
rect 118792 39992 118844 40044
rect 365444 39992 365496 40044
rect 63224 39924 63276 39976
rect 369400 39924 369452 39976
rect 59636 39856 59688 39908
rect 366640 39856 366692 39908
rect 56048 39788 56100 39840
rect 368112 39788 368164 39840
rect 52552 39720 52604 39772
rect 366548 39720 366600 39772
rect 48964 39652 49016 39704
rect 363880 39652 363932 39704
rect 40684 39584 40736 39636
rect 363788 39584 363840 39636
rect 37188 39516 37240 39568
rect 362500 39516 362552 39568
rect 33600 39448 33652 39500
rect 363972 39448 364024 39500
rect 26516 39380 26568 39432
rect 362408 39380 362460 39432
rect 4068 39312 4120 39364
rect 365352 39312 365404 39364
rect 122288 39244 122340 39296
rect 365168 39244 365220 39296
rect 102232 37204 102284 37256
rect 375104 37204 375156 37256
rect 98644 37136 98696 37188
rect 374920 37136 374972 37188
rect 95148 37068 95200 37120
rect 376300 37068 376352 37120
rect 87972 37000 88024 37052
rect 374828 37000 374880 37052
rect 91560 36932 91612 36984
rect 381452 36932 381504 36984
rect 84476 36864 84528 36916
rect 374736 36864 374788 36916
rect 80888 36796 80940 36848
rect 373632 36796 373684 36848
rect 77392 36728 77444 36780
rect 372160 36728 372212 36780
rect 73804 36660 73856 36712
rect 372252 36660 372304 36712
rect 70308 36592 70360 36644
rect 369308 36592 369360 36644
rect 66720 36524 66772 36576
rect 370688 36524 370740 36576
rect 105728 36456 105780 36508
rect 377772 36456 377824 36508
rect 119896 34416 119948 34468
rect 383476 34416 383528 34468
rect 116400 34348 116452 34400
rect 380532 34348 380584 34400
rect 112812 34280 112864 34332
rect 377680 34280 377732 34332
rect 109316 34212 109368 34264
rect 379060 34212 379112 34264
rect 50160 34144 50212 34196
rect 375012 34144 375064 34196
rect 45468 34076 45520 34128
rect 372344 34076 372396 34128
rect 41880 34008 41932 34060
rect 369216 34008 369268 34060
rect 34796 33940 34848 33992
rect 363696 33940 363748 33992
rect 31300 33872 31352 33924
rect 386052 33872 386104 33924
rect 18236 33804 18288 33856
rect 380440 33804 380492 33856
rect 23020 33736 23072 33788
rect 385960 33736 386012 33788
rect 123484 33668 123536 33720
rect 382924 33668 382976 33720
rect 2872 33056 2924 33108
rect 383200 33056 383252 33108
rect 566464 33056 566516 33108
rect 580172 33056 580224 33108
rect 3424 31696 3476 31748
rect 460296 31696 460348 31748
rect 96252 31628 96304 31680
rect 378968 31628 379020 31680
rect 386144 31628 386196 31680
rect 460388 31628 460440 31680
rect 92756 31560 92808 31612
rect 382188 31560 382240 31612
rect 85672 31492 85724 31544
rect 384764 31492 384816 31544
rect 78588 31424 78640 31476
rect 383292 31424 383344 31476
rect 71504 31356 71556 31408
rect 380256 31356 380308 31408
rect 67916 31288 67968 31340
rect 377496 31288 377548 31340
rect 64328 31220 64380 31272
rect 383384 31220 383436 31272
rect 60832 31152 60884 31204
rect 380348 31152 380400 31204
rect 57244 31084 57296 31136
rect 377588 31084 377640 31136
rect 14740 31016 14792 31068
rect 385868 31016 385920 31068
rect 99840 30948 99892 31000
rect 376116 30948 376168 31000
rect 117596 28908 117648 28960
rect 369124 28908 369176 28960
rect 121092 28840 121144 28892
rect 373264 28840 373316 28892
rect 114008 28772 114060 28824
rect 366456 28772 366508 28824
rect 106924 28704 106976 28756
rect 365260 28704 365312 28756
rect 35992 28636 36044 28688
rect 383108 28636 383160 28688
rect 32404 28568 32456 28620
rect 380164 28568 380216 28620
rect 28908 28500 28960 28552
rect 377404 28500 377456 28552
rect 109684 28432 109736 28484
rect 460940 28432 460992 28484
rect 19432 28364 19484 28416
rect 372068 28364 372120 28416
rect 5264 28296 5316 28348
rect 384948 28296 385000 28348
rect 43076 28228 43128 28280
rect 462320 28228 462372 28280
rect 124680 28160 124732 28212
rect 374644 28160 374696 28212
rect 3424 20612 3476 20664
rect 370504 20612 370556 20664
rect 570604 20612 570656 20664
rect 579988 20612 580040 20664
rect 3424 6808 3476 6860
rect 371884 6808 371936 6860
rect 562324 6808 562376 6860
rect 580172 6808 580224 6860
rect 82084 4088 82136 4140
rect 367744 4088 367796 4140
rect 75000 4020 75052 4072
rect 367836 4020 367888 4072
rect 53748 3952 53800 4004
rect 364984 3952 365036 4004
rect 46664 3884 46716 3936
rect 363604 3884 363656 3936
rect 39580 3816 39632 3868
rect 361212 3816 361264 3868
rect 38384 3748 38436 3800
rect 366364 3748 366416 3800
rect 30104 3680 30156 3732
rect 360936 3680 360988 3732
rect 44272 3612 44324 3664
rect 383016 3612 383068 3664
rect 21824 3544 21876 3596
rect 362316 3544 362368 3596
rect 27712 3476 27764 3528
rect 384304 3476 384356 3528
rect 24216 3408 24268 3460
rect 385684 3408 385736 3460
rect 89168 3340 89220 3392
rect 361120 3340 361172 3392
rect 103336 3272 103388 3324
rect 361028 3272 361080 3324
rect 6460 3204 6512 3256
rect 109684 3204 109736 3256
rect 110512 3204 110564 3256
rect 360844 3204 360896 3256
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 686526 8156 703520
rect 24320 689353 24348 703520
rect 40512 700330 40540 703520
rect 40500 700324 40552 700330
rect 40500 700266 40552 700272
rect 24306 689344 24362 689353
rect 24306 689279 24362 689288
rect 8116 686520 8168 686526
rect 8116 686462 8168 686468
rect 72988 685166 73016 703520
rect 89180 685234 89208 703520
rect 105464 700369 105492 703520
rect 137848 700505 137876 703520
rect 137834 700496 137890 700505
rect 154132 700466 154160 703520
rect 137834 700431 137890 700440
rect 154120 700460 154172 700466
rect 154120 700402 154172 700408
rect 170324 700398 170352 703520
rect 202800 700534 202828 703520
rect 218992 700670 219020 703520
rect 218980 700664 219032 700670
rect 218980 700606 219032 700612
rect 235184 700602 235212 703520
rect 235172 700596 235224 700602
rect 235172 700538 235224 700544
rect 202788 700528 202840 700534
rect 202788 700470 202840 700476
rect 170312 700392 170364 700398
rect 105450 700360 105506 700369
rect 170312 700334 170364 700340
rect 105450 700295 105506 700304
rect 267660 685302 267688 703520
rect 283852 692073 283880 703520
rect 283838 692064 283894 692073
rect 283838 691999 283894 692008
rect 300136 690674 300164 703520
rect 332520 700738 332548 703520
rect 332508 700732 332560 700738
rect 332508 700674 332560 700680
rect 300124 690668 300176 690674
rect 300124 690610 300176 690616
rect 348804 687954 348832 703520
rect 364996 700806 365024 703520
rect 397472 700874 397500 703520
rect 397460 700868 397512 700874
rect 397460 700810 397512 700816
rect 364984 700800 365036 700806
rect 364984 700742 365036 700748
rect 348792 687948 348844 687954
rect 348792 687890 348844 687896
rect 267648 685296 267700 685302
rect 267648 685238 267700 685244
rect 89168 685228 89220 685234
rect 89168 685170 89220 685176
rect 72976 685160 73028 685166
rect 72976 685102 73028 685108
rect 3792 684684 3844 684690
rect 3792 684626 3844 684632
rect 3424 684616 3476 684622
rect 3424 684558 3476 684564
rect 3332 683392 3384 683398
rect 3332 683334 3384 683340
rect 3240 682712 3292 682718
rect 3240 682654 3292 682660
rect 3148 633412 3200 633418
rect 3148 633354 3200 633360
rect 3160 632097 3188 633354
rect 3146 632088 3202 632097
rect 3146 632023 3202 632032
rect 3252 580009 3280 682654
rect 3238 580000 3294 580009
rect 3238 579935 3294 579944
rect 3344 566953 3372 683334
rect 3330 566944 3386 566953
rect 3330 566879 3386 566888
rect 3436 449585 3464 684558
rect 3608 683528 3660 683534
rect 3608 683470 3660 683476
rect 3516 683256 3568 683262
rect 3516 683198 3568 683204
rect 3528 658209 3556 683198
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3516 656192 3568 656198
rect 3516 656134 3568 656140
rect 3422 449576 3478 449585
rect 3422 449511 3478 449520
rect 3528 423609 3556 656134
rect 3620 462641 3648 683470
rect 3700 683460 3752 683466
rect 3700 683402 3752 683408
rect 3712 475697 3740 683402
rect 3804 501809 3832 684626
rect 3976 684548 4028 684554
rect 3976 684490 4028 684496
rect 3884 683596 3936 683602
rect 3884 683538 3936 683544
rect 3896 514865 3924 683538
rect 3988 527921 4016 684490
rect 24124 683732 24176 683738
rect 24124 683674 24176 683680
rect 359464 683732 359516 683738
rect 359464 683674 359516 683680
rect 21456 683664 21508 683670
rect 21456 683606 21508 683612
rect 21364 683324 21416 683330
rect 21364 683266 21416 683272
rect 4068 683188 4120 683194
rect 4068 683130 4120 683136
rect 4080 553897 4108 683130
rect 11060 682780 11112 682786
rect 11060 682722 11112 682728
rect 11072 680354 11100 682722
rect 10980 680326 11100 680354
rect 10980 675850 11008 680326
rect 6920 675844 6972 675850
rect 6920 675786 6972 675792
rect 10968 675844 11020 675850
rect 10968 675786 11020 675792
rect 6932 670698 6960 675786
rect 6840 670670 6960 670698
rect 6840 667962 6868 670670
rect 4804 667956 4856 667962
rect 4804 667898 4856 667904
rect 6828 667956 6880 667962
rect 6828 667898 6880 667904
rect 4066 553888 4122 553897
rect 4066 553823 4122 553832
rect 3974 527912 4030 527921
rect 3974 527847 4030 527856
rect 3882 514856 3938 514865
rect 4816 514826 4844 667898
rect 21376 663794 21404 683266
rect 21284 663766 21404 663794
rect 20902 656296 20958 656305
rect 20902 656231 20958 656240
rect 20916 656198 20944 656231
rect 20904 656192 20956 656198
rect 20904 656134 20956 656140
rect 21284 654134 21312 663766
rect 21468 656305 21496 683606
rect 24136 682786 24164 683674
rect 24124 682780 24176 682786
rect 24124 682722 24176 682728
rect 359476 672110 359504 683674
rect 362222 679008 362278 679017
rect 362222 678943 362278 678952
rect 359464 672104 359516 672110
rect 359464 672046 359516 672052
rect 360844 672104 360896 672110
rect 360844 672046 360896 672052
rect 21454 656296 21510 656305
rect 21454 656231 21510 656240
rect 21284 654106 21404 654134
rect 21376 634814 21404 654106
rect 20916 634786 21404 634814
rect 20916 633418 20944 634786
rect 20904 633412 20956 633418
rect 20904 633354 20956 633360
rect 360856 602342 360884 672046
rect 361762 667992 361818 668001
rect 361762 667927 361764 667936
rect 361816 667927 361818 667936
rect 361764 667898 361816 667904
rect 361762 656976 361818 656985
rect 361762 656911 361764 656920
rect 361816 656911 361818 656920
rect 361764 656882 361816 656888
rect 361762 645960 361818 645969
rect 361762 645895 361764 645904
rect 361816 645895 361818 645904
rect 361764 645866 361816 645872
rect 361578 634944 361634 634953
rect 361578 634879 361634 634888
rect 361592 634846 361620 634879
rect 361580 634840 361632 634846
rect 361580 634782 361632 634788
rect 361578 623928 361634 623937
rect 361578 623863 361634 623872
rect 361592 623830 361620 623863
rect 361580 623824 361632 623830
rect 361580 623766 361632 623772
rect 361578 612912 361634 612921
rect 361578 612847 361580 612856
rect 361632 612847 361634 612856
rect 361580 612818 361632 612824
rect 360844 602336 360896 602342
rect 360844 602278 360896 602284
rect 361762 601896 361818 601905
rect 361762 601831 361818 601840
rect 361776 601730 361804 601831
rect 361764 601724 361816 601730
rect 361764 601666 361816 601672
rect 361578 590880 361634 590889
rect 361578 590815 361580 590824
rect 361632 590815 361634 590824
rect 361580 590786 361632 590792
rect 361762 579864 361818 579873
rect 361762 579799 361818 579808
rect 361776 579698 361804 579799
rect 361764 579692 361816 579698
rect 361764 579634 361816 579640
rect 361578 568848 361634 568857
rect 361578 568783 361580 568792
rect 361632 568783 361634 568792
rect 361580 568754 361632 568760
rect 361670 557832 361726 557841
rect 361670 557767 361726 557776
rect 361684 557598 361712 557767
rect 361672 557592 361724 557598
rect 361672 557534 361724 557540
rect 361762 546816 361818 546825
rect 361762 546751 361818 546760
rect 361776 546514 361804 546751
rect 361764 546508 361816 546514
rect 361764 546450 361816 546456
rect 361762 535800 361818 535809
rect 361762 535735 361818 535744
rect 361776 535498 361804 535735
rect 361764 535492 361816 535498
rect 361764 535434 361816 535440
rect 361762 524784 361818 524793
rect 361762 524719 361818 524728
rect 361776 524482 361804 524719
rect 361764 524476 361816 524482
rect 361764 524418 361816 524424
rect 3882 514791 3938 514800
rect 3976 514820 4028 514826
rect 3976 514762 4028 514768
rect 4804 514820 4856 514826
rect 4804 514762 4856 514768
rect 3790 501800 3846 501809
rect 3790 501735 3846 501744
rect 3698 475688 3754 475697
rect 3698 475623 3754 475632
rect 3606 462632 3662 462641
rect 3606 462567 3662 462576
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3988 410553 4016 514762
rect 361762 513768 361818 513777
rect 361762 513703 361818 513712
rect 361776 513398 361804 513703
rect 361764 513392 361816 513398
rect 361764 513334 361816 513340
rect 361762 502752 361818 502761
rect 361762 502687 361818 502696
rect 361776 502382 361804 502687
rect 361764 502376 361816 502382
rect 361764 502318 361816 502324
rect 361762 491736 361818 491745
rect 361762 491671 361818 491680
rect 361776 491366 361804 491671
rect 361764 491360 361816 491366
rect 361764 491302 361816 491308
rect 361762 480720 361818 480729
rect 361762 480655 361818 480664
rect 361776 480282 361804 480655
rect 361764 480276 361816 480282
rect 361764 480218 361816 480224
rect 361762 469704 361818 469713
rect 361762 469639 361818 469648
rect 361776 469266 361804 469639
rect 361764 469260 361816 469266
rect 361764 469202 361816 469208
rect 361762 458688 361818 458697
rect 361762 458623 361818 458632
rect 361776 458250 361804 458623
rect 361764 458244 361816 458250
rect 361764 458186 361816 458192
rect 361762 447672 361818 447681
rect 361762 447607 361818 447616
rect 361776 447166 361804 447607
rect 361764 447160 361816 447166
rect 361764 447102 361816 447108
rect 361762 436656 361818 436665
rect 361762 436591 361818 436600
rect 361776 436150 361804 436591
rect 361764 436144 361816 436150
rect 361764 436086 361816 436092
rect 361762 425640 361818 425649
rect 361762 425575 361818 425584
rect 361776 425134 361804 425575
rect 361764 425128 361816 425134
rect 361764 425070 361816 425076
rect 361578 414624 361634 414633
rect 361578 414559 361634 414568
rect 361592 414050 361620 414559
rect 361580 414044 361632 414050
rect 361580 413986 361632 413992
rect 3974 410544 4030 410553
rect 3974 410479 4030 410488
rect 361578 403608 361634 403617
rect 361578 403543 361634 403552
rect 361592 403034 361620 403543
rect 361580 403028 361632 403034
rect 361580 402970 361632 402976
rect 3790 397488 3846 397497
rect 3790 397423 3846 397432
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 3436 307766 3464 358391
rect 3606 345400 3662 345409
rect 3606 345335 3662 345344
rect 3424 307760 3476 307766
rect 3424 307702 3476 307708
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 3344 292602 3372 293111
rect 3332 292596 3384 292602
rect 3332 292538 3384 292544
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3160 84250 3188 84623
rect 3148 84244 3200 84250
rect 3148 84186 3200 84192
rect 3146 71632 3202 71641
rect 3146 71567 3202 71576
rect 3160 70446 3188 71567
rect 3148 70440 3200 70446
rect 3148 70382 3200 70388
rect 3252 47054 3280 136711
rect 3240 47048 3292 47054
rect 3240 46990 3292 46996
rect 3344 46918 3372 149767
rect 3436 60042 3464 306167
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3424 60036 3476 60042
rect 3424 59978 3476 59984
rect 3422 58576 3478 58585
rect 3422 58511 3478 58520
rect 3332 46912 3384 46918
rect 3332 46854 3384 46860
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 3436 31754 3464 58511
rect 3528 46578 3556 267135
rect 3620 266422 3648 345335
rect 3608 266416 3660 266422
rect 3608 266358 3660 266364
rect 3606 254144 3662 254153
rect 3606 254079 3662 254088
rect 3620 46646 3648 254079
rect 3698 241088 3754 241097
rect 3698 241023 3754 241032
rect 3712 46714 3740 241023
rect 3804 233238 3832 397423
rect 361578 392592 361634 392601
rect 361578 392527 361634 392536
rect 361592 392018 361620 392527
rect 361580 392012 361632 392018
rect 361580 391954 361632 391960
rect 362236 383654 362264 678943
rect 378784 667956 378836 667962
rect 378784 667898 378836 667904
rect 376024 656940 376076 656946
rect 376024 656882 376076 656888
rect 374736 645924 374788 645930
rect 374736 645866 374788 645872
rect 371884 623824 371936 623830
rect 371884 623766 371936 623772
rect 363604 612876 363656 612882
rect 363604 612818 363656 612824
rect 362960 602336 363012 602342
rect 362960 602278 363012 602284
rect 362972 598398 363000 602278
rect 362960 598392 363012 598398
rect 362960 598334 363012 598340
rect 362224 383648 362276 383654
rect 362224 383590 362276 383596
rect 361578 381576 361634 381585
rect 361578 381511 361634 381520
rect 361592 380934 361620 381511
rect 361580 380928 361632 380934
rect 361580 380870 361632 380876
rect 363616 380866 363644 612818
rect 370504 601724 370556 601730
rect 370504 601666 370556 601672
rect 365444 598392 365496 598398
rect 365444 598334 365496 598340
rect 363696 590844 363748 590850
rect 363696 590786 363748 590792
rect 363604 380860 363656 380866
rect 363604 380802 363656 380808
rect 363708 379506 363736 590786
rect 365456 590646 365484 598334
rect 365444 590640 365496 590646
rect 365444 590582 365496 590588
rect 367744 590640 367796 590646
rect 367744 590582 367796 590588
rect 367756 582894 367784 590582
rect 367744 582888 367796 582894
rect 367744 582830 367796 582836
rect 367744 579692 367796 579698
rect 367744 579634 367796 579640
rect 363788 568812 363840 568818
rect 363788 568754 363840 568760
rect 363696 379500 363748 379506
rect 363696 379442 363748 379448
rect 363800 378146 363828 568754
rect 363788 378140 363840 378146
rect 363788 378082 363840 378088
rect 367756 378078 367784 579634
rect 369124 386436 369176 386442
rect 369124 386378 369176 386384
rect 367744 378072 367796 378078
rect 367744 378014 367796 378020
rect 3882 371376 3938 371385
rect 3882 371311 3938 371320
rect 3792 233232 3844 233238
rect 3792 233174 3844 233180
rect 3790 214976 3846 214985
rect 3790 214911 3846 214920
rect 3804 46782 3832 214911
rect 3896 205154 3924 371311
rect 361578 370560 361634 370569
rect 361578 370495 361634 370504
rect 361592 369918 361620 370495
rect 361580 369912 361632 369918
rect 361580 369854 361632 369860
rect 362222 359544 362278 359553
rect 362222 359479 362278 359488
rect 361762 348528 361818 348537
rect 361762 348463 361818 348472
rect 361776 347818 361804 348463
rect 361764 347812 361816 347818
rect 361764 347754 361816 347760
rect 362236 347750 362264 359479
rect 362224 347744 362276 347750
rect 362224 347686 362276 347692
rect 361764 340944 361816 340950
rect 361764 340886 361816 340892
rect 361776 337521 361804 340886
rect 361762 337512 361818 337521
rect 361762 337447 361818 337456
rect 362224 336048 362276 336054
rect 362224 335990 362276 335996
rect 362236 326505 362264 335990
rect 364064 334008 364116 334014
rect 364064 333950 364116 333956
rect 362222 326496 362278 326505
rect 362222 326431 362278 326440
rect 3974 319288 4030 319297
rect 3974 319223 4030 319232
rect 3988 241466 4016 319223
rect 361764 315988 361816 315994
rect 361764 315930 361816 315936
rect 361776 315489 361804 315930
rect 361762 315480 361818 315489
rect 361762 315415 361818 315424
rect 4804 307760 4856 307766
rect 4804 307702 4856 307708
rect 3976 241460 4028 241466
rect 3976 241402 4028 241408
rect 3884 205148 3936 205154
rect 3884 205090 3936 205096
rect 3882 201920 3938 201929
rect 3882 201855 3938 201864
rect 3792 46776 3844 46782
rect 3792 46718 3844 46724
rect 3700 46708 3752 46714
rect 3700 46650 3752 46656
rect 3608 46640 3660 46646
rect 3608 46582 3660 46588
rect 3516 46572 3568 46578
rect 3516 46514 3568 46520
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 3896 45422 3924 201855
rect 3974 188864 4030 188873
rect 3974 188799 4030 188808
rect 3988 45490 4016 188799
rect 4066 162888 4122 162897
rect 4066 162823 4122 162832
rect 4080 46850 4108 162823
rect 4816 59362 4844 307702
rect 360844 305652 360896 305658
rect 360844 305594 360896 305600
rect 19984 292596 20036 292602
rect 19984 292538 20036 292544
rect 4896 266416 4948 266422
rect 4896 266358 4948 266364
rect 4908 68950 4936 266358
rect 5080 241460 5132 241466
rect 5080 241402 5132 241408
rect 4988 233232 5040 233238
rect 4988 233174 5040 233180
rect 4896 68944 4948 68950
rect 4896 68886 4948 68892
rect 4804 59356 4856 59362
rect 4804 59298 4856 59304
rect 5000 57934 5028 233174
rect 5092 80102 5120 241402
rect 5172 205148 5224 205154
rect 5172 205090 5224 205096
rect 5080 80096 5132 80102
rect 5080 80038 5132 80044
rect 5184 69018 5212 205090
rect 8576 80028 8628 80034
rect 8576 79970 8628 79976
rect 8588 78538 8616 79970
rect 8576 78532 8628 78538
rect 8576 78474 8628 78480
rect 10324 78532 10376 78538
rect 10324 78474 10376 78480
rect 5172 69012 5224 69018
rect 5172 68954 5224 68960
rect 7564 69012 7616 69018
rect 7564 68954 7616 68960
rect 5540 68944 5592 68950
rect 5540 68886 5592 68892
rect 5552 66298 5580 68886
rect 5540 66292 5592 66298
rect 5540 66234 5592 66240
rect 7576 60722 7604 68954
rect 8300 66224 8352 66230
rect 8300 66166 8352 66172
rect 8312 62694 8340 66166
rect 10336 63918 10364 78474
rect 10324 63912 10376 63918
rect 10324 63854 10376 63860
rect 12072 63912 12124 63918
rect 12072 63854 12124 63860
rect 8300 62688 8352 62694
rect 8300 62630 8352 62636
rect 10416 62688 10468 62694
rect 10416 62630 10468 62636
rect 7564 60716 7616 60722
rect 7564 60658 7616 60664
rect 9588 60716 9640 60722
rect 9588 60658 9640 60664
rect 7564 59356 7616 59362
rect 7564 59298 7616 59304
rect 4988 57928 5040 57934
rect 4988 57870 5040 57876
rect 5540 57928 5592 57934
rect 5540 57870 5592 57876
rect 5552 54534 5580 57870
rect 7576 56642 7604 59298
rect 9600 57882 9628 60658
rect 9600 57854 9720 57882
rect 7564 56636 7616 56642
rect 7564 56578 7616 56584
rect 9692 56438 9720 57854
rect 10428 56506 10456 62630
rect 12084 56574 12112 63854
rect 10784 56568 10836 56574
rect 10784 56510 10836 56516
rect 12072 56568 12124 56574
rect 12072 56510 12124 56516
rect 13728 56568 13780 56574
rect 13728 56510 13780 56516
rect 17960 56568 18012 56574
rect 17960 56510 18012 56516
rect 10416 56500 10468 56506
rect 10416 56442 10468 56448
rect 9680 56432 9732 56438
rect 9680 56374 9732 56380
rect 10796 54670 10824 56510
rect 12440 56500 12492 56506
rect 12440 56442 12492 56448
rect 10784 54664 10836 54670
rect 10784 54606 10836 54612
rect 5540 54528 5592 54534
rect 5540 54470 5592 54476
rect 11704 54528 11756 54534
rect 11704 54470 11756 54476
rect 11716 51134 11744 54470
rect 12452 52766 12480 56442
rect 13636 54664 13688 54670
rect 13636 54606 13688 54612
rect 12440 52760 12492 52766
rect 12440 52702 12492 52708
rect 13648 52494 13676 54606
rect 13740 53038 13768 56510
rect 17972 54126 18000 56510
rect 17960 54120 18012 54126
rect 17960 54062 18012 54068
rect 13728 53032 13780 53038
rect 13728 52974 13780 52980
rect 15200 53032 15252 53038
rect 15200 52974 15252 52980
rect 14556 52760 14608 52766
rect 14556 52702 14608 52708
rect 13636 52488 13688 52494
rect 13636 52430 13688 52436
rect 11704 51128 11756 51134
rect 11704 51070 11756 51076
rect 4068 46844 4120 46850
rect 4068 46786 4120 46792
rect 14568 46306 14596 52702
rect 15212 49706 15240 52974
rect 19248 52420 19300 52426
rect 19248 52362 19300 52368
rect 15292 51060 15344 51066
rect 15292 51002 15344 51008
rect 15200 49700 15252 49706
rect 15200 49642 15252 49648
rect 15304 47326 15332 51002
rect 16856 49700 16908 49706
rect 16856 49642 16908 49648
rect 16868 48210 16896 49642
rect 19260 49609 19288 52362
rect 19246 49600 19302 49609
rect 19246 49535 19302 49544
rect 16856 48204 16908 48210
rect 16856 48146 16908 48152
rect 15292 47320 15344 47326
rect 15292 47262 15344 47268
rect 19248 47320 19300 47326
rect 19248 47262 19300 47268
rect 14556 46300 14608 46306
rect 14556 46242 14608 46248
rect 19260 46238 19288 47262
rect 19996 46374 20024 292538
rect 359464 155372 359516 155378
rect 359464 155314 359516 155320
rect 20904 84244 20956 84250
rect 20956 84192 21404 84194
rect 20904 84186 21404 84192
rect 20916 84166 21404 84186
rect 20076 70440 20128 70446
rect 20076 70382 20128 70388
rect 20088 46510 20116 70382
rect 21376 64874 21404 84166
rect 21284 64846 21404 64874
rect 20904 60036 20956 60042
rect 20904 59978 20956 59984
rect 20916 59945 20944 59978
rect 20902 59936 20958 59945
rect 20902 59871 20958 59880
rect 21284 55298 21312 64846
rect 21454 59936 21510 59945
rect 21454 59871 21510 59880
rect 21284 55270 21404 55298
rect 20628 54120 20680 54126
rect 20628 54062 20680 54068
rect 20640 48226 20668 54062
rect 20640 48198 20760 48226
rect 20076 46504 20128 46510
rect 20076 46446 20128 46452
rect 19984 46368 20036 46374
rect 19984 46310 20036 46316
rect 19248 46232 19300 46238
rect 19248 46174 19300 46180
rect 20732 46102 20760 48198
rect 20812 48204 20864 48210
rect 20812 48146 20864 48152
rect 20824 46170 20852 48146
rect 21376 46442 21404 55270
rect 21364 46436 21416 46442
rect 21364 46378 21416 46384
rect 20812 46164 20864 46170
rect 20812 46106 20864 46112
rect 20720 46096 20772 46102
rect 20720 46038 20772 46044
rect 3976 45484 4028 45490
rect 3976 45426 4028 45432
rect 3884 45416 3936 45422
rect 3884 45358 3936 45364
rect 21468 45354 21496 59871
rect 359476 46617 359504 155314
rect 359556 129056 359608 129062
rect 359556 128998 359608 129004
rect 359462 46608 359518 46617
rect 359462 46543 359518 46552
rect 359568 46306 359596 128998
rect 359556 46300 359608 46306
rect 359556 46242 359608 46248
rect 21456 45348 21508 45354
rect 21456 45290 21508 45296
rect 65524 45280 65576 45286
rect 65524 45222 65576 45228
rect 62028 45212 62080 45218
rect 62028 45154 62080 45160
rect 58440 45144 58492 45150
rect 58440 45086 58492 45092
rect 54944 45076 54996 45082
rect 54944 45018 54996 45024
rect 51356 45008 51408 45014
rect 51356 44950 51408 44956
rect 47860 44940 47912 44946
rect 47860 44882 47912 44888
rect 7656 44872 7708 44878
rect 7656 44814 7708 44820
rect 4068 39364 4120 39370
rect 4068 39306 4120 39312
rect 3424 31748 3476 31754
rect 3424 31690 3476 31696
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2870 3632 2926 3641
rect 2870 3567 2926 3576
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 570 3360 626 3369
rect 570 3295 626 3304
rect 584 480 612 3295
rect 1688 480 1716 3431
rect 2884 480 2912 3567
rect 4080 480 4108 39306
rect 5264 28348 5316 28354
rect 5264 28290 5316 28296
rect 5276 480 5304 28290
rect 6460 3256 6512 3262
rect 6460 3198 6512 3204
rect 6472 480 6500 3198
rect 7668 480 7696 44814
rect 12348 42084 12400 42090
rect 12348 42026 12400 42032
rect 8758 4040 8814 4049
rect 8758 3975 8814 3984
rect 8772 480 8800 3975
rect 9954 3768 10010 3777
rect 9954 3703 10010 3712
rect 9968 480 9996 3703
rect 12360 480 12388 42026
rect 40684 39636 40736 39642
rect 40684 39578 40736 39584
rect 37188 39568 37240 39574
rect 37188 39510 37240 39516
rect 33600 39500 33652 39506
rect 33600 39442 33652 39448
rect 26516 39432 26568 39438
rect 26516 39374 26568 39380
rect 18236 33856 18288 33862
rect 18236 33798 18288 33804
rect 14740 31068 14792 31074
rect 14740 31010 14792 31016
rect 13542 3904 13598 3913
rect 13542 3839 13598 3848
rect 13556 480 13584 3839
rect 14752 480 14780 31010
rect 17038 3224 17094 3233
rect 17038 3159 17094 3168
rect 17052 480 17080 3159
rect 18248 480 18276 33798
rect 23020 33788 23072 33794
rect 23020 33730 23072 33736
rect 19432 28416 19484 28422
rect 19432 28358 19484 28364
rect 19444 480 19472 28358
rect 21824 3596 21876 3602
rect 21824 3538 21876 3544
rect 21836 480 21864 3538
rect 23032 480 23060 33730
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24228 480 24256 3402
rect 26528 480 26556 39374
rect 31300 33924 31352 33930
rect 31300 33866 31352 33872
rect 28908 28552 28960 28558
rect 28908 28494 28960 28500
rect 27712 3528 27764 3534
rect 27712 3470 27764 3476
rect 27724 480 27752 3470
rect 28920 480 28948 28494
rect 30104 3732 30156 3738
rect 30104 3674 30156 3680
rect 30116 480 30144 3674
rect 31312 480 31340 33866
rect 32404 28620 32456 28626
rect 32404 28562 32456 28568
rect 32416 480 32444 28562
rect 33612 480 33640 39442
rect 34796 33992 34848 33998
rect 34796 33934 34848 33940
rect 34808 480 34836 33934
rect 35992 28688 36044 28694
rect 35992 28630 36044 28636
rect 36004 480 36032 28630
rect 37200 480 37228 39510
rect 39580 3868 39632 3874
rect 39580 3810 39632 3816
rect 38384 3800 38436 3806
rect 38384 3742 38436 3748
rect 38396 480 38424 3742
rect 39592 480 39620 3810
rect 40696 480 40724 39578
rect 45468 34128 45520 34134
rect 45468 34070 45520 34076
rect 41880 34060 41932 34066
rect 41880 34002 41932 34008
rect 41892 480 41920 34002
rect 43076 28280 43128 28286
rect 43076 28222 43128 28228
rect 43088 480 43116 28222
rect 44272 3664 44324 3670
rect 44272 3606 44324 3612
rect 44284 480 44312 3606
rect 45480 480 45508 34070
rect 46664 3936 46716 3942
rect 46664 3878 46716 3884
rect 46676 480 46704 3878
rect 47872 480 47900 44882
rect 48964 39704 49016 39710
rect 48964 39646 49016 39652
rect 48976 480 49004 39646
rect 50160 34196 50212 34202
rect 50160 34138 50212 34144
rect 50172 480 50200 34138
rect 51368 480 51396 44950
rect 52552 39772 52604 39778
rect 52552 39714 52604 39720
rect 52564 480 52592 39714
rect 53748 4004 53800 4010
rect 53748 3946 53800 3952
rect 53760 480 53788 3946
rect 54956 480 54984 45018
rect 56048 39840 56100 39846
rect 56048 39782 56100 39788
rect 56060 480 56088 39782
rect 57244 31136 57296 31142
rect 57244 31078 57296 31084
rect 57256 480 57284 31078
rect 58452 480 58480 45086
rect 59636 39908 59688 39914
rect 59636 39850 59688 39856
rect 59648 480 59676 39850
rect 60832 31204 60884 31210
rect 60832 31146 60884 31152
rect 60844 480 60872 31146
rect 62040 480 62068 45154
rect 63224 39976 63276 39982
rect 63224 39918 63276 39924
rect 63236 480 63264 39918
rect 64328 31272 64380 31278
rect 64328 31214 64380 31220
rect 64340 480 64368 31214
rect 65536 480 65564 45222
rect 69112 44804 69164 44810
rect 69112 44746 69164 44752
rect 66720 36576 66772 36582
rect 66720 36518 66772 36524
rect 66732 480 66760 36518
rect 67916 31340 67968 31346
rect 67916 31282 67968 31288
rect 67928 480 67956 31282
rect 69124 480 69152 44746
rect 72608 44736 72660 44742
rect 72608 44678 72660 44684
rect 70308 36644 70360 36650
rect 70308 36586 70360 36592
rect 70320 480 70348 36586
rect 71504 31408 71556 31414
rect 71504 31350 71556 31356
rect 71516 480 71544 31350
rect 72620 480 72648 44678
rect 76196 44668 76248 44674
rect 76196 44610 76248 44616
rect 73804 36712 73856 36718
rect 73804 36654 73856 36660
rect 73816 480 73844 36654
rect 75000 4072 75052 4078
rect 75000 4014 75052 4020
rect 75012 480 75040 4014
rect 76208 480 76236 44610
rect 111616 42764 111668 42770
rect 111616 42706 111668 42712
rect 108120 42696 108172 42702
rect 108120 42638 108172 42644
rect 104532 42628 104584 42634
rect 104532 42570 104584 42576
rect 101036 42560 101088 42566
rect 101036 42502 101088 42508
rect 97448 42492 97500 42498
rect 97448 42434 97500 42440
rect 93952 42424 94004 42430
rect 93952 42366 94004 42372
rect 90364 42356 90416 42362
rect 90364 42298 90416 42304
rect 86868 42288 86920 42294
rect 86868 42230 86920 42236
rect 83280 42220 83332 42226
rect 83280 42162 83332 42168
rect 79692 42152 79744 42158
rect 79692 42094 79744 42100
rect 77392 36780 77444 36786
rect 77392 36722 77444 36728
rect 77404 480 77432 36722
rect 78588 31476 78640 31482
rect 78588 31418 78640 31424
rect 78600 480 78628 31418
rect 79704 480 79732 42094
rect 80888 36848 80940 36854
rect 80888 36790 80940 36796
rect 80900 480 80928 36790
rect 82084 4140 82136 4146
rect 82084 4082 82136 4088
rect 82096 480 82124 4082
rect 83292 480 83320 42162
rect 84476 36916 84528 36922
rect 84476 36858 84528 36864
rect 84488 480 84516 36858
rect 85672 31544 85724 31550
rect 85672 31486 85724 31492
rect 85684 480 85712 31486
rect 86880 480 86908 42230
rect 87972 37052 88024 37058
rect 87972 36994 88024 37000
rect 87984 480 88012 36994
rect 89168 3392 89220 3398
rect 89168 3334 89220 3340
rect 89180 480 89208 3334
rect 90376 480 90404 42298
rect 91560 36984 91612 36990
rect 91560 36926 91612 36932
rect 91572 480 91600 36926
rect 92756 31612 92808 31618
rect 92756 31554 92808 31560
rect 92768 480 92796 31554
rect 93964 480 93992 42366
rect 95148 37120 95200 37126
rect 95148 37062 95200 37068
rect 95160 480 95188 37062
rect 96252 31680 96304 31686
rect 96252 31622 96304 31628
rect 96264 480 96292 31622
rect 97460 480 97488 42434
rect 98644 37188 98696 37194
rect 98644 37130 98696 37136
rect 98656 480 98684 37130
rect 99840 31000 99892 31006
rect 99840 30942 99892 30948
rect 99852 480 99880 30942
rect 101048 480 101076 42502
rect 102232 37256 102284 37262
rect 102232 37198 102284 37204
rect 102244 480 102272 37198
rect 103336 3324 103388 3330
rect 103336 3266 103388 3272
rect 103348 480 103376 3266
rect 104544 480 104572 42570
rect 105728 36508 105780 36514
rect 105728 36450 105780 36456
rect 105740 480 105768 36450
rect 106924 28756 106976 28762
rect 106924 28698 106976 28704
rect 106936 480 106964 28698
rect 108132 480 108160 42638
rect 109316 34264 109368 34270
rect 109316 34206 109368 34212
rect 109328 480 109356 34206
rect 109684 28484 109736 28490
rect 109684 28426 109736 28432
rect 109696 3262 109724 28426
rect 109684 3256 109736 3262
rect 109684 3198 109736 3204
rect 110512 3256 110564 3262
rect 110512 3198 110564 3204
rect 110524 480 110552 3198
rect 111628 480 111656 42706
rect 115204 42016 115256 42022
rect 115204 41958 115256 41964
rect 112812 34332 112864 34338
rect 112812 34274 112864 34280
rect 112824 480 112852 34274
rect 114008 28824 114060 28830
rect 114008 28766 114060 28772
rect 114020 480 114048 28766
rect 115216 480 115244 41958
rect 118792 40044 118844 40050
rect 118792 39986 118844 39992
rect 116400 34400 116452 34406
rect 116400 34342 116452 34348
rect 116412 480 116440 34342
rect 117596 28960 117648 28966
rect 117596 28902 117648 28908
rect 117608 480 117636 28902
rect 118804 480 118832 39986
rect 122288 39296 122340 39302
rect 122288 39238 122340 39244
rect 119896 34468 119948 34474
rect 119896 34410 119948 34416
rect 119908 480 119936 34410
rect 121092 28892 121144 28898
rect 121092 28834 121144 28840
rect 121104 480 121132 28834
rect 122300 480 122328 39238
rect 123484 33720 123536 33726
rect 123484 33662 123536 33668
rect 123496 480 123524 33662
rect 124680 28212 124732 28218
rect 124680 28154 124732 28160
rect 124692 480 124720 28154
rect 360856 3262 360884 305594
rect 361764 304972 361816 304978
rect 361764 304914 361816 304920
rect 361776 304473 361804 304914
rect 361762 304464 361818 304473
rect 361762 304399 361818 304408
rect 361028 304360 361080 304366
rect 361028 304302 361080 304308
rect 360936 304292 360988 304298
rect 360936 304234 360988 304240
rect 360948 3738 360976 304234
rect 360936 3732 360988 3738
rect 360936 3674 360988 3680
rect 361040 3330 361068 304302
rect 362222 302832 362278 302841
rect 362222 302767 362278 302776
rect 361120 300144 361172 300150
rect 361120 300086 361172 300092
rect 361132 3398 361160 300086
rect 361764 293956 361816 293962
rect 361764 293898 361816 293904
rect 361776 293457 361804 293898
rect 361762 293448 361818 293457
rect 361762 293383 361818 293392
rect 361764 282872 361816 282878
rect 361764 282814 361816 282820
rect 361776 282441 361804 282814
rect 361762 282432 361818 282441
rect 361762 282367 361818 282376
rect 361764 271856 361816 271862
rect 361764 271798 361816 271804
rect 361776 271425 361804 271798
rect 361762 271416 361818 271425
rect 361762 271351 361818 271360
rect 361212 268388 361264 268394
rect 361212 268330 361264 268336
rect 361224 3874 361252 268330
rect 361764 260840 361816 260846
rect 361764 260782 361816 260788
rect 361776 260409 361804 260782
rect 361762 260400 361818 260409
rect 361762 260335 361818 260344
rect 361764 249756 361816 249762
rect 361764 249698 361816 249704
rect 361776 249393 361804 249698
rect 361762 249384 361818 249393
rect 361762 249319 361818 249328
rect 361764 238740 361816 238746
rect 361764 238682 361816 238688
rect 361776 238377 361804 238682
rect 361762 238368 361818 238377
rect 361762 238303 361818 238312
rect 361764 227724 361816 227730
rect 361764 227666 361816 227672
rect 361776 227361 361804 227666
rect 361762 227352 361818 227361
rect 361762 227287 361818 227296
rect 361672 216368 361724 216374
rect 361670 216336 361672 216345
rect 361724 216336 361726 216345
rect 361670 216271 361726 216280
rect 361764 205624 361816 205630
rect 361764 205566 361816 205572
rect 361776 205329 361804 205566
rect 361762 205320 361818 205329
rect 361762 205255 361818 205264
rect 361764 194540 361816 194546
rect 361764 194482 361816 194488
rect 361776 194313 361804 194482
rect 361762 194304 361818 194313
rect 361762 194239 361818 194248
rect 361764 183524 361816 183530
rect 361764 183466 361816 183472
rect 361776 183297 361804 183466
rect 361762 183288 361818 183297
rect 361762 183223 361818 183232
rect 361764 172508 361816 172514
rect 361764 172450 361816 172456
rect 361776 172281 361804 172450
rect 361762 172272 361818 172281
rect 361762 172207 361818 172216
rect 361580 163532 361632 163538
rect 361580 163474 361632 163480
rect 361592 155378 361620 163474
rect 361764 161424 361816 161430
rect 361764 161366 361816 161372
rect 361776 161265 361804 161366
rect 361762 161256 361818 161265
rect 361762 161191 361818 161200
rect 361580 155372 361632 155378
rect 361580 155314 361632 155320
rect 361764 150408 361816 150414
rect 361764 150350 361816 150356
rect 361776 150249 361804 150350
rect 361762 150240 361818 150249
rect 361762 150175 361818 150184
rect 361764 139392 361816 139398
rect 361764 139334 361816 139340
rect 361776 139233 361804 139334
rect 361762 139224 361818 139233
rect 361762 139159 361818 139168
rect 361764 128308 361816 128314
rect 361764 128250 361816 128256
rect 361776 128217 361804 128250
rect 361762 128208 361818 128217
rect 361762 128143 361818 128152
rect 361304 118720 361356 118726
rect 361304 118662 361356 118668
rect 361316 46102 361344 118662
rect 361764 117292 361816 117298
rect 361764 117234 361816 117240
rect 361776 117201 361804 117234
rect 361762 117192 361818 117201
rect 361762 117127 361818 117136
rect 361396 111852 361448 111858
rect 361396 111794 361448 111800
rect 361408 46170 361436 111794
rect 361764 106276 361816 106282
rect 361764 106218 361816 106224
rect 361776 106185 361804 106218
rect 361762 106176 361818 106185
rect 361762 106111 361818 106120
rect 361764 95192 361816 95198
rect 361762 95160 361764 95169
rect 361816 95160 361818 95169
rect 361762 95095 361818 95104
rect 361764 84176 361816 84182
rect 361762 84144 361764 84153
rect 361816 84144 361818 84153
rect 361762 84079 361818 84088
rect 361764 73160 361816 73166
rect 361762 73128 361764 73137
rect 361816 73128 361818 73137
rect 361762 73063 361818 73072
rect 361762 62112 361818 62121
rect 361762 62047 361764 62056
rect 361816 62047 361818 62056
rect 361764 62018 361816 62024
rect 361764 51128 361816 51134
rect 361762 51096 361764 51105
rect 361816 51096 361818 51105
rect 361762 51031 361818 51040
rect 361396 46164 361448 46170
rect 361396 46106 361448 46112
rect 361304 46096 361356 46102
rect 361304 46038 361356 46044
rect 362236 4049 362264 302767
rect 363604 300280 363656 300286
rect 363604 300222 363656 300228
rect 362500 297832 362552 297838
rect 362500 297774 362552 297780
rect 362406 297664 362462 297673
rect 362316 297628 362368 297634
rect 362406 297599 362462 297608
rect 362316 297570 362368 297576
rect 362222 4040 362278 4049
rect 362222 3975 362278 3984
rect 361212 3868 361264 3874
rect 361212 3810 361264 3816
rect 362328 3602 362356 297570
rect 362420 39438 362448 297599
rect 362512 39574 362540 297774
rect 362960 124908 363012 124914
rect 362960 124850 363012 124856
rect 362972 122834 363000 124850
rect 362880 122806 363000 122834
rect 362880 118726 362908 122806
rect 362868 118720 362920 118726
rect 362868 118662 362920 118668
rect 362592 117972 362644 117978
rect 362592 117914 362644 117920
rect 362604 46238 362632 117914
rect 362592 46232 362644 46238
rect 362592 46174 362644 46180
rect 362500 39568 362552 39574
rect 362500 39510 362552 39516
rect 362408 39432 362460 39438
rect 362408 39374 362460 39380
rect 363616 3942 363644 300222
rect 363972 297900 364024 297906
rect 363972 297842 364024 297848
rect 363788 297560 363840 297566
rect 363788 297502 363840 297508
rect 363696 291848 363748 291854
rect 363696 291790 363748 291796
rect 363708 33998 363736 291790
rect 363800 39642 363828 297502
rect 363880 297424 363932 297430
rect 363880 297366 363932 297372
rect 363892 39710 363920 297366
rect 363880 39704 363932 39710
rect 363880 39646 363932 39652
rect 363788 39636 363840 39642
rect 363788 39578 363840 39584
rect 363984 39506 364012 297842
rect 364076 216374 364104 333950
rect 365168 305720 365220 305726
rect 365168 305662 365220 305668
rect 364984 301504 365036 301510
rect 364984 301446 365036 301452
rect 364064 216368 364116 216374
rect 364064 216310 364116 216316
rect 364064 116884 364116 116890
rect 364064 116826 364116 116832
rect 364076 111858 364104 116826
rect 364064 111852 364116 111858
rect 364064 111794 364116 111800
rect 363972 39500 364024 39506
rect 363972 39442 364024 39448
rect 363696 33992 363748 33998
rect 363696 33934 363748 33940
rect 364996 4010 365024 301446
rect 365074 297528 365130 297537
rect 365074 297463 365130 297472
rect 364984 4004 365036 4010
rect 364984 3946 365036 3952
rect 363604 3936 363656 3942
rect 363604 3878 363656 3884
rect 362316 3596 362368 3602
rect 362316 3538 362368 3544
rect 361120 3392 361172 3398
rect 361120 3334 361172 3340
rect 361028 3324 361080 3330
rect 361028 3266 361080 3272
rect 360844 3256 360896 3262
rect 365088 3233 365116 297463
rect 365180 39302 365208 305662
rect 367744 302932 367796 302938
rect 367744 302874 367796 302880
rect 366548 297696 366600 297702
rect 366548 297638 366600 297644
rect 365444 297492 365496 297498
rect 365444 297434 365496 297440
rect 365350 297392 365406 297401
rect 365350 297327 365406 297336
rect 365260 286340 365312 286346
rect 365260 286282 365312 286288
rect 365168 39296 365220 39302
rect 365168 39238 365220 39244
rect 365272 28762 365300 286282
rect 365364 39370 365392 297327
rect 365456 40050 365484 297434
rect 366364 291916 366416 291922
rect 366364 291858 366416 291864
rect 365444 40044 365496 40050
rect 365444 39986 365496 39992
rect 365352 39364 365404 39370
rect 365352 39306 365404 39312
rect 365260 28756 365312 28762
rect 365260 28698 365312 28704
rect 366376 3806 366404 291858
rect 366456 286408 366508 286414
rect 366456 286350 366508 286356
rect 366468 28830 366496 286350
rect 366560 39778 366588 297638
rect 366640 294704 366692 294710
rect 366640 294646 366692 294652
rect 366652 39914 366680 294646
rect 366916 118652 366968 118658
rect 366916 118594 366968 118600
rect 366928 116890 366956 118594
rect 366916 116884 366968 116890
rect 366916 116826 366968 116832
rect 366640 39908 366692 39914
rect 366640 39850 366692 39856
rect 366548 39772 366600 39778
rect 366548 39714 366600 39720
rect 366456 28824 366508 28830
rect 366456 28766 366508 28772
rect 367756 4146 367784 302874
rect 367836 301572 367888 301578
rect 367836 301514 367888 301520
rect 367744 4140 367796 4146
rect 367744 4082 367796 4088
rect 367848 4078 367876 301514
rect 367928 300416 367980 300422
rect 367928 300358 367980 300364
rect 367940 42022 367968 300358
rect 368204 300348 368256 300354
rect 368204 300290 368256 300296
rect 368020 300212 368072 300218
rect 368020 300154 368072 300160
rect 368032 42702 368060 300154
rect 368112 297764 368164 297770
rect 368112 297706 368164 297712
rect 368020 42696 368072 42702
rect 368020 42638 368072 42644
rect 367928 42016 367980 42022
rect 367928 41958 367980 41964
rect 368124 39846 368152 297706
rect 368216 42770 368244 300290
rect 369032 166320 369084 166326
rect 369032 166262 369084 166268
rect 369044 163538 369072 166262
rect 369032 163532 369084 163538
rect 369032 163474 369084 163480
rect 368296 126268 368348 126274
rect 368296 126210 368348 126216
rect 368308 117978 368336 126210
rect 368296 117972 368348 117978
rect 368296 117914 368348 117920
rect 368204 42764 368256 42770
rect 368204 42706 368256 42712
rect 368112 39840 368164 39846
rect 368112 39782 368164 39788
rect 369136 28966 369164 386378
rect 370516 379438 370544 601666
rect 371240 582888 371292 582894
rect 371240 582830 371292 582836
rect 371252 578950 371280 582830
rect 371240 578944 371292 578950
rect 371240 578886 371292 578892
rect 371896 380798 371924 623766
rect 374000 578944 374052 578950
rect 374000 578886 374052 578892
rect 374012 575550 374040 578886
rect 374000 575544 374052 575550
rect 374000 575486 374052 575492
rect 374644 386504 374696 386510
rect 374644 386446 374696 386452
rect 373264 385076 373316 385082
rect 373264 385018 373316 385024
rect 371884 380792 371936 380798
rect 371884 380734 371936 380740
rect 370504 379432 370556 379438
rect 370504 379374 370556 379380
rect 371884 339516 371936 339522
rect 371884 339458 371936 339464
rect 371896 315994 371924 339458
rect 371884 315988 371936 315994
rect 371884 315930 371936 315936
rect 370594 305688 370650 305697
rect 370594 305623 370650 305632
rect 369308 295180 369360 295186
rect 369308 295122 369360 295128
rect 369216 292120 369268 292126
rect 369216 292062 369268 292068
rect 369228 34066 369256 292062
rect 369320 36650 369348 295122
rect 369400 294636 369452 294642
rect 369400 294578 369452 294584
rect 369412 39982 369440 294578
rect 370504 286612 370556 286618
rect 370504 286554 370556 286560
rect 369400 39976 369452 39982
rect 369400 39918 369452 39924
rect 369308 36644 369360 36650
rect 369308 36586 369360 36592
rect 369216 34060 369268 34066
rect 369216 34002 369268 34008
rect 369124 28960 369176 28966
rect 369124 28902 369176 28908
rect 370516 20670 370544 286554
rect 370608 42566 370636 305623
rect 371884 303476 371936 303482
rect 371884 303418 371936 303424
rect 370872 300756 370924 300762
rect 370872 300698 370924 300704
rect 370780 300484 370832 300490
rect 370780 300426 370832 300432
rect 370688 294772 370740 294778
rect 370688 294714 370740 294720
rect 370596 42560 370648 42566
rect 370596 42502 370648 42508
rect 370700 36582 370728 294714
rect 370792 42634 370820 300426
rect 370780 42628 370832 42634
rect 370780 42570 370832 42576
rect 370884 42498 370912 300698
rect 370964 300552 371016 300558
rect 370964 300494 371016 300500
rect 370872 42492 370924 42498
rect 370872 42434 370924 42440
rect 370976 42430 371004 300494
rect 371240 122120 371292 122126
rect 371240 122062 371292 122068
rect 371252 118726 371280 122062
rect 371240 118720 371292 118726
rect 371240 118662 371292 118668
rect 370964 42424 371016 42430
rect 370964 42366 371016 42372
rect 370688 36576 370740 36582
rect 370688 36518 370740 36524
rect 370504 20664 370556 20670
rect 370504 20606 370556 20612
rect 371896 6866 371924 303418
rect 372252 294840 372304 294846
rect 372252 294782 372304 294788
rect 372160 294568 372212 294574
rect 371974 294536 372030 294545
rect 372160 294510 372212 294516
rect 371974 294471 372030 294480
rect 371884 6860 371936 6866
rect 371884 6802 371936 6808
rect 367836 4072 367888 4078
rect 367836 4014 367888 4020
rect 371988 3913 372016 294471
rect 372068 286544 372120 286550
rect 372068 286486 372120 286492
rect 372080 28422 372108 286486
rect 372172 36786 372200 294510
rect 372160 36780 372212 36786
rect 372160 36722 372212 36728
rect 372264 36718 372292 294782
rect 372344 289128 372396 289134
rect 372344 289070 372396 289076
rect 372252 36712 372304 36718
rect 372252 36654 372304 36660
rect 372356 34134 372384 289070
rect 372344 34128 372396 34134
rect 372344 34070 372396 34076
rect 373276 28898 373304 385018
rect 373724 302864 373776 302870
rect 373724 302806 373776 302812
rect 373356 300824 373408 300830
rect 373356 300766 373408 300772
rect 373368 42226 373396 300766
rect 373540 300688 373592 300694
rect 373540 300630 373592 300636
rect 373448 300620 373500 300626
rect 373448 300562 373500 300568
rect 373460 42294 373488 300562
rect 373552 42362 373580 300630
rect 373632 294908 373684 294914
rect 373632 294850 373684 294856
rect 373540 42356 373592 42362
rect 373540 42298 373592 42304
rect 373448 42288 373500 42294
rect 373448 42230 373500 42236
rect 373356 42220 373408 42226
rect 373356 42162 373408 42168
rect 373644 36854 373672 294850
rect 373736 45354 373764 302806
rect 373724 45348 373776 45354
rect 373724 45290 373776 45296
rect 373632 36848 373684 36854
rect 373632 36790 373684 36796
rect 373264 28892 373316 28898
rect 373264 28834 373316 28840
rect 372068 28416 372120 28422
rect 372068 28358 372120 28364
rect 374656 28218 374684 386446
rect 374748 382226 374776 645866
rect 374736 382220 374788 382226
rect 374736 382162 374788 382168
rect 376036 382158 376064 656882
rect 378140 575476 378192 575482
rect 378140 575418 378192 575424
rect 378152 569906 378180 575418
rect 378140 569900 378192 569906
rect 378140 569842 378192 569848
rect 378796 383586 378824 667898
rect 400864 634840 400916 634846
rect 400864 634782 400916 634788
rect 380348 569900 380400 569906
rect 380348 569842 380400 569848
rect 380360 563038 380388 569842
rect 380348 563032 380400 563038
rect 380348 562974 380400 562980
rect 382280 563032 382332 563038
rect 382280 562974 382332 562980
rect 382292 559774 382320 562974
rect 382280 559768 382332 559774
rect 382280 559710 382332 559716
rect 385040 559768 385092 559774
rect 385040 559710 385092 559716
rect 385052 555626 385080 559710
rect 385040 555620 385092 555626
rect 385040 555562 385092 555568
rect 387064 555620 387116 555626
rect 387064 555562 387116 555568
rect 387076 553450 387104 555562
rect 387064 553444 387116 553450
rect 387064 553386 387116 553392
rect 389824 553376 389876 553382
rect 389824 553318 389876 553324
rect 389836 541006 389864 553318
rect 389824 541000 389876 541006
rect 389824 540942 389876 540948
rect 392308 540932 392360 540938
rect 392308 540874 392360 540880
rect 392320 536858 392348 540874
rect 392308 536852 392360 536858
rect 392308 536794 392360 536800
rect 394700 536784 394752 536790
rect 394700 536726 394752 536732
rect 394712 529922 394740 536726
rect 394700 529916 394752 529922
rect 394700 529858 394752 529864
rect 396724 529916 396776 529922
rect 396724 529858 396776 529864
rect 396736 511970 396764 529858
rect 396724 511964 396776 511970
rect 396724 511906 396776 511912
rect 381544 491360 381596 491366
rect 381544 491302 381596 491308
rect 378784 383580 378836 383586
rect 378784 383522 378836 383528
rect 376024 382152 376076 382158
rect 376024 382094 376076 382100
rect 381556 372570 381584 491302
rect 396724 469260 396776 469266
rect 396724 469202 396776 469208
rect 382924 386572 382976 386578
rect 382924 386514 382976 386520
rect 381544 372564 381596 372570
rect 381544 372506 381596 372512
rect 380164 307080 380216 307086
rect 380164 307022 380216 307028
rect 378876 306196 378928 306202
rect 378876 306138 378928 306144
rect 378784 305992 378836 305998
rect 378784 305934 378836 305940
rect 378600 303612 378652 303618
rect 378600 303554 378652 303560
rect 375840 303544 375892 303550
rect 375840 303486 375892 303492
rect 374920 295316 374972 295322
rect 374920 295258 374972 295264
rect 374828 295112 374880 295118
rect 374828 295054 374880 295060
rect 374736 295044 374788 295050
rect 374736 294986 374788 294992
rect 374748 36922 374776 294986
rect 374840 37058 374868 295054
rect 374932 37194 374960 295258
rect 375104 292188 375156 292194
rect 375104 292130 375156 292136
rect 375012 289808 375064 289814
rect 375012 289750 375064 289756
rect 374920 37188 374972 37194
rect 374920 37130 374972 37136
rect 374828 37052 374880 37058
rect 374828 36994 374880 37000
rect 374736 36916 374788 36922
rect 374736 36858 374788 36864
rect 375024 34202 375052 289750
rect 375116 37262 375144 292130
rect 375196 161560 375248 161566
rect 375196 161502 375248 161508
rect 375208 73166 375236 161502
rect 375196 73160 375248 73166
rect 375196 73102 375248 73108
rect 375852 46374 375880 303486
rect 376024 303340 376076 303346
rect 376024 303282 376076 303288
rect 375932 302728 375984 302734
rect 375932 302670 375984 302676
rect 375944 46578 375972 302670
rect 375932 46572 375984 46578
rect 375932 46514 375984 46520
rect 375840 46368 375892 46374
rect 375840 46310 375892 46316
rect 376036 42158 376064 303282
rect 376484 303272 376536 303278
rect 376484 303214 376536 303220
rect 376392 303068 376444 303074
rect 376392 303010 376444 303016
rect 376208 300076 376260 300082
rect 376208 300018 376260 300024
rect 376116 289196 376168 289202
rect 376116 289138 376168 289144
rect 376024 42152 376076 42158
rect 376024 42094 376076 42100
rect 375104 37256 375156 37262
rect 375104 37198 375156 37204
rect 375012 34196 375064 34202
rect 375012 34138 375064 34144
rect 376128 31006 376156 289138
rect 376220 42090 376248 300018
rect 376300 294976 376352 294982
rect 376300 294918 376352 294924
rect 376208 42084 376260 42090
rect 376208 42026 376260 42032
rect 376312 37126 376340 294918
rect 376404 44742 376432 303010
rect 376392 44736 376444 44742
rect 376392 44678 376444 44684
rect 376496 44674 376524 303214
rect 376576 303000 376628 303006
rect 376576 302942 376628 302948
rect 376588 44810 376616 302942
rect 376668 302796 376720 302802
rect 376668 302738 376720 302744
rect 376680 46646 376708 302738
rect 377680 292324 377732 292330
rect 377680 292266 377732 292272
rect 377588 289468 377640 289474
rect 377588 289410 377640 289416
rect 377496 289264 377548 289270
rect 377496 289206 377548 289212
rect 377404 286476 377456 286482
rect 377404 286418 377456 286424
rect 376668 46640 376720 46646
rect 376668 46582 376720 46588
rect 376576 44804 376628 44810
rect 376576 44746 376628 44752
rect 376484 44668 376536 44674
rect 376484 44610 376536 44616
rect 376300 37120 376352 37126
rect 376300 37062 376352 37068
rect 376116 31000 376168 31006
rect 376116 30942 376168 30948
rect 377416 28558 377444 286418
rect 377508 31346 377536 289206
rect 377496 31340 377548 31346
rect 377496 31282 377548 31288
rect 377600 31142 377628 289410
rect 377692 34338 377720 292266
rect 377772 291984 377824 291990
rect 377772 291926 377824 291932
rect 377784 36514 377812 291926
rect 378612 46714 378640 303554
rect 378690 302968 378746 302977
rect 378690 302903 378746 302912
rect 378600 46708 378652 46714
rect 378600 46650 378652 46656
rect 378704 45218 378732 302903
rect 378796 45422 378824 305934
rect 378888 46782 378916 306138
rect 379150 303240 379206 303249
rect 379150 303175 379206 303184
rect 379428 303204 379480 303210
rect 379060 292256 379112 292262
rect 379060 292198 379112 292204
rect 378968 289332 379020 289338
rect 378968 289274 379020 289280
rect 378876 46776 378928 46782
rect 378876 46718 378928 46724
rect 378784 45416 378836 45422
rect 378784 45358 378836 45364
rect 378692 45212 378744 45218
rect 378692 45154 378744 45160
rect 377772 36508 377824 36514
rect 377772 36450 377824 36456
rect 377680 34332 377732 34338
rect 377680 34274 377732 34280
rect 378980 31686 379008 289274
rect 379072 34270 379100 292198
rect 379164 45014 379192 303175
rect 379428 303146 379480 303152
rect 379244 303136 379296 303142
rect 379244 303078 379296 303084
rect 379334 303104 379390 303113
rect 379256 45150 379284 303078
rect 379334 303039 379390 303048
rect 379244 45144 379296 45150
rect 379244 45086 379296 45092
rect 379348 45082 379376 303039
rect 379440 45286 379468 303146
rect 379428 45280 379480 45286
rect 379428 45222 379480 45228
rect 379336 45076 379388 45082
rect 379336 45018 379388 45024
rect 379152 45008 379204 45014
rect 379152 44950 379204 44956
rect 379060 34264 379112 34270
rect 379060 34206 379112 34212
rect 378968 31680 379020 31686
rect 378968 31622 379020 31628
rect 377588 31136 377640 31142
rect 377588 31078 377640 31084
rect 380176 28626 380204 307022
rect 382004 306264 382056 306270
rect 382004 306206 382056 306212
rect 382094 306232 382150 306241
rect 381910 306096 381966 306105
rect 381820 306060 381872 306066
rect 381910 306031 381966 306040
rect 381820 306002 381872 306008
rect 381726 305960 381782 305969
rect 381726 305895 381782 305904
rect 381542 305824 381598 305833
rect 381542 305759 381598 305768
rect 381636 305788 381688 305794
rect 381452 295248 381504 295254
rect 381452 295190 381504 295196
rect 380532 292052 380584 292058
rect 380532 291994 380584 292000
rect 380438 291816 380494 291825
rect 380438 291751 380494 291760
rect 380256 289672 380308 289678
rect 380256 289614 380308 289620
rect 380268 31414 380296 289614
rect 380348 289400 380400 289406
rect 380348 289342 380400 289348
rect 380256 31408 380308 31414
rect 380256 31350 380308 31356
rect 380360 31210 380388 289342
rect 380452 33862 380480 291751
rect 380544 34406 380572 291994
rect 381360 278044 381412 278050
rect 381360 277986 381412 277992
rect 381372 45558 381400 277986
rect 381360 45552 381412 45558
rect 381360 45494 381412 45500
rect 381464 36990 381492 295190
rect 381452 36984 381504 36990
rect 381452 36926 381504 36932
rect 380532 34400 380584 34406
rect 380532 34342 380584 34348
rect 380440 33856 380492 33862
rect 380440 33798 380492 33804
rect 380348 31204 380400 31210
rect 380348 31146 380400 31152
rect 380164 28620 380216 28626
rect 380164 28562 380216 28568
rect 377404 28552 377456 28558
rect 377404 28494 377456 28500
rect 374644 28212 374696 28218
rect 374644 28154 374696 28160
rect 371974 3904 372030 3913
rect 371974 3839 372030 3848
rect 366364 3800 366416 3806
rect 366364 3742 366416 3748
rect 381556 3641 381584 305759
rect 381636 305730 381688 305736
rect 381648 45490 381676 305730
rect 381636 45484 381688 45490
rect 381636 45426 381688 45432
rect 381542 3632 381598 3641
rect 381542 3567 381598 3576
rect 381740 3505 381768 305895
rect 381832 46918 381860 306002
rect 381820 46912 381872 46918
rect 381820 46854 381872 46860
rect 381924 44946 381952 306031
rect 382016 46850 382044 306206
rect 382094 306167 382150 306176
rect 382004 46844 382056 46850
rect 382004 46786 382056 46792
rect 381912 44940 381964 44946
rect 381912 44882 381964 44888
rect 382108 44878 382136 306167
rect 382188 289604 382240 289610
rect 382188 289546 382240 289552
rect 382096 44872 382148 44878
rect 382096 44814 382148 44820
rect 382200 31618 382228 289546
rect 382936 33726 382964 386514
rect 396736 371210 396764 469202
rect 399484 447160 399536 447166
rect 399484 447102 399536 447108
rect 396724 371204 396776 371210
rect 396724 371146 396776 371152
rect 399496 369850 399524 447102
rect 400876 380730 400904 634782
rect 403624 557592 403676 557598
rect 403624 557534 403676 557540
rect 400956 511964 401008 511970
rect 400956 511906 401008 511912
rect 400968 495514 400996 511906
rect 400956 495508 401008 495514
rect 400956 495450 401008 495456
rect 402244 495508 402296 495514
rect 402244 495450 402296 495456
rect 402256 462398 402284 495450
rect 402244 462392 402296 462398
rect 402244 462334 402296 462340
rect 400864 380724 400916 380730
rect 400864 380666 400916 380672
rect 403636 376718 403664 557534
rect 406384 535492 406436 535498
rect 406384 535434 406436 535440
rect 405004 462392 405056 462398
rect 405004 462334 405056 462340
rect 405016 454034 405044 462334
rect 405004 454028 405056 454034
rect 405004 453970 405056 453976
rect 403624 376712 403676 376718
rect 403624 376654 403676 376660
rect 406396 375358 406424 535434
rect 407764 524476 407816 524482
rect 407764 524418 407816 524424
rect 406384 375352 406436 375358
rect 406384 375294 406436 375300
rect 407776 375290 407804 524418
rect 410524 513392 410576 513398
rect 410524 513334 410576 513340
rect 408408 454028 408460 454034
rect 408408 453970 408460 453976
rect 408420 448594 408448 453970
rect 408408 448588 408460 448594
rect 408408 448530 408460 448536
rect 410432 448520 410484 448526
rect 410432 448462 410484 448468
rect 410444 445738 410472 448462
rect 410432 445732 410484 445738
rect 410432 445674 410484 445680
rect 407764 375284 407816 375290
rect 407764 375226 407816 375232
rect 410536 373998 410564 513334
rect 411904 502376 411956 502382
rect 411904 502318 411956 502324
rect 410524 373992 410576 373998
rect 410524 373934 410576 373940
rect 411916 373930 411944 502318
rect 413284 445732 413336 445738
rect 413284 445674 413336 445680
rect 413296 433294 413324 445674
rect 413284 433288 413336 433294
rect 413284 433230 413336 433236
rect 411904 373924 411956 373930
rect 411904 373866 411956 373872
rect 409880 369912 409932 369918
rect 409880 369854 409932 369860
rect 399484 369844 399536 369850
rect 399484 369786 399536 369792
rect 409892 365702 409920 369854
rect 409880 365696 409932 365702
rect 409880 365638 409932 365644
rect 407028 350600 407080 350606
rect 407028 350542 407080 350548
rect 402244 347812 402296 347818
rect 402244 347754 402296 347760
rect 402256 337414 402284 347754
rect 402244 337408 402296 337414
rect 402244 337350 402296 337356
rect 399484 335368 399536 335374
rect 399484 335310 399536 335316
rect 385682 306912 385738 306921
rect 385682 306847 385738 306856
rect 383200 306332 383252 306338
rect 383200 306274 383252 306280
rect 383108 304428 383160 304434
rect 383108 304370 383160 304376
rect 383016 297968 383068 297974
rect 383016 297910 383068 297916
rect 382924 33720 382976 33726
rect 382924 33662 382976 33668
rect 382188 31612 382240 31618
rect 382188 31554 382240 31560
rect 383028 3670 383056 297910
rect 383120 28694 383148 304370
rect 383212 33114 383240 306274
rect 384672 306128 384724 306134
rect 384672 306070 384724 306076
rect 384488 305856 384540 305862
rect 384488 305798 384540 305804
rect 384396 305584 384448 305590
rect 384396 305526 384448 305532
rect 384304 292528 384356 292534
rect 384304 292470 384356 292476
rect 383476 292392 383528 292398
rect 383476 292334 383528 292340
rect 383292 289536 383344 289542
rect 383292 289478 383344 289484
rect 383200 33108 383252 33114
rect 383200 33050 383252 33056
rect 383304 31482 383332 289478
rect 383384 289060 383436 289066
rect 383384 289002 383436 289008
rect 383292 31476 383344 31482
rect 383292 31418 383344 31424
rect 383396 31278 383424 289002
rect 383488 34474 383516 292334
rect 384212 159452 384264 159458
rect 384212 159394 384264 159400
rect 384224 84182 384252 159394
rect 384212 84176 384264 84182
rect 384212 84118 384264 84124
rect 383476 34468 383528 34474
rect 383476 34410 383528 34416
rect 383384 31272 383436 31278
rect 383384 31214 383436 31220
rect 383108 28688 383160 28694
rect 383108 28630 383160 28636
rect 383016 3664 383068 3670
rect 383016 3606 383068 3612
rect 384316 3534 384344 292470
rect 384408 46753 384436 305526
rect 384394 46744 384450 46753
rect 384394 46679 384450 46688
rect 384500 46442 384528 305798
rect 384580 305516 384632 305522
rect 384580 305458 384632 305464
rect 384592 46510 384620 305458
rect 384684 46889 384712 306070
rect 384856 305924 384908 305930
rect 384856 305866 384908 305872
rect 384764 289740 384816 289746
rect 384764 289682 384816 289688
rect 384670 46880 384726 46889
rect 384670 46815 384726 46824
rect 384580 46504 384632 46510
rect 384580 46446 384632 46452
rect 384488 46436 384540 46442
rect 384488 46378 384540 46384
rect 384776 31550 384804 289682
rect 384868 47054 384896 305866
rect 384948 119400 385000 119406
rect 384948 119342 385000 119348
rect 384856 47048 384908 47054
rect 384856 46990 384908 46996
rect 384764 31544 384816 31550
rect 384764 31486 384816 31492
rect 384960 28354 384988 119342
rect 384948 28348 385000 28354
rect 384948 28290 385000 28296
rect 384304 3528 384356 3534
rect 381726 3496 381782 3505
rect 384304 3470 384356 3476
rect 385696 3466 385724 306847
rect 385776 304496 385828 304502
rect 385776 304438 385828 304444
rect 385788 3777 385816 304438
rect 386052 292460 386104 292466
rect 386052 292402 386104 292408
rect 385960 291780 386012 291786
rect 385960 291722 386012 291728
rect 385868 288992 385920 288998
rect 385868 288934 385920 288940
rect 385880 31074 385908 288934
rect 385972 33794 386000 291722
rect 386064 33930 386092 292402
rect 399496 249762 399524 335310
rect 402256 334914 402284 337350
rect 407040 335354 407068 350542
rect 413100 336864 413152 336870
rect 413100 336806 413152 336812
rect 409420 336796 409472 336802
rect 409420 336738 409472 336744
rect 406120 335326 407068 335354
rect 406120 334914 406148 335326
rect 402086 334886 402284 334914
rect 405766 334886 406148 334914
rect 409432 334900 409460 336738
rect 413112 334900 413140 336806
rect 413664 336122 413692 703520
rect 418804 700664 418856 700670
rect 418804 700606 418856 700612
rect 416044 685228 416096 685234
rect 416044 685170 416096 685176
rect 414664 458244 414716 458250
rect 414664 458186 414716 458192
rect 414676 371142 414704 458186
rect 414756 433288 414808 433294
rect 414756 433230 414808 433236
rect 414768 420986 414796 433230
rect 414756 420980 414808 420986
rect 414756 420922 414808 420928
rect 414664 371136 414716 371142
rect 414664 371078 414716 371084
rect 416056 336190 416084 685170
rect 416136 436144 416188 436150
rect 416136 436086 416188 436092
rect 416148 369782 416176 436086
rect 417424 425128 417476 425134
rect 417424 425070 417476 425076
rect 416136 369776 416188 369782
rect 416136 369718 416188 369724
rect 417436 368490 417464 425070
rect 417424 368484 417476 368490
rect 417424 368426 417476 368432
rect 416780 336932 416832 336938
rect 416780 336874 416832 336880
rect 416044 336184 416096 336190
rect 416044 336126 416096 336132
rect 413652 336116 413704 336122
rect 413652 336058 413704 336064
rect 416792 334900 416820 336874
rect 418816 336258 418844 700606
rect 418896 700460 418948 700466
rect 418896 700402 418948 700408
rect 418908 336394 418936 700402
rect 418988 685296 419040 685302
rect 418988 685238 419040 685244
rect 418896 336388 418948 336394
rect 418896 336330 418948 336336
rect 419000 336326 419028 685238
rect 420276 684684 420328 684690
rect 420276 684626 420328 684632
rect 420184 684616 420236 684622
rect 420184 684558 420236 684564
rect 419080 546508 419132 546514
rect 419080 546450 419132 546456
rect 419092 376650 419120 546450
rect 419172 480276 419224 480282
rect 419172 480218 419224 480224
rect 419080 376644 419132 376650
rect 419080 376586 419132 376592
rect 419184 372502 419212 480218
rect 419172 372496 419224 372502
rect 419172 372438 419224 372444
rect 418988 336320 419040 336326
rect 418988 336262 419040 336268
rect 418804 336252 418856 336258
rect 418804 336194 418856 336200
rect 420196 334830 420224 684558
rect 420288 334898 420316 684626
rect 420828 683664 420880 683670
rect 420828 683606 420880 683612
rect 420368 683596 420420 683602
rect 420368 683538 420420 683544
rect 420276 334892 420328 334898
rect 420276 334834 420328 334840
rect 420184 334824 420236 334830
rect 420380 334778 420408 683538
rect 420644 683528 420696 683534
rect 420644 683470 420696 683476
rect 420552 683392 420604 683398
rect 420552 683334 420604 683340
rect 420564 335034 420592 683334
rect 420552 335028 420604 335034
rect 420552 334970 420604 334976
rect 420184 334766 420236 334772
rect 420288 334762 420408 334778
rect 420276 334756 420408 334762
rect 420328 334750 420408 334756
rect 420276 334698 420328 334704
rect 420656 334694 420684 683470
rect 420736 683460 420788 683466
rect 420736 683402 420788 683408
rect 420644 334688 420696 334694
rect 420644 334630 420696 334636
rect 420748 334626 420776 683402
rect 420840 334966 420868 683606
rect 422484 447432 422536 447438
rect 422484 447374 422536 447380
rect 422496 444924 422524 447374
rect 427452 447228 427504 447234
rect 427452 447170 427504 447176
rect 427464 444924 427492 447170
rect 429856 445058 429884 703520
rect 445024 700868 445076 700874
rect 445024 700810 445076 700816
rect 444104 700732 444156 700738
rect 444104 700674 444156 700680
rect 437388 447364 437440 447370
rect 437388 447306 437440 447312
rect 432420 447296 432472 447302
rect 432420 447238 432472 447244
rect 429844 445052 429896 445058
rect 429844 444994 429896 445000
rect 432432 444924 432460 447238
rect 437400 444924 437428 447306
rect 442382 444378 442672 444394
rect 442382 444372 442684 444378
rect 442382 444366 442632 444372
rect 442632 444314 442684 444320
rect 420920 420912 420972 420918
rect 420920 420854 420972 420860
rect 420932 417586 420960 420854
rect 421484 417722 421512 420036
rect 421472 417716 421524 417722
rect 421472 417658 421524 417664
rect 420920 417580 420972 417586
rect 420920 417522 420972 417528
rect 422128 417518 422156 420036
rect 422786 420022 423168 420050
rect 423430 420022 423536 420050
rect 422116 417512 422168 417518
rect 422116 417454 422168 417460
rect 423140 416362 423168 420022
rect 423128 416356 423180 416362
rect 423128 416298 423180 416304
rect 423508 393990 423536 420022
rect 424060 417450 424088 420036
rect 424704 417790 424732 420036
rect 424692 417784 424744 417790
rect 424692 417726 424744 417732
rect 425348 417586 425376 420036
rect 425992 417654 426020 420036
rect 442816 419552 442868 419558
rect 442816 419494 442868 419500
rect 425980 417648 426032 417654
rect 425980 417590 426032 417596
rect 425060 417580 425112 417586
rect 425060 417522 425112 417528
rect 425336 417580 425388 417586
rect 425336 417522 425388 417528
rect 424048 417444 424100 417450
rect 424048 417386 424100 417392
rect 423588 416356 423640 416362
rect 423588 416298 423640 416304
rect 423496 393984 423548 393990
rect 423496 393926 423548 393932
rect 423600 391270 423628 416298
rect 425072 413982 425100 417522
rect 425060 413976 425112 413982
rect 425060 413918 425112 413924
rect 427084 413976 427136 413982
rect 427084 413918 427136 413924
rect 427096 397458 427124 413918
rect 439504 403028 439556 403034
rect 439504 402970 439556 402976
rect 427084 397452 427136 397458
rect 427084 397394 427136 397400
rect 428464 397452 428516 397458
rect 428464 397394 428516 397400
rect 423588 391264 423640 391270
rect 423588 391206 423640 391212
rect 428476 387802 428504 397394
rect 428464 387796 428516 387802
rect 428464 387738 428516 387744
rect 431224 387796 431276 387802
rect 431224 387738 431276 387744
rect 431236 369714 431264 387738
rect 431224 369708 431276 369714
rect 431224 369650 431276 369656
rect 432880 369708 432932 369714
rect 432880 369650 432932 369656
rect 432696 363044 432748 363050
rect 432696 362986 432748 362992
rect 432604 361616 432656 361622
rect 432604 361558 432656 361564
rect 431224 339584 431276 339590
rect 431224 339526 431276 339532
rect 427818 336832 427874 336841
rect 427818 336767 427874 336776
rect 420828 334960 420880 334966
rect 420828 334902 420880 334908
rect 427832 334900 427860 336767
rect 420736 334620 420788 334626
rect 420736 334562 420788 334568
rect 420458 334384 420514 334393
rect 420458 334319 420514 334328
rect 424138 334384 424194 334393
rect 424138 334319 424194 334328
rect 431236 304978 431264 339526
rect 431868 328500 431920 328506
rect 431868 328442 431920 328448
rect 431224 304972 431276 304978
rect 431224 304914 431276 304920
rect 420184 262880 420236 262886
rect 420184 262822 420236 262828
rect 420196 256766 420224 262822
rect 414664 256760 414716 256766
rect 414664 256702 414716 256708
rect 420184 256760 420236 256766
rect 420184 256702 420236 256708
rect 399484 249756 399536 249762
rect 399484 249698 399536 249704
rect 414676 203454 414704 256702
rect 429844 253224 429896 253230
rect 429844 253166 429896 253172
rect 429856 241466 429884 253166
rect 427084 241460 427136 241466
rect 427084 241402 427136 241408
rect 429844 241460 429896 241466
rect 429844 241402 429896 241408
rect 427096 229770 427124 241402
rect 421564 229764 421616 229770
rect 421564 229706 421616 229712
rect 427084 229764 427136 229770
rect 427084 229706 427136 229712
rect 410524 203448 410576 203454
rect 410524 203390 410576 203396
rect 414664 203448 414716 203454
rect 414664 203390 414716 203396
rect 407028 186992 407080 186998
rect 407028 186934 407080 186940
rect 407040 184210 407068 186934
rect 395344 184204 395396 184210
rect 395344 184146 395396 184152
rect 407028 184204 407080 184210
rect 407028 184146 407080 184152
rect 395356 174622 395384 184146
rect 389824 174616 389876 174622
rect 389824 174558 389876 174564
rect 395344 174616 395396 174622
rect 395344 174558 395396 174564
rect 389836 166326 389864 174558
rect 389824 166320 389876 166326
rect 389824 166262 389876 166268
rect 408500 164212 408552 164218
rect 408500 164154 408552 164160
rect 386144 160200 386196 160206
rect 386144 160142 386196 160148
rect 386156 62082 386184 160142
rect 408512 159866 408540 164154
rect 409512 160132 409564 160138
rect 409512 160074 409564 160080
rect 401600 159860 401652 159866
rect 401600 159802 401652 159808
rect 408500 159860 408552 159866
rect 408500 159802 408552 159808
rect 386236 159384 386288 159390
rect 386236 159326 386288 159332
rect 386248 95198 386276 159326
rect 400864 156664 400916 156670
rect 400864 156606 400916 156612
rect 396724 156188 396776 156194
rect 396724 156130 396776 156136
rect 395160 150476 395212 150482
rect 395160 150418 395212 150424
rect 395172 147694 395200 150418
rect 391204 147688 391256 147694
rect 391204 147630 391256 147636
rect 395160 147688 395212 147694
rect 395160 147630 395212 147636
rect 391216 137358 391244 147630
rect 389456 137352 389508 137358
rect 389456 137294 389508 137300
rect 391204 137352 391256 137358
rect 391204 137294 391256 137300
rect 388444 137284 388496 137290
rect 388444 137226 388496 137232
rect 387800 135244 387852 135250
rect 387800 135186 387852 135192
rect 387064 129804 387116 129810
rect 387064 129746 387116 129752
rect 387076 122126 387104 129746
rect 387812 128466 387840 135186
rect 388456 129062 388484 137226
rect 389468 135250 389496 137294
rect 396736 136678 396764 156130
rect 396908 153196 396960 153202
rect 396908 153138 396960 153144
rect 396920 150482 396948 153138
rect 396908 150476 396960 150482
rect 396908 150418 396960 150424
rect 400876 145178 400904 156606
rect 401612 153270 401640 159802
rect 409420 159792 409472 159798
rect 409420 159734 409472 159740
rect 409144 159724 409196 159730
rect 409144 159666 409196 159672
rect 406108 159520 406160 159526
rect 406108 159462 406160 159468
rect 406120 157554 406148 159462
rect 404268 157548 404320 157554
rect 404268 157490 404320 157496
rect 406108 157548 406160 157554
rect 406108 157490 406160 157496
rect 404280 156194 404308 157490
rect 404268 156188 404320 156194
rect 404268 156130 404320 156136
rect 401600 153264 401652 153270
rect 401600 153206 401652 153212
rect 407120 147688 407172 147694
rect 407120 147630 407172 147636
rect 407132 145178 407160 147630
rect 396816 145172 396868 145178
rect 396816 145114 396868 145120
rect 400864 145172 400916 145178
rect 400864 145114 400916 145120
rect 404820 145172 404872 145178
rect 404820 145114 404872 145120
rect 407120 145172 407172 145178
rect 407120 145114 407172 145120
rect 396828 137290 396856 145114
rect 404832 142186 404860 145114
rect 401600 142180 401652 142186
rect 401600 142122 401652 142128
rect 404820 142180 404872 142186
rect 404820 142122 404872 142128
rect 396816 137284 396868 137290
rect 396816 137226 396868 137232
rect 401612 136762 401640 142122
rect 401520 136734 401640 136762
rect 394700 136672 394752 136678
rect 394700 136614 394752 136620
rect 396724 136672 396776 136678
rect 396724 136614 396776 136620
rect 391204 135924 391256 135930
rect 391204 135866 391256 135872
rect 389456 135244 389508 135250
rect 389456 135186 389508 135192
rect 391216 129878 391244 135866
rect 394712 132530 394740 136614
rect 401520 135930 401548 136734
rect 401508 135924 401560 135930
rect 401508 135866 401560 135872
rect 394700 132524 394752 132530
rect 394700 132466 394752 132472
rect 391940 132456 391992 132462
rect 391940 132398 391992 132404
rect 389180 129872 389232 129878
rect 389180 129814 389232 129820
rect 391204 129872 391256 129878
rect 391204 129814 391256 129820
rect 388444 129056 388496 129062
rect 388444 128998 388496 129004
rect 387720 128438 387840 128466
rect 387720 126274 387748 128438
rect 387708 126268 387760 126274
rect 387708 126210 387760 126216
rect 389192 125610 389220 129814
rect 391952 129810 391980 132398
rect 391940 129804 391992 129810
rect 391940 129746 391992 129752
rect 389100 125582 389220 125610
rect 389100 124914 389128 125582
rect 389088 124908 389140 124914
rect 389088 124850 389140 124856
rect 387064 122120 387116 122126
rect 387064 122062 387116 122068
rect 389824 106956 389876 106962
rect 389824 106898 389876 106904
rect 389836 104938 389864 106898
rect 409156 106282 409184 159666
rect 409236 159656 409288 159662
rect 409236 159598 409288 159604
rect 409248 128314 409276 159598
rect 409328 159588 409380 159594
rect 409328 159530 409380 159536
rect 409340 139398 409368 159530
rect 409432 147694 409460 159734
rect 409524 150414 409552 160074
rect 410536 156670 410564 203390
rect 421576 193186 421604 229706
rect 418528 193180 418580 193186
rect 418528 193122 418580 193128
rect 421564 193180 421616 193186
rect 421564 193122 421616 193128
rect 418540 186998 418568 193122
rect 431224 190528 431276 190534
rect 431224 190470 431276 190476
rect 418528 186992 418580 186998
rect 418528 186934 418580 186940
rect 431236 175982 431264 190470
rect 419540 175976 419592 175982
rect 419540 175918 419592 175924
rect 431224 175976 431276 175982
rect 431224 175918 431276 175924
rect 419552 173942 419580 175918
rect 414664 173936 414716 173942
rect 414664 173878 414716 173884
rect 419540 173936 419592 173942
rect 419540 173878 419592 173884
rect 414676 169794 414704 173878
rect 414664 169788 414716 169794
rect 414664 169730 414716 169736
rect 411260 169720 411312 169726
rect 411260 169662 411312 169668
rect 411272 164286 411300 169662
rect 429844 168360 429896 168366
rect 429844 168302 429896 168308
rect 411260 164280 411312 164286
rect 411260 164222 411312 164228
rect 421838 162752 421894 162761
rect 421838 162687 421894 162696
rect 425886 162752 425942 162761
rect 425886 162687 425942 162696
rect 428646 162752 428702 162761
rect 428646 162687 428702 162696
rect 418712 162240 418764 162246
rect 418712 162182 418764 162188
rect 415124 162172 415176 162178
rect 415124 162114 415176 162120
rect 412088 161492 412140 161498
rect 412088 161434 412140 161440
rect 412100 159882 412128 161434
rect 415136 160206 415164 162114
rect 418724 161566 418752 162182
rect 418712 161560 418764 161566
rect 418712 161502 418764 161508
rect 415124 160200 415176 160206
rect 411792 159854 412128 159882
rect 415090 160148 415124 160154
rect 415090 160142 415176 160148
rect 415090 160126 415164 160142
rect 415090 159868 415118 160126
rect 418724 159882 418752 161502
rect 421852 160342 421880 162687
rect 425900 160478 425928 162687
rect 425336 160472 425388 160478
rect 425336 160414 425388 160420
rect 425888 160472 425940 160478
rect 425888 160414 425940 160420
rect 421840 160336 421892 160342
rect 421840 160278 421892 160284
rect 418416 159854 418752 159882
rect 421380 159452 421432 159458
rect 421380 159394 421432 159400
rect 421392 159338 421420 159394
rect 421852 159338 421880 160278
rect 425348 159882 425376 160414
rect 428660 160410 428688 162687
rect 428648 160404 428700 160410
rect 428648 160346 428700 160352
rect 427820 160200 427872 160206
rect 427820 160142 427872 160148
rect 425040 159854 425376 159882
rect 425164 159390 425192 159854
rect 427832 159798 427860 160142
rect 427820 159792 427872 159798
rect 428660 159746 428688 160346
rect 429856 160206 429884 168302
rect 431880 161566 431908 328442
rect 432616 325553 432644 361558
rect 432708 329225 432736 362986
rect 432788 362976 432840 362982
rect 432788 362918 432840 362924
rect 432800 332897 432828 362918
rect 432892 349110 432920 369650
rect 439516 367062 439544 402970
rect 442724 387796 442776 387802
rect 442724 387738 442776 387744
rect 441528 387116 441580 387122
rect 441528 387058 441580 387064
rect 439504 367056 439556 367062
rect 439504 366998 439556 367004
rect 439780 360324 439832 360330
rect 439780 360266 439832 360272
rect 436928 360256 436980 360262
rect 436928 360198 436980 360204
rect 435456 358828 435508 358834
rect 435456 358770 435508 358776
rect 432880 349104 432932 349110
rect 432880 349046 432932 349052
rect 435364 338156 435416 338162
rect 435364 338098 435416 338104
rect 432786 332888 432842 332897
rect 432786 332823 432842 332832
rect 432788 330268 432840 330274
rect 432788 330210 432840 330216
rect 432694 329216 432750 329225
rect 432694 329151 432750 329160
rect 432602 325544 432658 325553
rect 432602 325479 432658 325488
rect 432604 322992 432656 322998
rect 432604 322934 432656 322940
rect 432052 318300 432104 318306
rect 432052 318242 432104 318248
rect 432064 310865 432092 318242
rect 432616 314537 432644 322934
rect 432800 318209 432828 330210
rect 432880 324964 432932 324970
rect 432880 324906 432932 324912
rect 432892 321881 432920 324906
rect 432878 321872 432934 321881
rect 432878 321807 432934 321816
rect 432786 318200 432842 318209
rect 432786 318135 432842 318144
rect 432602 314528 432658 314537
rect 432602 314463 432658 314472
rect 432696 313948 432748 313954
rect 432696 313890 432748 313896
rect 432050 310856 432106 310865
rect 432050 310791 432106 310800
rect 432708 307193 432736 313890
rect 432694 307184 432750 307193
rect 432694 307119 432750 307128
rect 435376 293962 435404 338098
rect 435468 318306 435496 358770
rect 436836 338224 436888 338230
rect 436836 338166 436888 338172
rect 436744 332648 436796 332654
rect 436744 332590 436796 332596
rect 436008 328568 436060 328574
rect 436008 328510 436060 328516
rect 435456 318300 435508 318306
rect 435456 318242 435508 318248
rect 435364 293956 435416 293962
rect 435364 293898 435416 293904
rect 433340 202836 433392 202842
rect 433340 202778 433392 202784
rect 433352 196058 433380 202778
rect 433260 196030 433380 196058
rect 433260 190534 433288 196030
rect 433248 190528 433300 190534
rect 433248 190470 433300 190476
rect 432236 169788 432288 169794
rect 432236 169730 432288 169736
rect 432248 168434 432276 169730
rect 432236 168428 432288 168434
rect 432236 168370 432288 168376
rect 431868 161560 431920 161566
rect 431868 161502 431920 161508
rect 429844 160200 429896 160206
rect 429844 160142 429896 160148
rect 431880 159882 431908 161502
rect 436020 160274 436048 328510
rect 436756 194546 436784 332590
rect 436848 282878 436876 338166
rect 436940 322998 436968 360198
rect 437020 349104 437072 349110
rect 437020 349046 437072 349052
rect 437032 325038 437060 349046
rect 439688 335096 439740 335102
rect 439688 335038 439740 335044
rect 439596 332716 439648 332722
rect 439596 332658 439648 332664
rect 439504 330472 439556 330478
rect 439504 330414 439556 330420
rect 437020 325032 437072 325038
rect 437020 324974 437072 324980
rect 439320 325032 439372 325038
rect 439320 324974 439372 324980
rect 436928 322992 436980 322998
rect 436928 322934 436980 322940
rect 439332 322250 439360 324974
rect 439320 322244 439372 322250
rect 439320 322186 439372 322192
rect 436836 282872 436888 282878
rect 436836 282814 436888 282820
rect 437756 258732 437808 258738
rect 437756 258674 437808 258680
rect 437768 253230 437796 258674
rect 437756 253224 437808 253230
rect 437756 253166 437808 253172
rect 437480 208412 437532 208418
rect 437480 208354 437532 208360
rect 437492 202910 437520 208354
rect 437480 202904 437532 202910
rect 437480 202846 437532 202852
rect 436744 194540 436796 194546
rect 436744 194482 436796 194488
rect 436744 175228 436796 175234
rect 436744 175170 436796 175176
rect 436756 169794 436784 175170
rect 436744 169788 436796 169794
rect 436744 169730 436796 169736
rect 439516 163674 439544 330414
rect 439608 205630 439636 332658
rect 439700 271862 439728 335038
rect 439792 330274 439820 360266
rect 440884 337000 440936 337006
rect 440884 336942 440936 336948
rect 439872 335028 439924 335034
rect 439872 334970 439924 334976
rect 439780 330268 439832 330274
rect 439780 330210 439832 330216
rect 439884 322386 439912 334970
rect 439872 322380 439924 322386
rect 439872 322322 439924 322328
rect 439688 271856 439740 271862
rect 439688 271798 439740 271804
rect 440896 260846 440924 336942
rect 440976 336388 441028 336394
rect 440976 336330 441028 336336
rect 440988 319394 441016 336330
rect 441252 336320 441304 336326
rect 441252 336262 441304 336268
rect 441160 336252 441212 336258
rect 441160 336194 441212 336200
rect 441068 336184 441120 336190
rect 441068 336126 441120 336132
rect 441080 320686 441108 336126
rect 441172 320958 441200 336194
rect 441160 320952 441212 320958
rect 441160 320894 441212 320900
rect 441068 320680 441120 320686
rect 441068 320622 441120 320628
rect 441264 320550 441292 336262
rect 441252 320544 441304 320550
rect 441252 320486 441304 320492
rect 441540 320482 441568 387058
rect 442264 361684 442316 361690
rect 442264 361626 442316 361632
rect 442276 324970 442304 361626
rect 442356 334960 442408 334966
rect 442356 334902 442408 334908
rect 442264 324964 442316 324970
rect 442264 324906 442316 324912
rect 442368 322318 442396 334902
rect 442448 334892 442500 334898
rect 442448 334834 442500 334840
rect 442356 322312 442408 322318
rect 442356 322254 442408 322260
rect 442460 322182 442488 334834
rect 442448 322176 442500 322182
rect 442448 322118 442500 322124
rect 441528 320476 441580 320482
rect 441528 320418 441580 320424
rect 442736 320074 442764 387738
rect 442724 320068 442776 320074
rect 442724 320010 442776 320016
rect 440976 319388 441028 319394
rect 440976 319330 441028 319336
rect 442828 319190 442856 419494
rect 443644 414044 443696 414050
rect 443644 413986 443696 413992
rect 443656 368422 443684 413986
rect 443736 392012 443788 392018
rect 443736 391954 443788 391960
rect 443644 368416 443696 368422
rect 443644 368358 443696 368364
rect 443748 366994 443776 391954
rect 443828 380928 443880 380934
rect 443828 380870 443880 380876
rect 443736 366988 443788 366994
rect 443736 366930 443788 366936
rect 443840 365634 443868 380870
rect 443828 365628 443880 365634
rect 443828 365570 443880 365576
rect 443828 358896 443880 358902
rect 443828 358838 443880 358844
rect 443736 335708 443788 335714
rect 443736 335650 443788 335656
rect 443644 334076 443696 334082
rect 443644 334018 443696 334024
rect 442908 330404 442960 330410
rect 442908 330346 442960 330352
rect 442816 319184 442868 319190
rect 442816 319126 442868 319132
rect 440884 260840 440936 260846
rect 440884 260782 440936 260788
rect 442264 237448 442316 237454
rect 442264 237390 442316 237396
rect 440884 226636 440936 226642
rect 440884 226578 440936 226584
rect 440896 213926 440924 226578
rect 439688 213920 439740 213926
rect 439688 213862 439740 213868
rect 440884 213920 440936 213926
rect 440884 213862 440936 213868
rect 439700 208418 439728 213862
rect 439688 208412 439740 208418
rect 439688 208354 439740 208360
rect 439596 205624 439648 205630
rect 439596 205566 439648 205572
rect 442276 204270 442304 237390
rect 442448 230036 442500 230042
rect 442448 229978 442500 229984
rect 442460 226642 442488 229978
rect 442448 226636 442500 226642
rect 442448 226578 442500 226584
rect 440884 204264 440936 204270
rect 440884 204206 440936 204212
rect 442264 204264 442316 204270
rect 442264 204206 442316 204212
rect 440896 191826 440924 204206
rect 439596 191820 439648 191826
rect 439596 191762 439648 191768
rect 440884 191820 440936 191826
rect 440884 191762 440936 191768
rect 439608 175302 439636 191762
rect 439596 175296 439648 175302
rect 439596 175238 439648 175244
rect 440240 165980 440292 165986
rect 440240 165922 440292 165928
rect 438584 163668 438636 163674
rect 438584 163610 438636 163616
rect 439504 163668 439556 163674
rect 439504 163610 439556 163616
rect 437572 162308 437624 162314
rect 437572 162250 437624 162256
rect 435272 160268 435324 160274
rect 435272 160210 435324 160216
rect 436008 160268 436060 160274
rect 436008 160210 436060 160216
rect 435284 159882 435312 160210
rect 431664 159854 431908 159882
rect 434824 159854 435312 159882
rect 427820 159734 427872 159740
rect 428016 159730 428688 159746
rect 428004 159724 428688 159730
rect 428056 159718 428688 159724
rect 428004 159666 428056 159672
rect 434824 159662 434852 159854
rect 434812 159656 434864 159662
rect 434812 159598 434864 159604
rect 437584 159526 437612 162250
rect 438596 160206 438624 163610
rect 440252 162314 440280 165922
rect 440240 162308 440292 162314
rect 440240 162250 440292 162256
rect 438584 160200 438636 160206
rect 438584 160142 438636 160148
rect 438596 159610 438624 160142
rect 442920 160138 442948 330346
rect 443184 241188 443236 241194
rect 443184 241130 443236 241136
rect 443196 237454 443224 241130
rect 443184 237448 443236 237454
rect 443184 237390 443236 237396
rect 443656 227730 443684 334018
rect 443748 238746 443776 335650
rect 443840 313954 443868 358838
rect 444116 320822 444144 700674
rect 444288 422952 444340 422958
rect 444288 422894 444340 422900
rect 444196 341012 444248 341018
rect 444196 340954 444248 340960
rect 444208 336054 444236 340954
rect 444196 336048 444248 336054
rect 444196 335990 444248 335996
rect 444104 320816 444156 320822
rect 444104 320758 444156 320764
rect 444300 320006 444328 422894
rect 444932 334824 444984 334830
rect 444932 334766 444984 334772
rect 444944 321230 444972 334766
rect 445036 322522 445064 700810
rect 446496 700800 446548 700806
rect 446496 700742 446548 700748
rect 446404 700596 446456 700602
rect 446404 700538 446456 700544
rect 445116 687948 445168 687954
rect 445116 687890 445168 687896
rect 445024 322516 445076 322522
rect 445024 322458 445076 322464
rect 444932 321224 444984 321230
rect 444932 321166 444984 321172
rect 444288 320000 444340 320006
rect 444288 319942 444340 319948
rect 445128 319734 445156 687890
rect 445208 686520 445260 686526
rect 445208 686462 445260 686468
rect 445220 320113 445248 686462
rect 445300 685160 445352 685166
rect 445300 685102 445352 685108
rect 445206 320104 445262 320113
rect 445206 320039 445262 320048
rect 445116 319728 445168 319734
rect 445116 319670 445168 319676
rect 445312 319258 445340 685102
rect 445574 683360 445630 683369
rect 445484 683324 445536 683330
rect 445574 683295 445630 683304
rect 445484 683266 445536 683272
rect 445392 683256 445444 683262
rect 445392 683198 445444 683204
rect 445404 319530 445432 683198
rect 445496 319598 445524 683266
rect 445588 322794 445616 683295
rect 446312 682712 446364 682718
rect 446312 682654 446364 682660
rect 445668 447228 445720 447234
rect 445668 447170 445720 447176
rect 445680 353326 445708 447170
rect 446220 444372 446272 444378
rect 446220 444314 446272 444320
rect 445668 353320 445720 353326
rect 445668 353262 445720 353268
rect 446232 353122 446260 444314
rect 446220 353116 446272 353122
rect 446220 353058 446272 353064
rect 445668 334756 445720 334762
rect 445668 334698 445720 334704
rect 445576 322788 445628 322794
rect 445576 322730 445628 322736
rect 445484 319592 445536 319598
rect 445484 319534 445536 319540
rect 445392 319524 445444 319530
rect 445392 319466 445444 319472
rect 445680 319326 445708 334698
rect 446324 327486 446352 682654
rect 446312 327480 446364 327486
rect 446312 327422 446364 327428
rect 446416 320890 446444 700538
rect 446508 321434 446536 700742
rect 446588 700528 446640 700534
rect 446588 700470 446640 700476
rect 446600 322454 446628 700470
rect 447876 700460 447928 700466
rect 447876 700402 447928 700408
rect 446680 700324 446732 700330
rect 446680 700266 446732 700272
rect 446692 322833 446720 700266
rect 446864 684548 446916 684554
rect 446864 684490 446916 684496
rect 446770 683224 446826 683233
rect 446770 683159 446826 683168
rect 446678 322824 446734 322833
rect 446678 322759 446734 322768
rect 446588 322448 446640 322454
rect 446588 322390 446640 322396
rect 446496 321428 446548 321434
rect 446496 321370 446548 321376
rect 446404 320884 446456 320890
rect 446404 320826 446456 320832
rect 446784 319841 446812 683159
rect 446876 320618 446904 684490
rect 447048 683188 447100 683194
rect 447048 683130 447100 683136
rect 446954 682816 447010 682825
rect 446954 682751 447010 682760
rect 446864 320612 446916 320618
rect 446864 320554 446916 320560
rect 446770 319832 446826 319841
rect 446770 319767 446826 319776
rect 445668 319320 445720 319326
rect 445668 319262 445720 319268
rect 445300 319252 445352 319258
rect 445300 319194 445352 319200
rect 446968 319122 446996 682751
rect 447060 321094 447088 683130
rect 447784 669996 447836 670002
rect 447784 669938 447836 669944
rect 447324 447976 447376 447982
rect 447324 447918 447376 447924
rect 447232 447908 447284 447914
rect 447232 447850 447284 447856
rect 447140 447840 447192 447846
rect 447140 447782 447192 447788
rect 447152 447370 447180 447782
rect 447140 447364 447192 447370
rect 447140 447306 447192 447312
rect 447244 447302 447272 447850
rect 447336 447438 447364 447918
rect 447692 447840 447744 447846
rect 447692 447782 447744 447788
rect 447324 447432 447376 447438
rect 447324 447374 447376 447380
rect 447232 447296 447284 447302
rect 447232 447238 447284 447244
rect 447140 445052 447192 445058
rect 447140 444994 447192 445000
rect 447152 387802 447180 444994
rect 447140 387796 447192 387802
rect 447140 387738 447192 387744
rect 447416 387320 447468 387326
rect 447416 387262 447468 387268
rect 447140 383648 447192 383654
rect 447138 383616 447140 383625
rect 447192 383616 447194 383625
rect 447138 383551 447194 383560
rect 447232 383580 447284 383586
rect 447232 383522 447284 383528
rect 447244 382945 447272 383522
rect 447230 382936 447286 382945
rect 447230 382871 447286 382880
rect 447138 382256 447194 382265
rect 447138 382191 447194 382200
rect 447232 382220 447284 382226
rect 447152 382158 447180 382191
rect 447232 382162 447284 382168
rect 447140 382152 447192 382158
rect 447140 382094 447192 382100
rect 447244 381585 447272 382162
rect 447230 381576 447286 381585
rect 447230 381511 447286 381520
rect 447230 380896 447286 380905
rect 447230 380831 447286 380840
rect 447140 380792 447192 380798
rect 447140 380734 447192 380740
rect 447152 380225 447180 380734
rect 447244 380730 447272 380831
rect 447232 380724 447284 380730
rect 447232 380666 447284 380672
rect 447138 380216 447194 380225
rect 447138 380151 447194 380160
rect 447324 379500 447376 379506
rect 447324 379442 447376 379448
rect 447140 379432 447192 379438
rect 447140 379374 447192 379380
rect 447152 378865 447180 379374
rect 447138 378856 447194 378865
rect 447138 378791 447194 378800
rect 447336 378185 447364 379442
rect 447322 378176 447378 378185
rect 447232 378140 447284 378146
rect 447322 378111 447378 378120
rect 447232 378082 447284 378088
rect 447140 378072 447192 378078
rect 447140 378014 447192 378020
rect 447152 377505 447180 378014
rect 447138 377496 447194 377505
rect 447138 377431 447194 377440
rect 447244 376825 447272 378082
rect 447230 376816 447286 376825
rect 447230 376751 447286 376760
rect 447140 376712 447192 376718
rect 447140 376654 447192 376660
rect 447152 376145 447180 376654
rect 447232 376644 447284 376650
rect 447232 376586 447284 376592
rect 447138 376136 447194 376145
rect 447138 376071 447194 376080
rect 447244 375465 447272 376586
rect 447230 375456 447286 375465
rect 447230 375391 447286 375400
rect 447140 375352 447192 375358
rect 447140 375294 447192 375300
rect 447152 374785 447180 375294
rect 447232 375284 447284 375290
rect 447232 375226 447284 375232
rect 447138 374776 447194 374785
rect 447138 374711 447194 374720
rect 447244 374105 447272 375226
rect 447230 374096 447286 374105
rect 447230 374031 447286 374040
rect 447140 373992 447192 373998
rect 447140 373934 447192 373940
rect 447152 373425 447180 373934
rect 447232 373924 447284 373930
rect 447232 373866 447284 373872
rect 447138 373416 447194 373425
rect 447138 373351 447194 373360
rect 447244 372745 447272 373866
rect 447230 372736 447286 372745
rect 447230 372671 447286 372680
rect 447140 372564 447192 372570
rect 447140 372506 447192 372512
rect 447152 372065 447180 372506
rect 447232 372496 447284 372502
rect 447232 372438 447284 372444
rect 447138 372056 447194 372065
rect 447138 371991 447194 372000
rect 447244 371385 447272 372438
rect 447230 371376 447286 371385
rect 447230 371311 447286 371320
rect 447140 371204 447192 371210
rect 447140 371146 447192 371152
rect 447152 370705 447180 371146
rect 447232 371136 447284 371142
rect 447232 371078 447284 371084
rect 447138 370696 447194 370705
rect 447138 370631 447194 370640
rect 447244 370025 447272 371078
rect 447230 370016 447286 370025
rect 447230 369951 447286 369960
rect 447140 369844 447192 369850
rect 447140 369786 447192 369792
rect 447152 369345 447180 369786
rect 447232 369776 447284 369782
rect 447232 369718 447284 369724
rect 447138 369336 447194 369345
rect 447138 369271 447194 369280
rect 447244 368665 447272 369718
rect 447230 368656 447286 368665
rect 447230 368591 447286 368600
rect 447140 368484 447192 368490
rect 447140 368426 447192 368432
rect 447152 367985 447180 368426
rect 447232 368416 447284 368422
rect 447232 368358 447284 368364
rect 447138 367976 447194 367985
rect 447138 367911 447194 367920
rect 447244 367305 447272 368358
rect 447230 367296 447286 367305
rect 447230 367231 447286 367240
rect 447140 367056 447192 367062
rect 447140 366998 447192 367004
rect 447152 366625 447180 366998
rect 447232 366988 447284 366994
rect 447232 366930 447284 366936
rect 447138 366616 447194 366625
rect 447138 366551 447194 366560
rect 447244 365945 447272 366930
rect 447230 365936 447286 365945
rect 447230 365871 447286 365880
rect 447140 365696 447192 365702
rect 447140 365638 447192 365644
rect 447152 364585 447180 365638
rect 447232 365628 447284 365634
rect 447232 365570 447284 365576
rect 447244 365265 447272 365570
rect 447230 365256 447286 365265
rect 447230 365191 447286 365200
rect 447138 364576 447194 364585
rect 447138 364511 447194 364520
rect 447230 363896 447286 363905
rect 447230 363831 447286 363840
rect 447138 363216 447194 363225
rect 447138 363151 447194 363160
rect 447152 363050 447180 363151
rect 447140 363044 447192 363050
rect 447140 362986 447192 362992
rect 447244 362982 447272 363831
rect 447232 362976 447284 362982
rect 447232 362918 447284 362924
rect 447138 362536 447194 362545
rect 447138 362471 447194 362480
rect 447152 361622 447180 362471
rect 447230 361856 447286 361865
rect 447230 361791 447286 361800
rect 447244 361690 447272 361791
rect 447232 361684 447284 361690
rect 447232 361626 447284 361632
rect 447140 361616 447192 361622
rect 447140 361558 447192 361564
rect 447230 361176 447286 361185
rect 447230 361111 447286 361120
rect 447138 360496 447194 360505
rect 447138 360431 447194 360440
rect 447152 360262 447180 360431
rect 447244 360330 447272 361111
rect 447232 360324 447284 360330
rect 447232 360266 447284 360272
rect 447140 360256 447192 360262
rect 447140 360198 447192 360204
rect 447138 359816 447194 359825
rect 447138 359751 447194 359760
rect 447152 358834 447180 359751
rect 447230 359136 447286 359145
rect 447230 359071 447286 359080
rect 447244 358902 447272 359071
rect 447232 358896 447284 358902
rect 447232 358838 447284 358844
rect 447140 358828 447192 358834
rect 447140 358770 447192 358776
rect 447428 354385 447456 387262
rect 447600 387252 447652 387258
rect 447600 387194 447652 387200
rect 447508 380860 447560 380866
rect 447508 380802 447560 380808
rect 447520 379545 447548 380802
rect 447506 379536 447562 379545
rect 447506 379471 447562 379480
rect 447414 354376 447470 354385
rect 447414 354311 447470 354320
rect 447612 353705 447640 387194
rect 447598 353696 447654 353705
rect 447598 353631 447654 353640
rect 447322 351656 447378 351665
rect 447322 351591 447378 351600
rect 447138 350976 447194 350985
rect 447138 350911 447194 350920
rect 447152 350606 447180 350911
rect 447140 350600 447192 350606
rect 447140 350542 447192 350548
rect 447140 347744 447192 347750
rect 447140 347686 447192 347692
rect 447152 347585 447180 347686
rect 447138 347576 447194 347585
rect 447138 347511 447194 347520
rect 447138 342136 447194 342145
rect 447138 342071 447194 342080
rect 447152 340950 447180 342071
rect 447230 341456 447286 341465
rect 447230 341391 447286 341400
rect 447244 341018 447272 341391
rect 447232 341012 447284 341018
rect 447232 340954 447284 340960
rect 447140 340944 447192 340950
rect 447140 340886 447192 340892
rect 447230 340776 447286 340785
rect 447230 340711 447286 340720
rect 447138 340096 447194 340105
rect 447138 340031 447194 340040
rect 447152 339590 447180 340031
rect 447140 339584 447192 339590
rect 447140 339526 447192 339532
rect 447244 339522 447272 340711
rect 447232 339516 447284 339522
rect 447232 339458 447284 339464
rect 447230 339416 447286 339425
rect 447230 339351 447286 339360
rect 447138 338736 447194 338745
rect 447138 338671 447194 338680
rect 447152 338230 447180 338671
rect 447140 338224 447192 338230
rect 447140 338166 447192 338172
rect 447244 338162 447272 339351
rect 447232 338156 447284 338162
rect 447232 338098 447284 338104
rect 447138 337376 447194 337385
rect 447138 337311 447194 337320
rect 447152 337006 447180 337311
rect 447140 337000 447192 337006
rect 447140 336942 447192 336948
rect 447138 336696 447194 336705
rect 447138 336631 447194 336640
rect 447152 335374 447180 336631
rect 447230 336016 447286 336025
rect 447230 335951 447286 335960
rect 447244 335714 447272 335951
rect 447232 335708 447284 335714
rect 447232 335650 447284 335656
rect 447140 335368 447192 335374
rect 447140 335310 447192 335316
rect 447230 335336 447286 335345
rect 447230 335271 447286 335280
rect 447138 334656 447194 334665
rect 447138 334591 447194 334600
rect 447152 334014 447180 334591
rect 447244 334082 447272 335271
rect 447232 334076 447284 334082
rect 447232 334018 447284 334024
rect 447140 334008 447192 334014
rect 447140 333950 447192 333956
rect 447230 333976 447286 333985
rect 447230 333911 447286 333920
rect 447138 333296 447194 333305
rect 447138 333231 447194 333240
rect 447152 332654 447180 333231
rect 447244 332722 447272 333911
rect 447232 332716 447284 332722
rect 447232 332658 447284 332664
rect 447140 332648 447192 332654
rect 447140 332590 447192 332596
rect 447230 330576 447286 330585
rect 447140 330540 447192 330546
rect 447230 330511 447286 330520
rect 447140 330482 447192 330488
rect 447048 321088 447100 321094
rect 447048 321030 447100 321036
rect 446956 319116 447008 319122
rect 446956 319058 447008 319064
rect 443828 313948 443880 313954
rect 443828 313890 443880 313896
rect 447152 249762 447180 330482
rect 447244 330410 447272 330511
rect 447232 330404 447284 330410
rect 447232 330346 447284 330352
rect 447140 249756 447192 249762
rect 447140 249698 447192 249704
rect 447152 248946 447180 249698
rect 446404 248940 446456 248946
rect 446404 248882 446456 248888
rect 447140 248940 447192 248946
rect 447140 248882 447192 248888
rect 445760 247036 445812 247042
rect 445760 246978 445812 246984
rect 445668 245608 445720 245614
rect 445668 245550 445720 245556
rect 445680 241194 445708 245550
rect 445668 241188 445720 241194
rect 445668 241130 445720 241136
rect 445772 239834 445800 246978
rect 445208 239828 445260 239834
rect 445208 239770 445260 239776
rect 445760 239828 445812 239834
rect 445760 239770 445812 239776
rect 443736 238740 443788 238746
rect 443736 238682 443788 238688
rect 445220 237454 445248 239770
rect 443920 237448 443972 237454
rect 443920 237390 443972 237396
rect 445208 237448 445260 237454
rect 445208 237390 445260 237396
rect 443932 230042 443960 237390
rect 443920 230036 443972 230042
rect 443920 229978 443972 229984
rect 443644 227724 443696 227730
rect 443644 227666 443696 227672
rect 444012 169788 444064 169794
rect 444012 169730 444064 169736
rect 444024 165986 444052 169730
rect 444012 165980 444064 165986
rect 444012 165922 444064 165928
rect 446416 163674 446444 248882
rect 447232 247716 447284 247722
rect 447232 247658 447284 247664
rect 447244 245682 447272 247658
rect 447232 245676 447284 245682
rect 447232 245618 447284 245624
rect 447336 199442 447364 351591
rect 447506 338056 447562 338065
rect 447506 337991 447562 338000
rect 447520 335102 447548 337991
rect 447508 335096 447560 335102
rect 447508 335038 447560 335044
rect 447704 330585 447732 447782
rect 447796 387122 447824 669938
rect 447888 419558 447916 700402
rect 449164 700392 449216 700398
rect 449164 700334 449216 700340
rect 447968 700324 448020 700330
rect 447968 700266 448020 700272
rect 447980 422958 448008 700266
rect 448980 461100 449032 461106
rect 448980 461042 449032 461048
rect 448428 447976 448480 447982
rect 448428 447918 448480 447924
rect 448060 447908 448112 447914
rect 448060 447850 448112 447856
rect 447968 422952 448020 422958
rect 447968 422894 448020 422900
rect 447876 419552 447928 419558
rect 447876 419494 447928 419500
rect 447876 388544 447928 388550
rect 447876 388486 447928 388492
rect 447784 387116 447836 387122
rect 447784 387058 447836 387064
rect 447888 355065 447916 388486
rect 447968 385688 448020 385694
rect 447968 385630 448020 385636
rect 447874 355056 447930 355065
rect 447874 354991 447930 355000
rect 447876 353320 447928 353326
rect 447876 353262 447928 353268
rect 447784 353116 447836 353122
rect 447784 353058 447836 353064
rect 447796 331265 447824 353058
rect 447888 344865 447916 353262
rect 447980 352345 448008 385630
rect 447966 352336 448022 352345
rect 447966 352271 448022 352280
rect 447966 345536 448022 345545
rect 447966 345471 448022 345480
rect 447874 344856 447930 344865
rect 447874 344791 447930 344800
rect 447876 337408 447928 337414
rect 447876 337350 447928 337356
rect 447782 331256 447838 331265
rect 447782 331191 447838 331200
rect 447690 330576 447746 330585
rect 447888 330546 447916 337350
rect 447690 330511 447746 330520
rect 447876 330540 447928 330546
rect 447876 330482 447928 330488
rect 447416 330472 447468 330478
rect 447416 330414 447468 330420
rect 447428 329905 447456 330414
rect 447414 329896 447470 329905
rect 447414 329831 447470 329840
rect 447508 321156 447560 321162
rect 447508 321098 447560 321104
rect 447520 320618 447548 321098
rect 447508 320612 447560 320618
rect 447508 320554 447560 320560
rect 447980 309806 448008 345471
rect 448072 330478 448100 447850
rect 448336 388476 448388 388482
rect 448336 388418 448388 388424
rect 448152 386028 448204 386034
rect 448152 385970 448204 385976
rect 448164 353025 448192 385970
rect 448244 385416 448296 385422
rect 448244 385358 448296 385364
rect 448150 353016 448206 353025
rect 448150 352951 448206 352960
rect 448256 348945 448284 385358
rect 448348 349625 448376 388418
rect 448440 386646 448468 447918
rect 448428 386640 448480 386646
rect 448428 386582 448480 386588
rect 448334 349616 448390 349625
rect 448334 349551 448390 349560
rect 448242 348936 448298 348945
rect 448242 348871 448298 348880
rect 448440 343505 448468 386582
rect 448992 346905 449020 461042
rect 449070 387016 449126 387025
rect 449070 386951 449126 386960
rect 449084 357105 449112 386951
rect 449070 357096 449126 357105
rect 449070 357031 449126 357040
rect 448978 346896 449034 346905
rect 448978 346831 449034 346840
rect 448426 343496 448482 343505
rect 448426 343431 448482 343440
rect 448440 337414 448468 343431
rect 448428 337408 448480 337414
rect 448428 337350 448480 337356
rect 448150 332616 448206 332625
rect 448150 332551 448206 332560
rect 448060 330472 448112 330478
rect 448060 330414 448112 330420
rect 447968 309800 448020 309806
rect 447968 309742 448020 309748
rect 447784 201340 447836 201346
rect 447784 201282 447836 201288
rect 447324 199436 447376 199442
rect 447324 199378 447376 199384
rect 447232 183524 447284 183530
rect 447232 183466 447284 183472
rect 447244 182850 447272 183466
rect 447232 182844 447284 182850
rect 447232 182786 447284 182792
rect 447232 172508 447284 172514
rect 447232 172450 447284 172456
rect 447244 171834 447272 172450
rect 447232 171828 447284 171834
rect 447232 171770 447284 171776
rect 447796 169794 447824 201282
rect 448164 182850 448192 332551
rect 448334 331936 448390 331945
rect 448334 331871 448390 331880
rect 448152 182844 448204 182850
rect 448152 182786 448204 182792
rect 448348 171834 448376 331871
rect 448426 331256 448482 331265
rect 448426 331191 448482 331200
rect 448336 171828 448388 171834
rect 448336 171770 448388 171776
rect 448440 171134 448468 331191
rect 449176 321366 449204 700334
rect 449256 690668 449308 690674
rect 449256 690610 449308 690616
rect 449164 321360 449216 321366
rect 449164 321302 449216 321308
rect 449268 319870 449296 690610
rect 462332 670002 462360 703520
rect 478524 700466 478552 703520
rect 478512 700460 478564 700466
rect 478512 700402 478564 700408
rect 494808 700330 494836 703520
rect 494796 700324 494848 700330
rect 494796 700266 494848 700272
rect 527192 699825 527220 703520
rect 543476 700369 543504 703520
rect 543462 700360 543518 700369
rect 543462 700295 543518 700304
rect 559668 699825 559696 703520
rect 527178 699816 527234 699825
rect 527178 699751 527234 699760
rect 559654 699816 559710 699825
rect 559654 699751 559710 699760
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 576124 696992 576176 696998
rect 576124 696934 576176 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 462320 669996 462372 670002
rect 462320 669938 462372 669944
rect 457810 667992 457866 668001
rect 457810 667927 457866 667936
rect 457718 652896 457774 652905
rect 457718 652831 457774 652840
rect 457626 650176 457682 650185
rect 457626 650111 457682 650120
rect 457534 645960 457590 645969
rect 457534 645895 457590 645904
rect 457442 643240 457498 643249
rect 457442 643175 457498 643184
rect 457350 640384 457406 640393
rect 457350 640319 457406 640328
rect 457258 637936 457314 637945
rect 457258 637871 457314 637880
rect 457272 599622 457300 637871
rect 457364 599690 457392 640319
rect 457352 599684 457404 599690
rect 457352 599626 457404 599632
rect 457260 599616 457312 599622
rect 457260 599558 457312 599564
rect 457456 598806 457484 643175
rect 457444 598800 457496 598806
rect 457444 598742 457496 598748
rect 457548 597582 457576 645895
rect 457536 597576 457588 597582
rect 457536 597518 457588 597524
rect 457640 596970 457668 650111
rect 457628 596964 457680 596970
rect 457628 596906 457680 596912
rect 450544 596828 450596 596834
rect 450544 596770 450596 596776
rect 449808 518220 449860 518226
rect 449808 518162 449860 518168
rect 449820 503509 449848 518162
rect 450360 517540 450412 517546
rect 450360 517482 450412 517488
rect 449992 516792 450044 516798
rect 449992 516734 450044 516740
rect 450004 507657 450032 516734
rect 450372 510241 450400 517482
rect 450450 516896 450506 516905
rect 450450 516831 450506 516840
rect 450464 514729 450492 516831
rect 450450 514720 450506 514729
rect 450450 514655 450506 514664
rect 450556 512417 450584 596770
rect 457732 595474 457760 652831
rect 457824 600234 457852 667927
rect 458086 662552 458142 662561
rect 458086 662487 458142 662496
rect 457994 659968 458050 659977
rect 457994 659903 458050 659912
rect 457902 657520 457958 657529
rect 457902 657455 457958 657464
rect 457812 600228 457864 600234
rect 457812 600170 457864 600176
rect 457720 595468 457772 595474
rect 457720 595410 457772 595416
rect 457916 551342 457944 657455
rect 457904 551336 457956 551342
rect 457904 551278 457956 551284
rect 458008 523734 458036 659903
rect 457996 523728 458048 523734
rect 457996 523670 458048 523676
rect 458100 518294 458128 662487
rect 571984 643136 572036 643142
rect 571984 643078 572036 643084
rect 458822 635488 458878 635497
rect 458822 635423 458878 635432
rect 458730 611416 458786 611425
rect 458730 611351 458786 611360
rect 458640 604036 458692 604042
rect 458640 603978 458692 603984
rect 458652 596902 458680 603978
rect 458744 599826 458772 611351
rect 458732 599820 458784 599826
rect 458732 599762 458784 599768
rect 458640 596896 458692 596902
rect 458640 596838 458692 596844
rect 458088 518288 458140 518294
rect 458088 518230 458140 518236
rect 458836 518129 458864 635423
rect 459006 633448 459062 633457
rect 459006 633383 459062 633392
rect 458914 623928 458970 623937
rect 458914 623863 458970 623872
rect 458928 604042 458956 623863
rect 458916 604036 458968 604042
rect 458916 603978 458968 603984
rect 459020 603922 459048 633383
rect 459098 630728 459154 630737
rect 459098 630663 459154 630672
rect 458928 603894 459048 603922
rect 458928 599593 458956 603894
rect 459008 603764 459060 603770
rect 459008 603706 459060 603712
rect 459020 599758 459048 603706
rect 459008 599752 459060 599758
rect 459008 599694 459060 599700
rect 458914 599584 458970 599593
rect 458914 599519 458970 599528
rect 459112 589937 459140 630663
rect 459190 628144 459246 628153
rect 459190 628079 459246 628088
rect 459098 589928 459154 589937
rect 459098 589863 459154 589872
rect 459204 587178 459232 628079
rect 459282 625832 459338 625841
rect 459282 625767 459338 625776
rect 459192 587172 459244 587178
rect 459192 587114 459244 587120
rect 459296 584458 459324 625767
rect 459374 621072 459430 621081
rect 459374 621007 459430 621016
rect 459284 584452 459336 584458
rect 459284 584394 459336 584400
rect 459388 519586 459416 621007
rect 460202 618352 460258 618361
rect 460202 618287 460258 618296
rect 459466 616040 459522 616049
rect 459466 615975 459522 615984
rect 459480 603770 459508 615975
rect 460110 613864 460166 613873
rect 460110 613799 460166 613808
rect 460018 608696 460074 608705
rect 460018 608631 460074 608640
rect 459926 606384 459982 606393
rect 459926 606319 459982 606328
rect 459468 603764 459520 603770
rect 459468 603706 459520 603712
rect 459466 603664 459522 603673
rect 459466 603599 459522 603608
rect 459480 598466 459508 603599
rect 459836 602132 459888 602138
rect 459836 602074 459888 602080
rect 459468 598460 459520 598466
rect 459468 598402 459520 598408
rect 459848 597038 459876 602074
rect 459836 597032 459888 597038
rect 459836 596974 459888 596980
rect 459940 594114 459968 606319
rect 459928 594108 459980 594114
rect 459928 594050 459980 594056
rect 460032 592686 460060 608631
rect 460124 602138 460152 613799
rect 460112 602132 460164 602138
rect 460112 602074 460164 602080
rect 460110 602032 460166 602041
rect 460110 601967 460166 601976
rect 460124 600302 460152 601967
rect 460112 600296 460164 600302
rect 460112 600238 460164 600244
rect 460216 598262 460244 618287
rect 570604 616888 570656 616894
rect 570604 616830 570656 616836
rect 462320 600296 462372 600302
rect 462320 600238 462372 600244
rect 461584 600228 461636 600234
rect 461584 600170 461636 600176
rect 460204 598256 460256 598262
rect 460204 598198 460256 598204
rect 460020 592680 460072 592686
rect 460020 592622 460072 592628
rect 459376 519580 459428 519586
rect 459376 519522 459428 519528
rect 458822 518120 458878 518129
rect 458822 518055 458878 518064
rect 450636 516860 450688 516866
rect 450636 516802 450688 516808
rect 450542 512408 450598 512417
rect 450542 512343 450598 512352
rect 450358 510232 450414 510241
rect 450358 510167 450414 510176
rect 450372 509234 450400 510167
rect 450372 509206 450492 509234
rect 449990 507648 450046 507657
rect 449990 507583 450046 507592
rect 449806 503500 449862 503509
rect 449806 503435 449862 503444
rect 449624 457496 449676 457502
rect 449624 457438 449676 457444
rect 449532 454708 449584 454714
rect 449532 454650 449584 454656
rect 449440 387116 449492 387122
rect 449440 387058 449492 387064
rect 449348 385144 449400 385150
rect 449348 385086 449400 385092
rect 449360 348265 449388 385086
rect 449346 348256 449402 348265
rect 449346 348191 449402 348200
rect 449346 344176 449402 344185
rect 449346 344111 449402 344120
rect 449256 319864 449308 319870
rect 449256 319806 449308 319812
rect 448520 262948 448572 262954
rect 448520 262890 448572 262896
rect 448532 258738 448560 262890
rect 448520 258732 448572 258738
rect 448520 258674 448572 258680
rect 449164 258120 449216 258126
rect 449164 258062 449216 258068
rect 449176 247110 449204 258062
rect 449164 247104 449216 247110
rect 449164 247046 449216 247052
rect 449164 243568 449216 243574
rect 449164 243510 449216 243516
rect 449176 201346 449204 243510
rect 449164 201340 449216 201346
rect 449164 201282 449216 201288
rect 448348 171106 448468 171134
rect 447784 169788 447836 169794
rect 447784 169730 447836 169736
rect 445208 163668 445260 163674
rect 445208 163610 445260 163616
rect 446404 163668 446456 163674
rect 446404 163610 446456 163616
rect 445220 161634 445248 163610
rect 445208 161628 445260 161634
rect 445208 161570 445260 161576
rect 441574 160132 441626 160138
rect 441574 160074 441626 160080
rect 442908 160132 442960 160138
rect 442908 160074 442960 160080
rect 441586 159868 441614 160074
rect 445220 159882 445248 161570
rect 448348 161430 448376 171106
rect 449360 164218 449388 344111
rect 449452 342825 449480 387058
rect 449544 356425 449572 454650
rect 449636 357785 449664 457438
rect 449716 454776 449768 454782
rect 449716 454718 449768 454724
rect 449622 357776 449678 357785
rect 449622 357711 449678 357720
rect 449530 356416 449586 356425
rect 449530 356351 449586 356360
rect 449728 355745 449756 454718
rect 449808 387184 449860 387190
rect 449808 387126 449860 387132
rect 449820 358465 449848 387126
rect 449806 358456 449862 358465
rect 449806 358391 449862 358400
rect 449714 355736 449770 355745
rect 449714 355671 449770 355680
rect 449806 350296 449862 350305
rect 449806 350231 449862 350240
rect 449438 342816 449494 342825
rect 449438 342751 449494 342760
rect 449440 336116 449492 336122
rect 449440 336058 449492 336064
rect 449452 319802 449480 336058
rect 449532 334688 449584 334694
rect 449532 334630 449584 334636
rect 449440 319796 449492 319802
rect 449440 319738 449492 319744
rect 449544 319666 449572 334630
rect 449624 334620 449676 334626
rect 449624 334562 449676 334568
rect 449636 319938 449664 334562
rect 449716 327480 449768 327486
rect 449716 327422 449768 327428
rect 449728 320618 449756 327422
rect 449716 320612 449768 320618
rect 449716 320554 449768 320560
rect 449624 319932 449676 319938
rect 449624 319874 449676 319880
rect 449532 319660 449584 319666
rect 449532 319602 449584 319608
rect 449820 263566 449848 350231
rect 450004 334121 450032 507583
rect 450082 505472 450138 505481
rect 450082 505407 450138 505416
rect 450096 338026 450124 505407
rect 450174 503296 450230 503305
rect 450174 503231 450230 503240
rect 450084 338020 450136 338026
rect 450084 337962 450136 337968
rect 450188 336870 450216 503231
rect 450360 338020 450412 338026
rect 450360 337962 450412 337968
rect 450266 337784 450322 337793
rect 450266 337719 450322 337728
rect 450176 336864 450228 336870
rect 450280 336841 450308 337719
rect 450372 336938 450400 337962
rect 450360 336932 450412 336938
rect 450360 336874 450412 336880
rect 450176 336806 450228 336812
rect 450266 336832 450322 336841
rect 449990 334112 450046 334121
rect 449990 334047 450046 334056
rect 449898 328944 449954 328953
rect 449898 328879 449954 328888
rect 449912 328574 449940 328879
rect 449900 328568 449952 328574
rect 449900 328510 449952 328516
rect 450004 326641 450032 334047
rect 450084 330540 450136 330546
rect 450084 330482 450136 330488
rect 449990 326632 450046 326641
rect 449990 326567 450046 326576
rect 450096 324601 450124 330482
rect 450188 325281 450216 336806
rect 450266 336767 450322 336776
rect 450280 328001 450308 336767
rect 450266 327992 450322 328001
rect 450266 327927 450322 327936
rect 450372 325694 450400 336874
rect 450464 335354 450492 509206
rect 450556 462398 450584 512343
rect 450648 505481 450676 516802
rect 450634 505472 450690 505481
rect 450634 505407 450690 505416
rect 450648 500126 450754 500154
rect 451936 500126 452226 500154
rect 450544 462392 450596 462398
rect 450544 462334 450596 462340
rect 450556 337793 450584 462334
rect 450648 402974 450676 500126
rect 450648 402946 450860 402974
rect 450728 387388 450780 387394
rect 450728 387330 450780 387336
rect 450542 337784 450598 337793
rect 450542 337719 450598 337728
rect 450740 336802 450768 387330
rect 450832 385900 450860 402946
rect 451936 385914 451964 500126
rect 453304 497480 453356 497486
rect 453304 497422 453356 497428
rect 452568 496868 452620 496874
rect 452568 496810 452620 496816
rect 452016 455524 452068 455530
rect 452016 455466 452068 455472
rect 451582 385886 451964 385914
rect 452028 385422 452056 455466
rect 452580 385914 452608 496810
rect 453028 389156 453080 389162
rect 453028 389098 453080 389104
rect 452318 385886 452608 385914
rect 453040 385900 453068 389098
rect 453316 386034 453344 497422
rect 453684 496874 453712 500140
rect 454052 500126 455170 500154
rect 453672 496868 453724 496874
rect 453672 496810 453724 496816
rect 453948 496868 454000 496874
rect 453948 496810 454000 496816
rect 453304 386028 453356 386034
rect 453304 385970 453356 385976
rect 453960 385914 453988 496810
rect 454052 389162 454080 500126
rect 455328 497072 455380 497078
rect 455328 497014 455380 497020
rect 455144 496936 455196 496942
rect 455144 496878 455196 496884
rect 454684 455456 454736 455462
rect 454684 455398 454736 455404
rect 454040 389156 454092 389162
rect 454040 389098 454092 389104
rect 454696 387394 454724 455398
rect 455156 393314 455184 496878
rect 455340 393314 455368 497014
rect 456524 497004 456576 497010
rect 456524 496946 456576 496952
rect 456536 393314 456564 496946
rect 456628 496874 456656 500140
rect 457628 497684 457680 497690
rect 457628 497626 457680 497632
rect 457444 497616 457496 497622
rect 457444 497558 457496 497564
rect 456616 496868 456668 496874
rect 456616 496810 456668 496816
rect 454880 393286 455184 393314
rect 455248 393286 455368 393314
rect 456352 393286 456564 393314
rect 454684 387388 454736 387394
rect 454684 387330 454736 387336
rect 454880 385914 454908 393286
rect 453790 385886 453988 385914
rect 454526 385886 454908 385914
rect 455248 385900 455276 393286
rect 456352 385914 456380 393286
rect 456708 389156 456760 389162
rect 456708 389098 456760 389104
rect 455998 385886 456380 385914
rect 456720 385900 456748 389098
rect 457456 387326 457484 497558
rect 457536 428460 457588 428466
rect 457536 428402 457588 428408
rect 457548 389162 457576 428402
rect 457536 389156 457588 389162
rect 457536 389098 457588 389104
rect 457444 387320 457496 387326
rect 457444 387262 457496 387268
rect 457640 386186 457668 497626
rect 458100 496942 458128 500140
rect 458824 497548 458876 497554
rect 458824 497490 458876 497496
rect 458088 496936 458140 496942
rect 458088 496878 458140 496884
rect 458088 430024 458140 430030
rect 458088 429966 458140 429972
rect 458100 393314 458128 429966
rect 457364 386158 457668 386186
rect 457824 393286 458128 393314
rect 457364 385694 457392 386158
rect 457824 385914 457852 393286
rect 458836 388550 458864 497490
rect 459572 497078 459600 500140
rect 459560 497072 459612 497078
rect 459560 497014 459612 497020
rect 461044 497010 461072 500140
rect 461032 497004 461084 497010
rect 461032 496946 461084 496952
rect 458916 460964 458968 460970
rect 458916 460906 458968 460912
rect 458928 447914 458956 460906
rect 459008 454096 459060 454102
rect 459008 454038 459060 454044
rect 459020 447982 459048 454038
rect 459008 447976 459060 447982
rect 459008 447918 459060 447924
rect 458916 447908 458968 447914
rect 458916 447850 458968 447856
rect 459376 429956 459428 429962
rect 459376 429898 459428 429904
rect 459388 393314 459416 429898
rect 459468 429888 459520 429894
rect 459468 429830 459520 429836
rect 459020 393286 459416 393314
rect 458824 388544 458876 388550
rect 458824 388486 458876 388492
rect 459020 386186 459048 393286
rect 458560 386158 459048 386186
rect 458560 385914 458588 386158
rect 459480 386050 459508 429830
rect 460756 395344 460808 395350
rect 460756 395286 460808 395292
rect 459652 389904 459704 389910
rect 459652 389846 459704 389852
rect 459296 386022 459508 386050
rect 459296 385914 459324 386022
rect 457470 385886 457852 385914
rect 458206 385886 458588 385914
rect 458942 385886 459324 385914
rect 459664 385900 459692 389846
rect 460768 385914 460796 395286
rect 461124 388952 461176 388958
rect 461124 388894 461176 388900
rect 460414 385886 460796 385914
rect 461136 385900 461164 388894
rect 461596 388074 461624 600170
rect 461676 598800 461728 598806
rect 461676 598742 461728 598748
rect 461688 388822 461716 598742
rect 461768 520328 461820 520334
rect 461768 520270 461820 520276
rect 461676 388816 461728 388822
rect 461676 388758 461728 388764
rect 461780 388482 461808 520270
rect 461860 497752 461912 497758
rect 461860 497694 461912 497700
rect 461768 388476 461820 388482
rect 461768 388418 461820 388424
rect 461584 388068 461636 388074
rect 461584 388010 461636 388016
rect 461872 387258 461900 497694
rect 462332 402974 462360 600238
rect 463160 600086 463266 600114
rect 469614 600086 469904 600114
rect 475962 600086 476068 600114
rect 462964 597576 463016 597582
rect 462964 597518 463016 597524
rect 462332 402946 462912 402974
rect 462596 388068 462648 388074
rect 462596 388010 462648 388016
rect 462136 387864 462188 387870
rect 462136 387806 462188 387812
rect 461860 387252 461912 387258
rect 461860 387194 461912 387200
rect 462148 385914 462176 387806
rect 461886 385886 462176 385914
rect 462608 385900 462636 388010
rect 462884 385914 462912 402946
rect 462976 388686 463004 597518
rect 463054 517576 463110 517585
rect 463054 517511 463110 517520
rect 462964 388680 463016 388686
rect 462964 388622 463016 388628
rect 463068 388482 463096 517511
rect 463160 501129 463188 600086
rect 465080 599820 465132 599826
rect 465080 599762 465132 599768
rect 463700 598460 463752 598466
rect 463700 598402 463752 598408
rect 463146 501120 463202 501129
rect 463146 501055 463202 501064
rect 463608 392624 463660 392630
rect 463608 392566 463660 392572
rect 463620 388958 463648 392566
rect 463608 388952 463660 388958
rect 463608 388894 463660 388900
rect 463056 388476 463108 388482
rect 463056 388418 463108 388424
rect 463712 385914 463740 598402
rect 464344 596964 464396 596970
rect 464344 596906 464396 596912
rect 463792 594108 463844 594114
rect 463792 594050 463844 594056
rect 463804 402974 463832 594050
rect 463804 402946 464292 402974
rect 464264 385914 464292 402946
rect 464356 388754 464384 596906
rect 464436 518288 464488 518294
rect 464436 518230 464488 518236
rect 464448 402974 464476 518230
rect 464448 402946 464568 402974
rect 464344 388748 464396 388754
rect 464344 388690 464396 388696
rect 464540 388550 464568 402946
rect 464896 389836 464948 389842
rect 464896 389778 464948 389784
rect 464528 388544 464580 388550
rect 464528 388486 464580 388492
rect 464908 387870 464936 389778
rect 465092 389298 465120 599762
rect 466460 599752 466512 599758
rect 466460 599694 466512 599700
rect 465172 592680 465224 592686
rect 465172 592622 465224 592628
rect 465080 389292 465132 389298
rect 465080 389234 465132 389240
rect 464896 387864 464948 387870
rect 464896 387806 464948 387812
rect 465184 385914 465212 592622
rect 465724 523728 465776 523734
rect 465724 523670 465776 523676
rect 465736 388618 465764 523670
rect 466472 389298 466500 599694
rect 467104 599684 467156 599690
rect 467104 599626 467156 599632
rect 466552 597032 466604 597038
rect 466552 596974 466604 596980
rect 465908 389292 465960 389298
rect 465908 389234 465960 389240
rect 466460 389292 466512 389298
rect 466460 389234 466512 389240
rect 465724 388612 465776 388618
rect 465724 388554 465776 388560
rect 465920 385914 465948 389234
rect 466564 385914 466592 596974
rect 467116 389026 467144 599626
rect 468484 599616 468536 599622
rect 468484 599558 468536 599564
rect 467932 598256 467984 598262
rect 467932 598198 467984 598204
rect 467196 551336 467248 551342
rect 467196 551278 467248 551284
rect 467104 389020 467156 389026
rect 467104 388962 467156 388968
rect 467208 388890 467236 551278
rect 467944 402974 467972 598198
rect 467944 402946 468064 402974
rect 467380 389292 467432 389298
rect 467380 389234 467432 389240
rect 467196 388884 467248 388890
rect 467196 388826 467248 388832
rect 467392 385914 467420 389234
rect 468036 385914 468064 402946
rect 468496 389094 468524 599558
rect 469404 596896 469456 596902
rect 469404 596838 469456 596844
rect 468576 595468 468628 595474
rect 468576 595410 468628 595416
rect 468484 389088 468536 389094
rect 468484 389030 468536 389036
rect 468588 388958 468616 595410
rect 469312 519580 469364 519586
rect 469312 519522 469364 519528
rect 468668 461032 468720 461038
rect 468668 460974 468720 460980
rect 468680 447846 468708 460974
rect 468668 447840 468720 447846
rect 468668 447782 468720 447788
rect 469324 393314 469352 519522
rect 469416 402974 469444 596838
rect 469876 518226 469904 600086
rect 470600 587172 470652 587178
rect 470600 587114 470652 587120
rect 469864 518220 469916 518226
rect 469864 518162 469916 518168
rect 469416 402946 469536 402974
rect 469232 393286 469352 393314
rect 468576 388952 468628 388958
rect 468576 388894 468628 388900
rect 462884 385886 463358 385914
rect 463712 385886 464094 385914
rect 464264 385886 464830 385914
rect 465184 385886 465566 385914
rect 465920 385886 466302 385914
rect 466564 385886 467038 385914
rect 467392 385886 467774 385914
rect 468036 385886 468510 385914
rect 469232 385900 469260 393286
rect 469508 385914 469536 402946
rect 470612 389298 470640 587114
rect 470692 584452 470744 584458
rect 470692 584394 470744 584400
rect 470600 389292 470652 389298
rect 470600 389234 470652 389240
rect 469508 385886 469982 385914
rect 470704 385900 470732 584394
rect 476040 517614 476068 600086
rect 476028 517608 476080 517614
rect 476028 517550 476080 517556
rect 476040 516866 476068 517550
rect 482296 517478 482324 600100
rect 488644 598330 488672 600100
rect 488632 598324 488684 598330
rect 488632 598266 488684 598272
rect 494336 598324 494388 598330
rect 494336 598266 494388 598272
rect 493324 598256 493376 598262
rect 493324 598198 493376 598204
rect 482928 520940 482980 520946
rect 482928 520882 482980 520888
rect 482742 517576 482798 517585
rect 482940 517562 482968 520882
rect 488632 520328 488684 520334
rect 488632 520270 488684 520276
rect 488644 517970 488672 520270
rect 488644 517942 488980 517970
rect 482798 517534 483000 517562
rect 482742 517511 482798 517520
rect 482284 517472 482336 517478
rect 482284 517414 482336 517420
rect 476028 516860 476080 516866
rect 476028 516802 476080 516808
rect 492128 516792 492180 516798
rect 492128 516734 492180 516740
rect 492140 512650 492168 516734
rect 492128 512644 492180 512650
rect 492128 512586 492180 512592
rect 492140 512485 492168 512586
rect 492126 512476 492182 512485
rect 492126 512411 492182 512420
rect 480272 500126 480608 500154
rect 481652 500126 481804 500154
rect 482664 500126 483000 500154
rect 483860 500126 484196 500154
rect 485056 500126 485392 500154
rect 485792 500126 486588 500154
rect 487172 500126 487784 500154
rect 488980 500126 489224 500154
rect 480272 497690 480300 500126
rect 480260 497684 480312 497690
rect 480260 497626 480312 497632
rect 481652 497486 481680 500126
rect 482664 497758 482692 500126
rect 482652 497752 482704 497758
rect 482652 497694 482704 497700
rect 483860 497622 483888 500126
rect 483848 497616 483900 497622
rect 483848 497558 483900 497564
rect 485056 497554 485084 500126
rect 485044 497548 485096 497554
rect 485044 497490 485096 497496
rect 481640 497480 481692 497486
rect 481640 497422 481692 497428
rect 473726 462904 473782 462913
rect 473726 462839 473782 462848
rect 473740 454102 473768 462839
rect 480996 455524 481048 455530
rect 480996 455466 481048 455472
rect 473728 454096 473780 454102
rect 473728 454038 473780 454044
rect 473740 453900 473768 454038
rect 481008 453900 481036 455466
rect 485792 454782 485820 500126
rect 485780 454776 485832 454782
rect 485780 454718 485832 454724
rect 487172 454714 487200 500126
rect 489196 496913 489224 500126
rect 489932 500126 490176 500154
rect 491312 500126 491372 500154
rect 489182 496904 489238 496913
rect 489182 496839 489238 496848
rect 489932 457502 489960 500126
rect 489920 457496 489972 457502
rect 489920 457438 489972 457444
rect 488264 456068 488316 456074
rect 488264 456010 488316 456016
rect 488276 455462 488304 456010
rect 488264 455456 488316 455462
rect 488264 455398 488316 455404
rect 487160 454708 487212 454714
rect 487160 454650 487212 454656
rect 488276 453900 488304 455398
rect 471624 428466 471652 432140
rect 474292 430030 474320 432140
rect 474280 430024 474332 430030
rect 474280 429966 474332 429972
rect 476960 429962 476988 432140
rect 476948 429956 477000 429962
rect 476948 429898 477000 429904
rect 479628 429894 479656 432140
rect 479616 429888 479668 429894
rect 479616 429830 479668 429836
rect 482296 429214 482324 432140
rect 484964 429214 484992 432140
rect 487172 432126 487646 432154
rect 489932 432126 490314 432154
rect 480904 429208 480956 429214
rect 480904 429150 480956 429156
rect 482284 429208 482336 429214
rect 482284 429150 482336 429156
rect 483664 429208 483716 429214
rect 483664 429150 483716 429156
rect 484952 429208 485004 429214
rect 484952 429150 485004 429156
rect 476118 428496 476174 428505
rect 471612 428460 471664 428466
rect 476118 428431 476174 428440
rect 471612 428402 471664 428408
rect 476132 402974 476160 428431
rect 476132 402946 476896 402974
rect 471060 389292 471112 389298
rect 471060 389234 471112 389240
rect 471072 385914 471100 389234
rect 474372 389088 474424 389094
rect 472162 389056 472218 389065
rect 472162 388991 472218 389000
rect 473634 389056 473690 389065
rect 474372 389030 474424 389036
rect 473634 388991 473690 389000
rect 471072 385886 471454 385914
rect 472176 385900 472204 388991
rect 472898 388920 472954 388929
rect 472898 388855 472954 388864
rect 472912 385900 472940 388855
rect 473648 385900 473676 388991
rect 474384 385900 474412 389030
rect 475108 389020 475160 389026
rect 475108 388962 475160 388968
rect 475120 385900 475148 388962
rect 475844 388816 475896 388822
rect 475844 388758 475896 388764
rect 475856 385900 475884 388758
rect 476580 388680 476632 388686
rect 476580 388622 476632 388628
rect 476592 385900 476620 388622
rect 476868 385914 476896 402946
rect 480916 389910 480944 429150
rect 483676 395350 483704 429150
rect 487068 423360 487120 423366
rect 487068 423302 487120 423308
rect 484308 421592 484360 421598
rect 484308 421534 484360 421540
rect 483664 395344 483716 395350
rect 483664 395286 483716 395292
rect 484320 393314 484348 421534
rect 486976 416084 487028 416090
rect 486976 416026 487028 416032
rect 486988 393314 487016 416026
rect 483584 393286 484348 393314
rect 486896 393286 487016 393314
rect 480904 389904 480956 389910
rect 480904 389846 480956 389852
rect 479522 389056 479578 389065
rect 479522 388991 479578 389000
rect 478788 388952 478840 388958
rect 478788 388894 478840 388900
rect 478052 388748 478104 388754
rect 478052 388690 478104 388696
rect 476868 385886 477342 385914
rect 478064 385900 478092 388690
rect 478800 385900 478828 388894
rect 479536 385900 479564 388991
rect 480260 388884 480312 388890
rect 480260 388826 480312 388832
rect 480272 385900 480300 388826
rect 480996 388612 481048 388618
rect 480996 388554 481048 388560
rect 481008 385900 481036 388554
rect 481732 388544 481784 388550
rect 481732 388486 481784 388492
rect 481744 385900 481772 388486
rect 482468 388476 482520 388482
rect 482468 388418 482520 388424
rect 482480 385900 482508 388418
rect 483584 385914 483612 393286
rect 486424 389292 486476 389298
rect 486424 389234 486476 389240
rect 483940 388884 483992 388890
rect 483940 388826 483992 388832
rect 483230 385886 483612 385914
rect 483952 385900 483980 388826
rect 484676 388680 484728 388686
rect 484676 388622 484728 388628
rect 484688 385900 484716 388622
rect 485412 388612 485464 388618
rect 485412 388554 485464 388560
rect 485424 385900 485452 388554
rect 486436 385914 486464 389234
rect 486174 385886 486464 385914
rect 486896 385900 486924 393286
rect 487080 389298 487108 423302
rect 487172 392630 487200 432126
rect 488264 423292 488316 423298
rect 488264 423234 488316 423240
rect 488276 393314 488304 423234
rect 489644 423224 489696 423230
rect 489644 423166 489696 423172
rect 489656 393314 489684 423166
rect 488000 393286 488304 393314
rect 489472 393286 489684 393314
rect 487160 392624 487212 392630
rect 487160 392566 487212 392572
rect 487068 389292 487120 389298
rect 487068 389234 487120 389240
rect 488000 385914 488028 393286
rect 488356 388476 488408 388482
rect 488356 388418 488408 388424
rect 487646 385886 488028 385914
rect 488368 385900 488396 388418
rect 489472 385914 489500 393286
rect 489932 389842 489960 432126
rect 489920 389836 489972 389842
rect 489920 389778 489972 389784
rect 490564 389836 490616 389842
rect 490564 389778 490616 389784
rect 489828 388544 489880 388550
rect 489828 388486 489880 388492
rect 489118 385886 489500 385914
rect 489840 385900 489868 388486
rect 490576 385900 490604 389778
rect 491312 387190 491340 500126
rect 493140 396772 493192 396778
rect 493140 396714 493192 396720
rect 492404 395344 492456 395350
rect 492404 395286 492456 395292
rect 491576 392624 491628 392630
rect 491576 392566 491628 392572
rect 491300 387184 491352 387190
rect 491300 387126 491352 387132
rect 491588 385914 491616 392566
rect 492416 385914 492444 395286
rect 493152 385914 493180 396714
rect 493336 395321 493364 598198
rect 494244 518220 494296 518226
rect 494244 518162 494296 518168
rect 494152 517608 494204 517614
rect 494152 517550 494204 517556
rect 494164 508881 494192 517550
rect 494150 508872 494206 508881
rect 494150 508807 494206 508816
rect 494164 508570 494192 508807
rect 494152 508564 494204 508570
rect 494152 508506 494204 508512
rect 494256 505753 494284 518162
rect 494348 517546 494376 598266
rect 494992 596834 495020 600100
rect 500972 600086 501354 600114
rect 507136 600086 507702 600114
rect 513392 600086 514050 600114
rect 520292 600086 520398 600114
rect 494980 596828 495032 596834
rect 494980 596770 495032 596776
rect 494336 517540 494388 517546
rect 494336 517482 494388 517488
rect 494348 515953 494376 517482
rect 500972 516905 501000 600086
rect 500958 516896 501014 516905
rect 500958 516831 501014 516840
rect 502246 516896 502302 516905
rect 502246 516831 502302 516840
rect 494334 515944 494390 515953
rect 494334 515879 494390 515888
rect 494348 509930 494376 515879
rect 502260 514078 502288 516831
rect 507136 516769 507164 600086
rect 511264 576904 511316 576910
rect 511264 576846 511316 576852
rect 507122 516760 507178 516769
rect 507122 516695 507178 516704
rect 502248 514072 502300 514078
rect 502248 514014 502300 514020
rect 494336 509924 494388 509930
rect 494336 509866 494388 509872
rect 495072 505776 495124 505782
rect 494242 505744 494298 505753
rect 494242 505679 494298 505688
rect 495070 505744 495072 505753
rect 495124 505744 495126 505753
rect 495070 505679 495126 505688
rect 494702 501256 494758 501265
rect 494702 501191 494758 501200
rect 494716 462466 494744 501191
rect 494704 462460 494756 462466
rect 494704 462402 494756 462408
rect 494716 456074 494744 462402
rect 494704 456068 494756 456074
rect 494704 456010 494756 456016
rect 502984 423428 503036 423434
rect 502984 423370 503036 423376
rect 498108 423156 498160 423162
rect 498108 423098 498160 423104
rect 495348 420232 495400 420238
rect 495348 420174 495400 420180
rect 494612 399492 494664 399498
rect 494612 399434 494664 399440
rect 493968 398132 494020 398138
rect 493968 398074 494020 398080
rect 493322 395312 493378 395321
rect 493322 395247 493378 395256
rect 493980 385914 494008 398074
rect 494624 385914 494652 399434
rect 495360 385914 495388 420174
rect 497924 400920 497976 400926
rect 497924 400862 497976 400868
rect 496728 394052 496780 394058
rect 496728 393994 496780 394000
rect 495716 391332 495768 391338
rect 495716 391274 495768 391280
rect 491326 385886 491616 385914
rect 492062 385886 492444 385914
rect 492798 385886 493180 385914
rect 493534 385886 494008 385914
rect 494270 385886 494652 385914
rect 495006 385886 495388 385914
rect 495728 385900 495756 391274
rect 496740 385914 496768 393994
rect 497464 389292 497516 389298
rect 497464 389234 497516 389240
rect 497476 385914 497504 389234
rect 496478 385886 496768 385914
rect 497214 385886 497504 385914
rect 497936 385900 497964 400862
rect 498120 389298 498148 423098
rect 499304 423088 499356 423094
rect 499304 423030 499356 423036
rect 499316 393314 499344 423030
rect 500684 423020 500736 423026
rect 500684 422962 500736 422968
rect 500696 393314 500724 422962
rect 502248 422952 502300 422958
rect 502248 422894 502300 422900
rect 502260 393314 502288 422894
rect 499040 393286 499344 393314
rect 500512 393286 500724 393314
rect 501984 393286 502288 393314
rect 498108 389292 498160 389298
rect 498108 389234 498160 389240
rect 499040 385914 499068 393286
rect 499396 388816 499448 388822
rect 499396 388758 499448 388764
rect 498686 385886 499068 385914
rect 499408 385900 499436 388758
rect 500512 385914 500540 393286
rect 500868 388748 500920 388754
rect 500868 388690 500920 388696
rect 500158 385886 500540 385914
rect 500880 385900 500908 388690
rect 501984 385914 502012 393286
rect 502340 388952 502392 388958
rect 502340 388894 502392 388900
rect 501630 385886 502012 385914
rect 502352 385900 502380 388894
rect 502996 388890 503024 423370
rect 506480 417784 506532 417790
rect 506480 417726 506532 417732
rect 503720 417716 503772 417722
rect 503720 417658 503772 417664
rect 503444 402280 503496 402286
rect 503444 402222 503496 402228
rect 502984 388884 503036 388890
rect 502984 388826 503036 388832
rect 503456 385914 503484 402222
rect 503102 385886 503484 385914
rect 503732 385914 503760 417658
rect 503996 417512 504048 417518
rect 503996 417454 504048 417460
rect 504008 402974 504036 417454
rect 504008 402946 504128 402974
rect 504100 385914 504128 402946
rect 505560 393984 505612 393990
rect 505560 393926 505612 393932
rect 505284 391264 505336 391270
rect 505284 391206 505336 391212
rect 503732 385886 503838 385914
rect 504100 385886 504574 385914
rect 505296 385900 505324 391206
rect 505572 385914 505600 393926
rect 506492 389298 506520 417726
rect 507860 417648 507912 417654
rect 507860 417590 507912 417596
rect 506572 417444 506624 417450
rect 506572 417386 506624 417392
rect 506480 389292 506532 389298
rect 506480 389234 506532 389240
rect 506584 385914 506612 417386
rect 507872 389298 507900 417590
rect 507952 417580 508004 417586
rect 507952 417522 508004 417528
rect 507124 389292 507176 389298
rect 507124 389234 507176 389240
rect 507860 389292 507912 389298
rect 507860 389234 507912 389240
rect 507136 385914 507164 389234
rect 507964 385914 507992 417522
rect 508596 389292 508648 389298
rect 508596 389234 508648 389240
rect 508608 385914 508636 389234
rect 505572 385886 506046 385914
rect 506584 385886 506782 385914
rect 507136 385886 507518 385914
rect 507964 385886 508254 385914
rect 508608 385886 508990 385914
rect 457352 385688 457404 385694
rect 457352 385630 457404 385636
rect 452016 385416 452068 385422
rect 452016 385358 452068 385364
rect 509330 365256 509386 365265
rect 509330 365191 509386 365200
rect 450728 336796 450780 336802
rect 450728 336738 450780 336744
rect 450464 335326 450584 335354
rect 450556 334257 450584 335326
rect 450542 334248 450598 334257
rect 450542 334183 450598 334192
rect 450450 328672 450506 328681
rect 450450 328607 450506 328616
rect 450464 328506 450492 328607
rect 450452 328500 450504 328506
rect 450452 328442 450504 328448
rect 450556 327321 450584 334183
rect 450740 330546 450768 336738
rect 450728 330540 450780 330546
rect 450728 330482 450780 330488
rect 450542 327312 450598 327321
rect 450542 327247 450598 327256
rect 509344 326466 509372 365191
rect 510618 359136 510674 359145
rect 510618 359071 510674 359080
rect 509514 357640 509570 357649
rect 509514 357575 509570 357584
rect 509422 356144 509478 356153
rect 509422 356079 509478 356088
rect 509332 326460 509384 326466
rect 509332 326402 509384 326408
rect 509436 326398 509464 356079
rect 509424 326392 509476 326398
rect 509424 326334 509476 326340
rect 450372 325666 450768 325694
rect 450648 325553 450676 325666
rect 450634 325544 450690 325553
rect 450634 325479 450690 325488
rect 450174 325272 450230 325281
rect 450174 325207 450230 325216
rect 450542 324864 450598 324873
rect 450542 324799 450598 324808
rect 450082 324592 450138 324601
rect 450082 324527 450138 324536
rect 449808 263560 449860 263566
rect 449808 263502 449860 263508
rect 450556 221474 450584 324799
rect 450634 324184 450690 324193
rect 450634 324119 450690 324128
rect 450544 221468 450596 221474
rect 450544 221410 450596 221416
rect 450648 207670 450676 324119
rect 450740 235278 450768 325666
rect 509422 325000 509478 325009
rect 509422 324935 509478 324944
rect 509330 322960 509386 322969
rect 509330 322895 509386 322904
rect 473314 322788 473366 322794
rect 473314 322730 473366 322736
rect 459652 322720 459704 322726
rect 459494 322668 459652 322674
rect 459494 322662 459704 322668
rect 461308 322720 461360 322726
rect 461308 322662 461360 322668
rect 462226 322688 462282 322697
rect 459494 322646 459692 322662
rect 459100 322584 459152 322590
rect 458638 322552 458694 322561
rect 458942 322532 459100 322538
rect 461320 322561 461348 322662
rect 462226 322623 462282 322632
rect 462964 322652 463016 322658
rect 462964 322594 463016 322600
rect 458942 322526 459152 322532
rect 461306 322552 461362 322561
rect 458942 322510 459140 322526
rect 458638 322487 458694 322496
rect 461306 322487 461362 322496
rect 451832 320884 451884 320890
rect 451832 320826 451884 320832
rect 451844 320770 451872 320826
rect 451844 320754 451964 320770
rect 451844 320748 451976 320754
rect 451844 320742 451924 320748
rect 451924 320690 451976 320696
rect 454684 318232 454736 318238
rect 454684 318174 454736 318180
rect 451924 318164 451976 318170
rect 451924 318106 451976 318112
rect 450728 235272 450780 235278
rect 450728 235214 450780 235220
rect 450636 207664 450688 207670
rect 450636 207606 450688 207612
rect 448428 164212 448480 164218
rect 448428 164154 448480 164160
rect 449348 164212 449400 164218
rect 449348 164154 449400 164160
rect 448336 161424 448388 161430
rect 448336 161366 448388 161372
rect 448348 160750 448376 161366
rect 448336 160744 448388 160750
rect 448336 160686 448388 160692
rect 448440 159882 448468 164154
rect 450544 161628 450596 161634
rect 450544 161570 450596 161576
rect 444912 159854 445248 159882
rect 448224 159854 448468 159882
rect 437952 159594 438624 159610
rect 437940 159588 438624 159594
rect 437992 159582 438624 159588
rect 437940 159530 437992 159536
rect 437572 159520 437624 159526
rect 437572 159462 437624 159468
rect 421392 159310 421880 159338
rect 425152 159384 425204 159390
rect 425152 159326 425204 159332
rect 410524 156664 410576 156670
rect 410524 156606 410576 156612
rect 409512 150408 409564 150414
rect 409512 150350 409564 150356
rect 409420 147688 409472 147694
rect 409420 147630 409472 147636
rect 450556 142186 450584 161570
rect 450636 161560 450688 161566
rect 450636 161502 450688 161508
rect 450648 142254 450676 161502
rect 451740 158296 451792 158302
rect 451738 158264 451740 158273
rect 451792 158264 451794 158273
rect 451738 158199 451794 158208
rect 451740 157344 451792 157350
rect 451740 157286 451792 157292
rect 451752 156913 451780 157286
rect 451738 156904 451794 156913
rect 451738 156839 451794 156848
rect 451936 155553 451964 318106
rect 452016 308508 452068 308514
rect 452016 308450 452068 308456
rect 451922 155544 451978 155553
rect 451922 155479 451978 155488
rect 451924 154216 451976 154222
rect 451922 154184 451924 154193
rect 451976 154184 451978 154193
rect 451922 154119 451978 154128
rect 452028 151473 452056 308450
rect 452108 286680 452160 286686
rect 452108 286622 452160 286628
rect 452014 151464 452070 151473
rect 452014 151399 452070 151408
rect 451740 147416 451792 147422
rect 451738 147384 451740 147393
rect 451792 147384 451794 147393
rect 451738 147319 451794 147328
rect 451464 144832 451516 144838
rect 451464 144774 451516 144780
rect 451476 144673 451504 144774
rect 451462 144664 451518 144673
rect 451462 144599 451518 144608
rect 450636 142248 450688 142254
rect 450636 142190 450688 142196
rect 450544 142180 450596 142186
rect 450544 142122 450596 142128
rect 409328 139392 409380 139398
rect 409328 139334 409380 139340
rect 409236 128308 409288 128314
rect 409236 128250 409288 128256
rect 450556 106962 450584 142122
rect 450648 117298 450676 142190
rect 452120 132433 452148 286622
rect 453304 284980 453356 284986
rect 453304 284922 453356 284928
rect 452384 283620 452436 283626
rect 452384 283562 452436 283568
rect 452200 273964 452252 273970
rect 452200 273906 452252 273912
rect 452106 132424 452162 132433
rect 452106 132359 452162 132368
rect 452212 131322 452240 273906
rect 452292 268524 452344 268530
rect 452292 268466 452344 268472
rect 452120 131294 452240 131322
rect 451740 126404 451792 126410
rect 451740 126346 451792 126352
rect 451752 125633 451780 126346
rect 451738 125624 451794 125633
rect 451738 125559 451794 125568
rect 452120 124273 452148 131294
rect 452304 131186 452332 268466
rect 452396 152833 452424 283562
rect 452382 152824 452438 152833
rect 452382 152759 452438 152768
rect 452476 150272 452528 150278
rect 452476 150214 452528 150220
rect 452488 150113 452516 150214
rect 452474 150104 452530 150113
rect 452474 150039 452530 150048
rect 452568 148776 452620 148782
rect 452566 148744 452568 148753
rect 452620 148744 452622 148753
rect 452566 148679 452622 148688
rect 452568 146056 452620 146062
rect 452566 146024 452568 146033
rect 452620 146024 452622 146033
rect 452566 145959 452622 145968
rect 452568 143336 452620 143342
rect 452566 143304 452568 143313
rect 452620 143304 452622 143313
rect 452566 143239 452622 143248
rect 452568 141976 452620 141982
rect 452566 141944 452568 141953
rect 452620 141944 452622 141953
rect 452566 141879 452622 141888
rect 452568 140616 452620 140622
rect 452566 140584 452568 140593
rect 452620 140584 452622 140593
rect 452566 140519 452622 140528
rect 452568 139256 452620 139262
rect 452566 139224 452568 139233
rect 452620 139224 452622 139233
rect 452566 139159 452622 139168
rect 452568 137896 452620 137902
rect 452566 137864 452568 137873
rect 452620 137864 452622 137873
rect 452566 137799 452622 137808
rect 452568 136536 452620 136542
rect 452566 136504 452568 136513
rect 452620 136504 452622 136513
rect 452566 136439 452622 136448
rect 452568 135176 452620 135182
rect 452566 135144 452568 135153
rect 452620 135144 452622 135153
rect 452566 135079 452622 135088
rect 452568 133816 452620 133822
rect 452566 133784 452568 133793
rect 452620 133784 452622 133793
rect 452566 133719 452622 133728
rect 452212 131158 452332 131186
rect 452212 128353 452240 131158
rect 452292 131096 452344 131102
rect 452290 131064 452292 131073
rect 452344 131064 452346 131073
rect 452290 130999 452346 131008
rect 452384 129736 452436 129742
rect 452382 129704 452384 129713
rect 452436 129704 452438 129713
rect 452382 129639 452438 129648
rect 452198 128344 452254 128353
rect 452198 128279 452254 128288
rect 452290 126984 452346 126993
rect 453316 126954 453344 284922
rect 453672 279540 453724 279546
rect 453672 279482 453724 279488
rect 453396 279472 453448 279478
rect 453396 279414 453448 279420
rect 453408 131102 453436 279414
rect 453488 278112 453540 278118
rect 453488 278054 453540 278060
rect 453396 131096 453448 131102
rect 453396 131038 453448 131044
rect 453500 129742 453528 278054
rect 453580 272604 453632 272610
rect 453580 272546 453632 272552
rect 453488 129736 453540 129742
rect 453488 129678 453540 129684
rect 452290 126919 452292 126928
rect 452344 126919 452346 126928
rect 453304 126948 453356 126954
rect 452292 126890 452344 126896
rect 453304 126890 453356 126896
rect 453592 126410 453620 272546
rect 453684 262886 453712 279482
rect 453948 263628 454000 263634
rect 453948 263570 454000 263576
rect 453672 262880 453724 262886
rect 453672 262822 453724 262828
rect 453960 258126 453988 263570
rect 453948 258120 454000 258126
rect 453948 258062 454000 258068
rect 453580 126404 453632 126410
rect 453580 126346 453632 126352
rect 452106 124264 452162 124273
rect 452106 124199 452162 124208
rect 451832 124160 451884 124166
rect 451832 124102 451884 124108
rect 451844 122913 451872 124102
rect 451830 122904 451886 122913
rect 451830 122839 451886 122848
rect 454696 122262 454724 318174
rect 455892 315314 455920 322116
rect 456182 322102 456380 322130
rect 456458 322102 456656 322130
rect 456062 321872 456118 321881
rect 456062 321807 456118 321816
rect 455880 315308 455932 315314
rect 455880 315250 455932 315256
rect 454776 314016 454828 314022
rect 454776 313958 454828 313964
rect 454788 137902 454816 313958
rect 454960 309868 455012 309874
rect 454960 309810 455012 309816
rect 454868 307216 454920 307222
rect 454868 307158 454920 307164
rect 454776 137896 454828 137902
rect 454776 137838 454828 137844
rect 454880 133822 454908 307158
rect 454972 148782 455000 309810
rect 455052 280832 455104 280838
rect 455052 280774 455104 280780
rect 454960 148776 455012 148782
rect 454960 148718 455012 148724
rect 455064 144838 455092 280774
rect 455236 276684 455288 276690
rect 455236 276626 455288 276632
rect 455144 272536 455196 272542
rect 455144 272478 455196 272484
rect 455052 144832 455104 144838
rect 455052 144774 455104 144780
rect 455156 141982 455184 272478
rect 455248 154222 455276 276626
rect 455236 154216 455288 154222
rect 455236 154158 455288 154164
rect 455144 141976 455196 141982
rect 455144 141918 455196 141924
rect 454868 133816 454920 133822
rect 454868 133758 454920 133764
rect 451740 122256 451792 122262
rect 451740 122198 451792 122204
rect 454684 122256 454736 122262
rect 454684 122198 454736 122204
rect 451752 121553 451780 122198
rect 451738 121544 451794 121553
rect 451738 121479 451794 121488
rect 456076 119406 456104 321807
rect 456352 303414 456380 322102
rect 456340 303408 456392 303414
rect 456340 303350 456392 303356
rect 456628 301646 456656 322102
rect 456616 301640 456668 301646
rect 456616 301582 456668 301588
rect 456720 298042 456748 322116
rect 457010 322102 457208 322130
rect 457286 322102 457484 322130
rect 457562 322102 457760 322130
rect 457180 308446 457208 322102
rect 457456 316130 457484 322102
rect 457444 316124 457496 316130
rect 457444 316066 457496 316072
rect 457444 315376 457496 315382
rect 457444 315318 457496 315324
rect 457168 308440 457220 308446
rect 457168 308382 457220 308388
rect 456708 298036 456760 298042
rect 456708 297978 456760 297984
rect 456248 271108 456300 271114
rect 456248 271050 456300 271056
rect 456156 269884 456208 269890
rect 456156 269826 456208 269832
rect 456168 158302 456196 269826
rect 456260 243574 456288 271050
rect 456708 269952 456760 269958
rect 456708 269894 456760 269900
rect 456720 262954 456748 269894
rect 456892 266416 456944 266422
rect 456892 266358 456944 266364
rect 456904 263634 456932 266358
rect 456892 263628 456944 263634
rect 456892 263570 456944 263576
rect 456800 263560 456852 263566
rect 456800 263502 456852 263508
rect 456708 262948 456760 262954
rect 456708 262890 456760 262896
rect 456812 262721 456840 263502
rect 456798 262712 456854 262721
rect 456798 262647 456854 262656
rect 456892 250980 456944 250986
rect 456892 250922 456944 250928
rect 456800 249756 456852 249762
rect 456800 249698 456852 249704
rect 456812 248849 456840 249698
rect 456798 248840 456854 248849
rect 456798 248775 456854 248784
rect 456904 247722 456932 250922
rect 456892 247716 456944 247722
rect 456892 247658 456944 247664
rect 456248 243568 456300 243574
rect 456248 243510 456300 243516
rect 456800 235272 456852 235278
rect 456800 235214 456852 235220
rect 456812 234977 456840 235214
rect 456798 234968 456854 234977
rect 456798 234903 456854 234912
rect 456156 158296 456208 158302
rect 456156 158238 456208 158244
rect 457456 136542 457484 315318
rect 457536 299940 457588 299946
rect 457536 299882 457588 299888
rect 457548 157350 457576 299882
rect 457732 294506 457760 322102
rect 457824 317082 457852 322116
rect 458100 321570 458128 322116
rect 458088 321564 458140 321570
rect 458088 321506 458140 321512
rect 458376 321502 458404 322116
rect 459218 322114 459416 322130
rect 459218 322108 459428 322114
rect 459218 322102 459376 322108
rect 459770 322102 459968 322130
rect 459376 322050 459428 322056
rect 458364 321496 458416 321502
rect 458364 321438 458416 321444
rect 459940 320890 459968 322102
rect 460032 321473 460060 322116
rect 460018 321464 460074 321473
rect 460018 321399 460074 321408
rect 459928 320884 459980 320890
rect 459928 320826 459980 320832
rect 460308 320006 460336 322116
rect 460584 320074 460612 322116
rect 460754 322008 460810 322017
rect 460754 321943 460810 321952
rect 460664 321020 460716 321026
rect 460664 320962 460716 320968
rect 460572 320068 460624 320074
rect 460572 320010 460624 320016
rect 460296 320000 460348 320006
rect 460296 319942 460348 319948
rect 460296 319456 460348 319462
rect 460202 319424 460258 319433
rect 460296 319398 460348 319404
rect 460202 319359 460258 319368
rect 457812 317076 457864 317082
rect 457812 317018 457864 317024
rect 458916 316736 458968 316742
rect 458916 316678 458968 316684
rect 457996 316124 458048 316130
rect 457996 316066 458048 316072
rect 458008 296002 458036 316066
rect 458824 305448 458876 305454
rect 458824 305390 458876 305396
rect 457996 295996 458048 296002
rect 457996 295938 458048 295944
rect 457720 294500 457772 294506
rect 457720 294442 457772 294448
rect 457628 274032 457680 274038
rect 457628 273974 457680 273980
rect 457536 157344 457588 157350
rect 457536 157286 457588 157292
rect 457640 140622 457668 273974
rect 457720 271176 457772 271182
rect 457720 271118 457772 271124
rect 457732 147422 457760 271118
rect 457810 234968 457866 234977
rect 457810 234903 457866 234912
rect 457824 162246 457852 234903
rect 457904 221468 457956 221474
rect 457904 221410 457956 221416
rect 457916 221105 457944 221410
rect 457902 221096 457958 221105
rect 457902 221031 457958 221040
rect 457812 162240 457864 162246
rect 457812 162182 457864 162188
rect 457916 162178 457944 221031
rect 457904 162172 457956 162178
rect 457904 162114 457956 162120
rect 457720 147416 457772 147422
rect 457720 147358 457772 147364
rect 457628 140616 457680 140622
rect 457628 140558 457680 140564
rect 457444 136536 457496 136542
rect 457444 136478 457496 136484
rect 458836 124166 458864 305390
rect 458928 135182 458956 316678
rect 459008 311228 459060 311234
rect 459008 311170 459060 311176
rect 459020 146062 459048 311170
rect 459376 304156 459428 304162
rect 459376 304098 459428 304104
rect 459284 282192 459336 282198
rect 459284 282134 459336 282140
rect 459192 275324 459244 275330
rect 459192 275266 459244 275272
rect 459100 271244 459152 271250
rect 459100 271186 459152 271192
rect 459008 146056 459060 146062
rect 459008 145998 459060 146004
rect 459112 139262 459140 271186
rect 459204 143342 459232 275266
rect 459296 150278 459324 282134
rect 459388 250986 459416 304098
rect 459468 282940 459520 282946
rect 459468 282882 459520 282888
rect 459480 271114 459508 282882
rect 459468 271108 459520 271114
rect 459468 271050 459520 271056
rect 459560 268592 459612 268598
rect 459560 268534 459612 268540
rect 459572 266422 459600 268534
rect 459560 266416 459612 266422
rect 459560 266358 459612 266364
rect 459376 250980 459428 250986
rect 459376 250922 459428 250928
rect 459560 207664 459612 207670
rect 459560 207606 459612 207612
rect 460020 207664 460072 207670
rect 460020 207606 460072 207612
rect 459572 161498 459600 207606
rect 460032 207369 460060 207606
rect 460018 207360 460074 207369
rect 460018 207295 460074 207304
rect 459560 161492 459612 161498
rect 459560 161434 459612 161440
rect 459284 150272 459336 150278
rect 459284 150214 459336 150220
rect 459192 143336 459244 143342
rect 459192 143278 459244 143284
rect 459100 139256 459152 139262
rect 459100 139198 459152 139204
rect 458916 135176 458968 135182
rect 458916 135118 458968 135124
rect 458824 124160 458876 124166
rect 458824 124102 458876 124108
rect 456064 119400 456116 119406
rect 456064 119342 456116 119348
rect 450636 117292 450688 117298
rect 450636 117234 450688 117240
rect 450544 106956 450596 106962
rect 450544 106898 450596 106904
rect 409144 106276 409196 106282
rect 409144 106218 409196 106224
rect 389528 104910 389864 104938
rect 386236 95192 386288 95198
rect 386236 95134 386288 95140
rect 386144 62076 386196 62082
rect 386144 62018 386196 62024
rect 386144 51128 386196 51134
rect 386144 51070 386196 51076
rect 386052 33924 386104 33930
rect 386052 33866 386104 33872
rect 385960 33788 386012 33794
rect 385960 33730 386012 33736
rect 386156 31686 386184 51070
rect 386144 31680 386196 31686
rect 386144 31622 386196 31628
rect 385868 31068 385920 31074
rect 385868 31010 385920 31016
rect 385774 3768 385830 3777
rect 385774 3703 385830 3712
rect 381726 3431 381782 3440
rect 385684 3460 385736 3466
rect 385684 3402 385736 3408
rect 460216 3369 460244 319359
rect 460308 31754 460336 319398
rect 460388 296744 460440 296750
rect 460388 296686 460440 296692
rect 460400 282946 460428 296686
rect 460388 282940 460440 282946
rect 460388 282882 460440 282888
rect 460676 200734 460704 320962
rect 460664 200728 460716 200734
rect 460664 200670 460716 200676
rect 460768 200138 460796 321943
rect 460860 321434 460888 322116
rect 460848 321428 460900 321434
rect 460848 321370 460900 321376
rect 461136 319870 461164 322116
rect 461412 320754 461440 322116
rect 461688 321366 461716 322116
rect 461676 321360 461728 321366
rect 461676 321302 461728 321308
rect 461964 321065 461992 322116
rect 462516 321337 462544 322116
rect 462502 321328 462558 321337
rect 462502 321263 462558 321272
rect 461950 321056 462006 321065
rect 461950 320991 462006 321000
rect 461400 320748 461452 320754
rect 461400 320690 461452 320696
rect 461124 319864 461176 319870
rect 461124 319806 461176 319812
rect 462792 319598 462820 322116
rect 462976 322114 463004 322594
rect 469036 322584 469088 322590
rect 473326 322538 473354 322730
rect 473452 322720 473504 322726
rect 480628 322720 480680 322726
rect 473452 322662 473504 322668
rect 480470 322668 480628 322674
rect 480470 322662 480680 322668
rect 480994 322688 481050 322697
rect 473464 322561 473492 322662
rect 478144 322652 478196 322658
rect 480470 322646 480668 322662
rect 480904 322652 480956 322658
rect 478144 322594 478196 322600
rect 480994 322623 481050 322632
rect 480904 322594 480956 322600
rect 469088 322532 469154 322538
rect 469036 322526 469154 322532
rect 469048 322510 469154 322526
rect 473294 322510 473354 322538
rect 473450 322552 473506 322561
rect 473450 322487 473506 322496
rect 473452 322448 473504 322454
rect 473450 322416 473452 322425
rect 473504 322416 473506 322425
rect 473450 322351 473506 322360
rect 478156 322318 478184 322594
rect 480628 322584 480680 322590
rect 480916 322561 480944 322594
rect 480628 322526 480680 322532
rect 480902 322552 480958 322561
rect 480640 322318 480668 322526
rect 480902 322487 480958 322496
rect 507400 322516 507452 322522
rect 507400 322458 507452 322464
rect 481546 322416 481602 322425
rect 482296 322386 482402 322402
rect 481546 322351 481602 322360
rect 482284 322380 482402 322386
rect 482336 322374 482402 322380
rect 482284 322322 482336 322328
rect 463792 322312 463844 322318
rect 473452 322312 473504 322318
rect 463844 322260 463910 322266
rect 463792 322254 463910 322260
rect 478144 322312 478196 322318
rect 473504 322260 473570 322266
rect 473452 322254 473570 322260
rect 463804 322238 463910 322254
rect 473464 322238 473570 322254
rect 474292 322250 474398 322266
rect 474280 322244 474398 322250
rect 474332 322238 474398 322244
rect 474950 322250 475148 322266
rect 478144 322254 478196 322260
rect 480628 322312 480680 322318
rect 506940 322312 506992 322318
rect 480628 322254 480680 322260
rect 490130 322250 490328 322266
rect 506940 322254 506992 322260
rect 474950 322244 475160 322250
rect 474950 322238 475108 322244
rect 474280 322186 474332 322192
rect 475108 322186 475160 322192
rect 475384 322244 475436 322250
rect 490130 322244 490340 322250
rect 490130 322238 490288 322244
rect 475384 322186 475436 322192
rect 490288 322186 490340 322192
rect 490564 322244 490616 322250
rect 490564 322186 490616 322192
rect 462964 322108 463016 322114
rect 462964 322050 463016 322056
rect 463068 320618 463096 322116
rect 463344 321162 463372 322116
rect 463332 321156 463384 321162
rect 463332 321098 463384 321104
rect 463056 320612 463108 320618
rect 463056 320554 463108 320560
rect 463620 319938 463648 322116
rect 463608 319932 463660 319938
rect 463608 319874 463660 319880
rect 462780 319592 462832 319598
rect 462780 319534 462832 319540
rect 464068 319048 464120 319054
rect 464068 318990 464120 318996
rect 463792 318980 463844 318986
rect 463792 318922 463844 318928
rect 461584 317076 461636 317082
rect 461584 317018 461636 317024
rect 461596 299470 461624 317018
rect 462964 311160 463016 311166
rect 462964 311102 463016 311108
rect 461676 310344 461728 310350
rect 461676 310286 461728 310292
rect 461688 304162 461716 310286
rect 461676 304156 461728 304162
rect 461676 304098 461728 304104
rect 461584 299464 461636 299470
rect 461584 299406 461636 299412
rect 462976 296750 463004 311102
rect 463804 306202 463832 318922
rect 463792 306196 463844 306202
rect 463792 306138 463844 306144
rect 464080 302734 464108 318990
rect 464172 310350 464200 322116
rect 464356 322102 464462 322130
rect 464632 322102 464738 322130
rect 464908 322102 465014 322130
rect 464356 311166 464384 322102
rect 464632 319054 464660 322102
rect 464620 319048 464672 319054
rect 464620 318990 464672 318996
rect 464908 318986 464936 322102
rect 465172 319048 465224 319054
rect 465172 318990 465224 318996
rect 464896 318980 464948 318986
rect 464896 318922 464948 318928
rect 464344 311160 464396 311166
rect 464344 311102 464396 311108
rect 464160 310344 464212 310350
rect 464160 310286 464212 310292
rect 465184 305522 465212 318990
rect 465276 316034 465304 322116
rect 465448 316124 465500 316130
rect 465448 316066 465500 316072
rect 465276 316006 465396 316034
rect 465368 306270 465396 316006
rect 465460 306338 465488 316066
rect 465448 306332 465500 306338
rect 465448 306274 465500 306280
rect 465356 306264 465408 306270
rect 465356 306206 465408 306212
rect 465552 305590 465580 322116
rect 465736 322102 465842 322130
rect 466012 322102 466118 322130
rect 465736 319054 465764 322102
rect 465724 319048 465776 319054
rect 465724 318990 465776 318996
rect 466012 316130 466040 322102
rect 466000 316124 466052 316130
rect 466000 316066 466052 316072
rect 465540 305584 465592 305590
rect 465540 305526 465592 305532
rect 465172 305516 465224 305522
rect 465172 305458 465224 305464
rect 464068 302728 464120 302734
rect 464068 302670 464120 302676
rect 462964 296744 463016 296750
rect 462964 296686 463016 296692
rect 461400 286748 461452 286754
rect 461400 286690 461452 286696
rect 461412 279546 461440 286690
rect 461400 279540 461452 279546
rect 461400 279482 461452 279488
rect 466380 268462 466408 322116
rect 466670 322102 466868 322130
rect 466946 322102 467144 322130
rect 466840 319054 466868 322102
rect 466828 319048 466880 319054
rect 466828 318990 466880 318996
rect 467116 318986 467144 322102
rect 467104 318980 467156 318986
rect 467104 318922 467156 318928
rect 467208 316034 467236 322116
rect 467380 319048 467432 319054
rect 467380 318990 467432 318996
rect 467208 316006 467328 316034
rect 467300 288930 467328 316006
rect 467392 312594 467420 318990
rect 467484 316034 467512 322116
rect 467656 318980 467708 318986
rect 467656 318922 467708 318928
rect 467484 316006 467604 316034
rect 467380 312588 467432 312594
rect 467380 312530 467432 312536
rect 467576 293282 467604 316006
rect 467564 293276 467616 293282
rect 467564 293218 467616 293224
rect 467668 290494 467696 318922
rect 467760 300014 467788 322116
rect 468050 322102 468248 322130
rect 468326 322102 468524 322130
rect 468220 316034 468248 322102
rect 468496 319138 468524 322102
rect 468588 321434 468616 322116
rect 468576 321428 468628 321434
rect 468576 321370 468628 321376
rect 468864 319938 468892 322116
rect 468852 319932 468904 319938
rect 468852 319874 468904 319880
rect 469416 319870 469444 322116
rect 469692 320006 469720 322116
rect 469968 321366 469996 322116
rect 469956 321360 470008 321366
rect 469956 321302 470008 321308
rect 469680 320000 469732 320006
rect 469680 319942 469732 319948
rect 469404 319864 469456 319870
rect 469404 319806 469456 319812
rect 470244 319598 470272 322116
rect 470520 321337 470548 322116
rect 470506 321328 470562 321337
rect 470506 321263 470562 321272
rect 470232 319592 470284 319598
rect 470232 319534 470284 319540
rect 470796 319190 470824 322116
rect 471072 319802 471100 322116
rect 471060 319796 471112 319802
rect 471060 319738 471112 319744
rect 471348 319734 471376 322116
rect 471336 319728 471388 319734
rect 471624 319705 471652 322116
rect 471900 320958 471928 322116
rect 471888 320952 471940 320958
rect 471888 320894 471940 320900
rect 471336 319670 471388 319676
rect 471610 319696 471666 319705
rect 471610 319631 471666 319640
rect 472176 319394 472204 322116
rect 472452 320686 472480 322116
rect 472440 320680 472492 320686
rect 472440 320622 472492 320628
rect 472728 319977 472756 322116
rect 472714 319968 472770 319977
rect 472714 319903 472770 319912
rect 473004 319841 473032 322116
rect 472990 319832 473046 319841
rect 472990 319767 473046 319776
rect 472164 319388 472216 319394
rect 472164 319330 472216 319336
rect 473832 319326 473860 322116
rect 474108 319666 474136 322116
rect 474568 322102 474674 322130
rect 475120 322102 475226 322130
rect 474096 319660 474148 319666
rect 474096 319602 474148 319608
rect 473820 319320 473872 319326
rect 473820 319262 473872 319268
rect 470784 319184 470836 319190
rect 468496 319110 469076 319138
rect 470784 319126 470836 319132
rect 468220 316006 468800 316034
rect 467748 300008 467800 300014
rect 467748 299950 467800 299956
rect 467656 290488 467708 290494
rect 467656 290430 467708 290436
rect 467288 288924 467340 288930
rect 467288 288866 467340 288872
rect 468772 269822 468800 316006
rect 469048 313274 469076 319110
rect 474568 316034 474596 322102
rect 475120 319138 475148 322102
rect 473740 316006 474596 316034
rect 474844 319110 475148 319138
rect 469036 313268 469088 313274
rect 469036 313210 469088 313216
rect 471244 291712 471296 291718
rect 471244 291654 471296 291660
rect 471256 286754 471284 291654
rect 471244 286748 471296 286754
rect 471244 286690 471296 286696
rect 473360 274712 473412 274718
rect 473360 274654 473412 274660
rect 468760 269816 468812 269822
rect 468760 269758 468812 269764
rect 473372 268598 473400 274654
rect 473740 269958 473768 316006
rect 474004 307828 474056 307834
rect 474004 307770 474056 307776
rect 474016 291718 474044 307770
rect 474844 302802 474872 319110
rect 475108 319048 475160 319054
rect 475108 318990 475160 318996
rect 475120 306066 475148 318990
rect 475108 306060 475160 306066
rect 475108 306002 475160 306008
rect 475396 302870 475424 322186
rect 484216 322176 484268 322182
rect 475488 305998 475516 322116
rect 475672 322102 475778 322130
rect 475948 322102 476054 322130
rect 475672 319054 475700 322102
rect 475660 319048 475712 319054
rect 475660 318990 475712 318996
rect 475948 316034 475976 322102
rect 476316 319462 476344 322116
rect 476500 322102 476606 322130
rect 476882 322102 477080 322130
rect 477158 322102 477356 322130
rect 476304 319456 476356 319462
rect 476304 319398 476356 319404
rect 475672 316006 475976 316034
rect 475672 306134 475700 316006
rect 475660 306128 475712 306134
rect 475660 306070 475712 306076
rect 475476 305992 475528 305998
rect 475476 305934 475528 305940
rect 475384 302864 475436 302870
rect 475384 302806 475436 302812
rect 474832 302796 474884 302802
rect 474832 302738 474884 302744
rect 474004 291712 474056 291718
rect 474004 291654 474056 291660
rect 475384 287836 475436 287842
rect 475384 287778 475436 287784
rect 475396 274718 475424 287778
rect 476500 286618 476528 322102
rect 477052 313954 477080 322102
rect 477040 313948 477092 313954
rect 477040 313890 477092 313896
rect 477328 307154 477356 322102
rect 477316 307148 477368 307154
rect 477316 307090 477368 307096
rect 477420 305998 477448 322116
rect 477696 318102 477724 322116
rect 477986 322102 478184 322130
rect 478262 322102 478460 322130
rect 484268 322124 484334 322130
rect 484216 322118 484334 322124
rect 477684 318096 477736 318102
rect 477684 318038 477736 318044
rect 478156 311166 478184 322102
rect 478144 311160 478196 311166
rect 478144 311102 478196 311108
rect 477408 305992 477460 305998
rect 477408 305934 477460 305940
rect 478144 298988 478196 298994
rect 478144 298930 478196 298936
rect 478156 295390 478184 298930
rect 476856 295384 476908 295390
rect 476856 295326 476908 295332
rect 478144 295384 478196 295390
rect 478144 295326 478196 295332
rect 476868 287842 476896 295326
rect 478432 291718 478460 322102
rect 478524 317422 478552 322116
rect 478800 319666 478828 322116
rect 479076 321162 479104 322116
rect 479352 321298 479380 322116
rect 479340 321292 479392 321298
rect 479340 321234 479392 321240
rect 479064 321156 479116 321162
rect 479064 321098 479116 321104
rect 479628 319734 479656 322116
rect 479904 320142 479932 322116
rect 479892 320136 479944 320142
rect 479892 320078 479944 320084
rect 480180 319802 480208 322116
rect 480732 320074 480760 322116
rect 481284 320482 481312 322116
rect 481836 320822 481864 322116
rect 481824 320816 481876 320822
rect 481824 320758 481876 320764
rect 482112 320550 482140 322116
rect 482664 321201 482692 322116
rect 482650 321192 482706 321201
rect 482650 321127 482706 321136
rect 482100 320544 482152 320550
rect 482100 320486 482152 320492
rect 481272 320476 481324 320482
rect 481272 320418 481324 320424
rect 480720 320068 480772 320074
rect 480720 320010 480772 320016
rect 480168 319796 480220 319802
rect 480168 319738 480220 319744
rect 479616 319728 479668 319734
rect 479616 319670 479668 319676
rect 478788 319660 478840 319666
rect 478788 319602 478840 319608
rect 482940 319258 482968 322116
rect 483216 320113 483244 322116
rect 483202 320104 483258 320113
rect 483202 320039 483258 320048
rect 483492 319530 483520 322116
rect 483480 319524 483532 319530
rect 483480 319466 483532 319472
rect 482928 319252 482980 319258
rect 482928 319194 482980 319200
rect 483664 319184 483716 319190
rect 483664 319126 483716 319132
rect 478512 317416 478564 317422
rect 478512 317358 478564 317364
rect 479524 317416 479576 317422
rect 479524 317358 479576 317364
rect 478880 301708 478932 301714
rect 478880 301650 478932 301656
rect 478892 298994 478920 301650
rect 478880 298988 478932 298994
rect 478880 298930 478932 298936
rect 478420 291712 478472 291718
rect 478420 291654 478472 291660
rect 476856 287836 476908 287842
rect 476856 287778 476908 287784
rect 476488 286612 476540 286618
rect 476488 286554 476540 286560
rect 475384 274712 475436 274718
rect 475384 274654 475436 274660
rect 479536 273222 479564 317358
rect 482652 313336 482704 313342
rect 482652 313278 482704 313284
rect 482468 310548 482520 310554
rect 482468 310490 482520 310496
rect 482480 307358 482508 310490
rect 482664 307834 482692 313278
rect 483676 310554 483704 319126
rect 483768 319122 483796 322116
rect 484044 321094 484072 322116
rect 484228 322102 484334 322118
rect 484596 321230 484624 322116
rect 484584 321224 484636 321230
rect 484584 321166 484636 321172
rect 484032 321088 484084 321094
rect 484032 321030 484084 321036
rect 484872 319190 484900 322116
rect 485056 322102 485162 322130
rect 485332 322102 485438 322130
rect 485608 322102 485714 322130
rect 484860 319184 484912 319190
rect 484860 319126 484912 319132
rect 483756 319116 483808 319122
rect 483756 319058 483808 319064
rect 484768 319116 484820 319122
rect 484768 319058 484820 319064
rect 484492 319048 484544 319054
rect 484492 318990 484544 318996
rect 483664 310548 483716 310554
rect 483664 310490 483716 310496
rect 482652 307828 482704 307834
rect 482652 307770 482704 307776
rect 481088 307352 481140 307358
rect 481088 307294 481140 307300
rect 482468 307352 482520 307358
rect 482468 307294 482520 307300
rect 481100 301714 481128 307294
rect 484504 303550 484532 318990
rect 484780 303618 484808 319058
rect 485056 313342 485084 322102
rect 485332 319054 485360 322102
rect 485608 319122 485636 322102
rect 485596 319116 485648 319122
rect 485596 319058 485648 319064
rect 485872 319116 485924 319122
rect 485872 319058 485924 319064
rect 485320 319048 485372 319054
rect 485320 318990 485372 318996
rect 485044 313336 485096 313342
rect 485044 313278 485096 313284
rect 484768 303612 484820 303618
rect 484768 303554 484820 303560
rect 484492 303544 484544 303550
rect 484492 303486 484544 303492
rect 485884 303482 485912 319058
rect 485976 316034 486004 322116
rect 486160 322102 486266 322130
rect 486436 322102 486542 322130
rect 486712 322102 486818 322130
rect 486988 322102 487094 322130
rect 485976 316006 486096 316034
rect 486068 305794 486096 316006
rect 486160 305930 486188 322102
rect 486436 319274 486464 322102
rect 486344 319246 486464 319274
rect 486344 316062 486372 319246
rect 486712 319002 486740 322102
rect 486988 319122 487016 322102
rect 487252 319252 487304 319258
rect 487252 319194 487304 319200
rect 486976 319116 487028 319122
rect 486976 319058 487028 319064
rect 486436 318974 486740 319002
rect 486332 316056 486384 316062
rect 486332 315998 486384 316004
rect 486148 305924 486200 305930
rect 486148 305866 486200 305872
rect 486056 305788 486108 305794
rect 486056 305730 486108 305736
rect 485872 303476 485924 303482
rect 485872 303418 485924 303424
rect 481088 301708 481140 301714
rect 481088 301650 481140 301656
rect 486436 278050 486464 318974
rect 486516 316056 486568 316062
rect 486516 315998 486568 316004
rect 486528 305862 486556 315998
rect 486516 305856 486568 305862
rect 486516 305798 486568 305804
rect 486424 278044 486476 278050
rect 486424 277986 486476 277992
rect 479524 273216 479576 273222
rect 479524 273158 479576 273164
rect 473728 269952 473780 269958
rect 473728 269894 473780 269900
rect 487264 269890 487292 319194
rect 487356 316810 487384 322116
rect 487646 322102 487844 322130
rect 487922 322102 488120 322130
rect 487816 319122 487844 322102
rect 487804 319116 487856 319122
rect 487804 319058 487856 319064
rect 487344 316804 487396 316810
rect 487344 316746 487396 316752
rect 488092 286618 488120 322102
rect 488184 316034 488212 322116
rect 488368 322102 488474 322130
rect 488368 319258 488396 322102
rect 488356 319252 488408 319258
rect 488356 319194 488408 319200
rect 488356 319116 488408 319122
rect 488356 319058 488408 319064
rect 488184 316006 488304 316034
rect 488276 304570 488304 316006
rect 488264 304564 488316 304570
rect 488264 304506 488316 304512
rect 488368 293350 488396 319058
rect 488632 319048 488684 319054
rect 488632 318990 488684 318996
rect 488356 293344 488408 293350
rect 488356 293286 488408 293292
rect 488080 286612 488132 286618
rect 488080 286554 488132 286560
rect 488644 273970 488672 318990
rect 488736 318238 488764 322116
rect 488908 319116 488960 319122
rect 488908 319058 488960 319064
rect 488724 318232 488776 318238
rect 488724 318174 488776 318180
rect 488632 273964 488684 273970
rect 488632 273906 488684 273912
rect 488920 272610 488948 319058
rect 489012 305454 489040 322116
rect 489196 322102 489302 322130
rect 489472 322102 489578 322130
rect 489748 322102 489854 322130
rect 490300 322102 490406 322130
rect 489196 319054 489224 322102
rect 489472 319122 489500 322102
rect 489460 319116 489512 319122
rect 489460 319058 489512 319064
rect 489184 319048 489236 319054
rect 489184 318990 489236 318996
rect 489748 316034 489776 322102
rect 490300 319410 490328 322102
rect 489196 316006 489776 316034
rect 490024 319382 490328 319410
rect 489000 305448 489052 305454
rect 489000 305390 489052 305396
rect 489196 284986 489224 316006
rect 489184 284980 489236 284986
rect 489184 284922 489236 284928
rect 490024 278118 490052 319382
rect 490288 318912 490340 318918
rect 490288 318854 490340 318860
rect 490300 307222 490328 318854
rect 490288 307216 490340 307222
rect 490288 307158 490340 307164
rect 490012 278112 490064 278118
rect 490012 278054 490064 278060
rect 488908 272604 488960 272610
rect 488908 272546 488960 272552
rect 487252 269884 487304 269890
rect 487252 269826 487304 269832
rect 473360 268592 473412 268598
rect 473360 268534 473412 268540
rect 490576 268530 490604 322186
rect 490668 279478 490696 322116
rect 490852 322102 490958 322130
rect 491128 322102 491234 322130
rect 490852 286686 490880 322102
rect 491128 318918 491156 322102
rect 491392 319048 491444 319054
rect 491392 318990 491444 318996
rect 491116 318912 491168 318918
rect 491116 318854 491168 318860
rect 490840 286680 490892 286686
rect 490840 286622 490892 286628
rect 490656 279472 490708 279478
rect 490656 279414 490708 279420
rect 491404 274038 491432 318990
rect 491496 316742 491524 322116
rect 491668 319116 491720 319122
rect 491668 319058 491720 319064
rect 491484 316736 491536 316742
rect 491484 316678 491536 316684
rect 491392 274032 491444 274038
rect 491392 273974 491444 273980
rect 491680 271250 491708 319058
rect 491772 315382 491800 322116
rect 491956 322102 492062 322130
rect 492232 322102 492338 322130
rect 492508 322102 492614 322130
rect 492784 322102 492890 322130
rect 491760 315376 491812 315382
rect 491760 315318 491812 315324
rect 491956 314022 491984 322102
rect 492232 319122 492260 322102
rect 492220 319116 492272 319122
rect 492220 319058 492272 319064
rect 492508 319054 492536 322102
rect 492496 319048 492548 319054
rect 492496 318990 492548 318996
rect 491944 314016 491996 314022
rect 491944 313958 491996 313964
rect 492784 272542 492812 322102
rect 493048 319048 493100 319054
rect 493048 318990 493100 318996
rect 493060 311234 493088 318990
rect 493048 311228 493100 311234
rect 493048 311170 493100 311176
rect 493152 275330 493180 322116
rect 493324 319116 493376 319122
rect 493324 319058 493376 319064
rect 493140 275324 493192 275330
rect 493140 275266 493192 275272
rect 492772 272536 492824 272542
rect 492772 272478 492824 272484
rect 491668 271244 491720 271250
rect 491668 271186 491720 271192
rect 493336 271182 493364 319058
rect 493428 280838 493456 322116
rect 493612 322102 493718 322130
rect 493888 322102 493994 322130
rect 493612 319054 493640 322102
rect 493888 319122 493916 322102
rect 494256 321554 494284 322116
rect 494440 322102 494546 322130
rect 494256 321526 494376 321554
rect 494152 319184 494204 319190
rect 494152 319126 494204 319132
rect 493876 319116 493928 319122
rect 493876 319058 493928 319064
rect 493600 319048 493652 319054
rect 493600 318990 493652 318996
rect 494164 282198 494192 319126
rect 494348 319002 494376 321526
rect 494440 319190 494468 322102
rect 494428 319184 494480 319190
rect 494428 319126 494480 319132
rect 494704 319116 494756 319122
rect 494704 319058 494756 319064
rect 494348 318974 494468 319002
rect 494440 309874 494468 318974
rect 494428 309868 494480 309874
rect 494428 309810 494480 309816
rect 494152 282192 494204 282198
rect 494152 282134 494204 282140
rect 493416 280832 493468 280838
rect 493416 280774 493468 280780
rect 494716 276690 494744 319058
rect 494808 308514 494836 322116
rect 494992 322102 495098 322130
rect 495268 322102 495374 322130
rect 494796 308508 494848 308514
rect 494796 308450 494848 308456
rect 494992 283626 495020 322102
rect 495268 319122 495296 322102
rect 495256 319116 495308 319122
rect 495256 319058 495308 319064
rect 495636 318170 495664 322116
rect 495820 322102 495926 322130
rect 495624 318164 495676 318170
rect 495624 318106 495676 318112
rect 495820 299946 495848 322102
rect 496188 318170 496216 322116
rect 496176 318164 496228 318170
rect 496176 318106 496228 318112
rect 496464 318073 496492 322116
rect 496450 318064 496506 318073
rect 496450 317999 496506 318008
rect 495808 299940 495860 299946
rect 495808 299882 495860 299888
rect 494980 283620 495032 283626
rect 494980 283562 495032 283568
rect 494704 276684 494756 276690
rect 494704 276626 494756 276632
rect 493324 271176 493376 271182
rect 493324 271118 493376 271124
rect 496740 269890 496768 322116
rect 497016 316742 497044 322116
rect 497306 322102 497504 322130
rect 497004 316736 497056 316742
rect 497004 316678 497056 316684
rect 497476 314022 497504 322102
rect 497568 316034 497596 322116
rect 497752 322102 497858 322130
rect 498028 322102 498134 322130
rect 498410 322102 498608 322130
rect 497568 316006 497688 316034
rect 497464 314016 497516 314022
rect 497464 313958 497516 313964
rect 497660 309874 497688 316006
rect 497648 309868 497700 309874
rect 497648 309810 497700 309816
rect 497752 273970 497780 322102
rect 498028 284986 498056 322102
rect 498580 316034 498608 322102
rect 498672 319530 498700 322116
rect 498660 319524 498712 319530
rect 498660 319466 498712 319472
rect 498948 316034 498976 322116
rect 499132 322102 499238 322130
rect 499408 322102 499514 322130
rect 499790 322102 499988 322130
rect 498580 316006 498884 316034
rect 498948 316006 499068 316034
rect 498856 308514 498884 316006
rect 498844 308508 498896 308514
rect 498844 308450 498896 308456
rect 498016 284980 498068 284986
rect 498016 284922 498068 284928
rect 499040 275330 499068 316006
rect 499028 275324 499080 275330
rect 499028 275266 499080 275272
rect 497740 273964 497792 273970
rect 497740 273906 497792 273912
rect 499132 271182 499160 322102
rect 499408 274038 499436 322102
rect 499960 319122 499988 322102
rect 499948 319116 500000 319122
rect 499948 319058 500000 319064
rect 500052 316034 500080 322116
rect 500224 319116 500276 319122
rect 500224 319058 500276 319064
rect 500052 316006 500172 316034
rect 500144 305794 500172 316006
rect 500132 305788 500184 305794
rect 500132 305730 500184 305736
rect 500236 276690 500264 319058
rect 500328 316878 500356 322116
rect 500512 322102 500618 322130
rect 500788 322102 500894 322130
rect 501170 322102 501368 322130
rect 500316 316872 500368 316878
rect 500316 316814 500368 316820
rect 500224 276684 500276 276690
rect 500224 276626 500276 276632
rect 499396 274032 499448 274038
rect 499396 273974 499448 273980
rect 500512 271250 500540 322102
rect 500788 272542 500816 322102
rect 501340 319122 501368 322102
rect 501328 319116 501380 319122
rect 501328 319058 501380 319064
rect 501432 316946 501460 322116
rect 501420 316940 501472 316946
rect 501420 316882 501472 316888
rect 501708 316034 501736 322116
rect 501984 319569 502012 322116
rect 502168 322102 502274 322130
rect 502550 322102 502748 322130
rect 501970 319560 502026 319569
rect 501970 319495 502026 319504
rect 502168 319462 502196 322102
rect 502248 320952 502300 320958
rect 502248 320894 502300 320900
rect 502260 319598 502288 320894
rect 502248 319592 502300 319598
rect 502248 319534 502300 319540
rect 502156 319456 502208 319462
rect 502156 319398 502208 319404
rect 501880 319116 501932 319122
rect 501880 319058 501932 319064
rect 501708 316006 501828 316034
rect 501800 278050 501828 316006
rect 501892 315450 501920 319058
rect 502720 316034 502748 322102
rect 502812 319598 502840 322116
rect 502800 319592 502852 319598
rect 502800 319534 502852 319540
rect 503088 316034 503116 322116
rect 503378 322102 503576 322130
rect 502720 316006 503024 316034
rect 503088 316006 503208 316034
rect 501880 315444 501932 315450
rect 501880 315386 501932 315392
rect 502996 315382 503024 316006
rect 502984 315376 503036 315382
rect 502984 315318 503036 315324
rect 503180 313993 503208 316006
rect 503166 313984 503222 313993
rect 503166 313919 503222 313928
rect 503548 311234 503576 322102
rect 503536 311228 503588 311234
rect 503536 311170 503588 311176
rect 503640 279478 503668 322116
rect 503930 322102 505048 322130
rect 503628 279472 503680 279478
rect 503628 279414 503680 279420
rect 501788 278044 501840 278050
rect 501788 277986 501840 277992
rect 500776 272536 500828 272542
rect 500776 272478 500828 272484
rect 500500 271244 500552 271250
rect 500500 271186 500552 271192
rect 499120 271176 499172 271182
rect 499120 271118 499172 271124
rect 505020 269958 505048 322102
rect 506952 307086 506980 322254
rect 507308 321088 507360 321094
rect 507308 321030 507360 321036
rect 507030 320920 507086 320929
rect 507030 320855 507086 320864
rect 506940 307080 506992 307086
rect 506940 307022 506992 307028
rect 507044 304502 507072 320855
rect 507214 320784 507270 320793
rect 507124 320748 507176 320754
rect 507214 320719 507270 320728
rect 507124 320690 507176 320696
rect 507032 304496 507084 304502
rect 507032 304438 507084 304444
rect 507136 286550 507164 320690
rect 507228 288998 507256 320719
rect 507320 289814 507348 321030
rect 507412 292534 507440 322458
rect 507492 321836 507544 321842
rect 507492 321778 507544 321784
rect 507400 292528 507452 292534
rect 507400 292470 507452 292476
rect 507504 292126 507532 321778
rect 507676 321224 507728 321230
rect 507676 321166 507728 321172
rect 507584 320816 507636 320822
rect 507584 320758 507636 320764
rect 507492 292120 507544 292126
rect 507492 292062 507544 292068
rect 507596 291786 507624 320758
rect 507688 297906 507716 321166
rect 507768 320272 507820 320278
rect 507768 320214 507820 320220
rect 507676 297900 507728 297906
rect 507676 297842 507728 297848
rect 507780 297838 507808 320214
rect 509344 319433 509372 322895
rect 509436 322153 509464 324935
rect 509422 322144 509478 322153
rect 509422 322079 509478 322088
rect 509424 322040 509476 322046
rect 509424 321982 509476 321988
rect 509330 319424 509386 319433
rect 509330 319359 509386 319368
rect 509436 319274 509464 321982
rect 509344 319246 509464 319274
rect 509344 300762 509372 319246
rect 509424 319184 509476 319190
rect 509424 319126 509476 319132
rect 509332 300756 509384 300762
rect 509332 300698 509384 300704
rect 507768 297832 507820 297838
rect 507768 297774 507820 297780
rect 509436 294574 509464 319126
rect 509528 303346 509556 357575
rect 509606 344040 509662 344049
rect 509606 343975 509662 343984
rect 509516 303340 509568 303346
rect 509516 303282 509568 303288
rect 509620 303249 509648 343975
rect 509698 335880 509754 335889
rect 509698 335815 509754 335824
rect 509712 331214 509740 335815
rect 509882 333160 509938 333169
rect 509882 333095 509938 333104
rect 509712 331186 509832 331214
rect 509700 326392 509752 326398
rect 509700 326334 509752 326340
rect 509712 319190 509740 326334
rect 509804 321554 509832 331186
rect 509896 322522 509924 333095
rect 510158 328128 510214 328137
rect 510158 328063 510214 328072
rect 509976 326460 510028 326466
rect 509976 326402 510028 326408
rect 509884 322516 509936 322522
rect 509884 322458 509936 322464
rect 509988 322046 510016 326402
rect 509976 322040 510028 322046
rect 509976 321982 510028 321988
rect 509804 321526 510016 321554
rect 509988 321230 510016 321526
rect 509976 321224 510028 321230
rect 509976 321166 510028 321172
rect 509700 319184 509752 319190
rect 509700 319126 509752 319132
rect 509606 303240 509662 303249
rect 509606 303175 509662 303184
rect 510172 300082 510200 328063
rect 510436 324964 510488 324970
rect 510436 324906 510488 324912
rect 510448 319938 510476 324906
rect 510528 323604 510580 323610
rect 510528 323546 510580 323552
rect 510436 319932 510488 319938
rect 510436 319874 510488 319880
rect 510540 319870 510568 323546
rect 510528 319864 510580 319870
rect 510528 319806 510580 319812
rect 510632 300830 510660 359071
rect 510802 355872 510858 355881
rect 510802 355807 510858 355816
rect 510710 353152 510766 353161
rect 510710 353087 510766 353096
rect 510620 300824 510672 300830
rect 510620 300766 510672 300772
rect 510160 300076 510212 300082
rect 510160 300018 510212 300024
rect 510724 295186 510752 353087
rect 510816 303278 510844 355807
rect 510894 346080 510950 346089
rect 510894 346015 510950 346024
rect 510804 303272 510856 303278
rect 510804 303214 510856 303220
rect 510908 303113 510936 346015
rect 510986 342816 511042 342825
rect 510986 342751 511042 342760
rect 511000 306105 511028 342751
rect 511170 340096 511226 340105
rect 511170 340031 511226 340040
rect 511078 337920 511134 337929
rect 511078 337855 511134 337864
rect 511092 320278 511120 337855
rect 511184 321842 511212 340031
rect 511172 321836 511224 321842
rect 511172 321778 511224 321784
rect 511080 320272 511132 320278
rect 511080 320214 511132 320220
rect 511276 320006 511304 576846
rect 511356 423564 511408 423570
rect 511356 423506 511408 423512
rect 511368 388686 511396 423506
rect 511356 388680 511408 388686
rect 511356 388622 511408 388628
rect 513392 387122 513420 600086
rect 519544 590708 519596 590714
rect 519544 590650 519596 590656
rect 515404 563100 515456 563106
rect 515404 563042 515456 563048
rect 513380 387116 513432 387122
rect 513380 387058 513432 387064
rect 512092 386572 512144 386578
rect 512092 386514 512144 386520
rect 512000 386436 512052 386442
rect 512000 386378 512052 386384
rect 512012 374921 512040 386378
rect 512104 377641 512132 386514
rect 512276 386504 512328 386510
rect 512276 386446 512328 386452
rect 512184 385076 512236 385082
rect 512184 385018 512236 385024
rect 512090 377632 512146 377641
rect 512090 377567 512146 377576
rect 512196 376553 512224 385018
rect 512288 378185 512316 386446
rect 513286 384704 513342 384713
rect 513286 384639 513342 384648
rect 512458 384160 512514 384169
rect 512458 384095 512514 384104
rect 512472 383722 512500 384095
rect 513300 383790 513328 384639
rect 513288 383784 513340 383790
rect 513288 383726 513340 383732
rect 512460 383716 512512 383722
rect 512460 383658 512512 383664
rect 512642 383616 512698 383625
rect 512642 383551 512698 383560
rect 512656 383042 512684 383551
rect 513286 383072 513342 383081
rect 512644 383036 512696 383042
rect 513286 383007 513342 383016
rect 512644 382978 512696 382984
rect 513300 382634 513328 383007
rect 513288 382628 513340 382634
rect 513288 382570 513340 382576
rect 512458 382528 512514 382537
rect 512458 382463 512460 382472
rect 512512 382463 512514 382472
rect 512460 382434 512512 382440
rect 513102 381984 513158 381993
rect 513102 381919 513158 381928
rect 512458 381440 512514 381449
rect 512458 381375 512514 381384
rect 512472 380934 512500 381375
rect 512460 380928 512512 380934
rect 512460 380870 512512 380876
rect 512550 379808 512606 379817
rect 512550 379743 512552 379752
rect 512604 379743 512606 379752
rect 512552 379714 512604 379720
rect 512826 379264 512882 379273
rect 512826 379199 512882 379208
rect 512840 378282 512868 379199
rect 512828 378276 512880 378282
rect 512828 378218 512880 378224
rect 512274 378176 512330 378185
rect 512274 378111 512330 378120
rect 512826 377088 512882 377097
rect 512826 377023 512882 377032
rect 512840 376786 512868 377023
rect 512828 376780 512880 376786
rect 512828 376722 512880 376728
rect 512182 376544 512238 376553
rect 512182 376479 512238 376488
rect 513116 376038 513144 381919
rect 513194 380896 513250 380905
rect 513194 380831 513250 380840
rect 513208 377466 513236 380831
rect 513286 380352 513342 380361
rect 513286 380287 513342 380296
rect 513300 379574 513328 380287
rect 513288 379568 513340 379574
rect 513288 379510 513340 379516
rect 513286 378720 513342 378729
rect 513286 378655 513342 378664
rect 513300 378350 513328 378655
rect 513288 378344 513340 378350
rect 513288 378286 513340 378292
rect 514024 378208 514076 378214
rect 514024 378150 514076 378156
rect 513196 377460 513248 377466
rect 513196 377402 513248 377408
rect 513104 376032 513156 376038
rect 513104 375974 513156 375980
rect 513286 376000 513342 376009
rect 513286 375935 513288 375944
rect 513340 375935 513342 375944
rect 513288 375906 513340 375912
rect 513286 375456 513342 375465
rect 513286 375391 513288 375400
rect 513340 375391 513342 375400
rect 513288 375362 513340 375368
rect 511998 374912 512054 374921
rect 511998 374847 512054 374856
rect 512090 374368 512146 374377
rect 512090 374303 512146 374312
rect 512104 374066 512132 374303
rect 512092 374060 512144 374066
rect 512092 374002 512144 374008
rect 511998 373824 512054 373833
rect 511998 373759 512054 373768
rect 512012 372638 512040 373759
rect 512458 373280 512514 373289
rect 512458 373215 512514 373224
rect 512472 372774 512500 373215
rect 512460 372768 512512 372774
rect 512090 372736 512146 372745
rect 512460 372710 512512 372716
rect 512090 372671 512092 372680
rect 512144 372671 512146 372680
rect 512092 372642 512144 372648
rect 512000 372632 512052 372638
rect 512000 372574 512052 372580
rect 512458 372192 512514 372201
rect 512458 372127 512514 372136
rect 512472 371958 512500 372127
rect 512460 371952 512512 371958
rect 512460 371894 512512 371900
rect 512090 371648 512146 371657
rect 512090 371583 512146 371592
rect 511998 367840 512054 367849
rect 511998 367775 512054 367784
rect 512012 367130 512040 367775
rect 512000 367124 512052 367130
rect 512000 367066 512052 367072
rect 511998 366208 512054 366217
rect 511998 366143 512054 366152
rect 512012 365906 512040 366143
rect 512000 365900 512052 365906
rect 512000 365842 512052 365848
rect 511998 362400 512054 362409
rect 511998 362335 512000 362344
rect 512052 362335 512054 362344
rect 512000 362306 512052 362312
rect 511998 354240 512054 354249
rect 511998 354175 512054 354184
rect 512012 354006 512040 354175
rect 512000 354000 512052 354006
rect 512000 353942 512052 353948
rect 511998 352608 512054 352617
rect 511998 352543 512054 352552
rect 512012 352442 512040 352543
rect 512000 352436 512052 352442
rect 512000 352378 512052 352384
rect 511998 350432 512054 350441
rect 511998 350367 512054 350376
rect 512012 349450 512040 350367
rect 512000 349444 512052 349450
rect 512000 349386 512052 349392
rect 511998 349344 512054 349353
rect 511998 349279 512000 349288
rect 512052 349279 512054 349288
rect 512000 349250 512052 349256
rect 511998 339008 512054 339017
rect 511998 338943 512054 338952
rect 511446 335744 511502 335753
rect 511446 335679 511502 335688
rect 511460 322318 511488 335679
rect 511814 327176 511870 327185
rect 511814 327111 511870 327120
rect 511448 322312 511500 322318
rect 511448 322254 511500 322260
rect 511828 320929 511856 327111
rect 511908 323672 511960 323678
rect 511908 323614 511960 323620
rect 511814 320920 511870 320929
rect 511814 320855 511870 320864
rect 511264 320000 511316 320006
rect 511264 319942 511316 319948
rect 511920 319666 511948 323614
rect 511908 319660 511960 319666
rect 511908 319602 511960 319608
rect 510986 306096 511042 306105
rect 510986 306031 511042 306040
rect 510894 303104 510950 303113
rect 510894 303039 510950 303048
rect 510712 295180 510764 295186
rect 510712 295122 510764 295128
rect 509424 294568 509476 294574
rect 509424 294510 509476 294516
rect 507584 291780 507636 291786
rect 507584 291722 507636 291728
rect 507308 289808 507360 289814
rect 507308 289750 507360 289756
rect 507216 288992 507268 288998
rect 507216 288934 507268 288940
rect 507124 286544 507176 286550
rect 507124 286486 507176 286492
rect 505008 269952 505060 269958
rect 505008 269894 505060 269900
rect 496728 269884 496780 269890
rect 496728 269826 496780 269832
rect 490564 268524 490616 268530
rect 490564 268466 490616 268472
rect 466368 268456 466420 268462
rect 466368 268398 466420 268404
rect 512012 268394 512040 338943
rect 512104 305658 512132 371583
rect 512826 371104 512882 371113
rect 512826 371039 512882 371048
rect 512458 370560 512514 370569
rect 512458 370495 512514 370504
rect 512472 370394 512500 370495
rect 512460 370388 512512 370394
rect 512460 370330 512512 370336
rect 512840 369986 512868 371039
rect 513286 370016 513342 370025
rect 512828 369980 512880 369986
rect 513286 369951 513342 369960
rect 512828 369922 512880 369928
rect 513300 369918 513328 369951
rect 513288 369912 513340 369918
rect 513288 369854 513340 369860
rect 513286 369472 513342 369481
rect 513286 369407 513342 369416
rect 512826 368928 512882 368937
rect 512826 368863 512882 368872
rect 512840 368626 512868 368863
rect 512828 368620 512880 368626
rect 512828 368562 512880 368568
rect 513300 368558 513328 369407
rect 513288 368552 513340 368558
rect 513288 368494 513340 368500
rect 512182 368384 512238 368393
rect 512182 368319 512238 368328
rect 512092 305652 512144 305658
rect 512092 305594 512144 305600
rect 512196 304366 512224 368319
rect 513286 367296 513342 367305
rect 513286 367231 513288 367240
rect 513340 367231 513342 367240
rect 513288 367202 513340 367208
rect 513286 366752 513342 366761
rect 513286 366687 513342 366696
rect 513300 365770 513328 366687
rect 513288 365764 513340 365770
rect 513288 365706 513340 365712
rect 512644 365220 512696 365226
rect 512644 365162 512696 365168
rect 512656 364585 512684 365162
rect 513286 365120 513342 365129
rect 513286 365055 513342 365064
rect 512642 364576 512698 364585
rect 512642 364511 512698 364520
rect 513300 364410 513328 365055
rect 513288 364404 513340 364410
rect 513288 364346 513340 364352
rect 513286 363624 513342 363633
rect 513342 363582 513512 363610
rect 513286 363559 513342 363568
rect 512458 363488 512514 363497
rect 512458 363423 512514 363432
rect 512472 363050 512500 363423
rect 512460 363044 512512 363050
rect 512460 362986 512512 362992
rect 513010 362944 513066 362953
rect 513010 362879 513066 362888
rect 512274 361856 512330 361865
rect 512274 361791 512330 361800
rect 512184 304360 512236 304366
rect 512184 304302 512236 304308
rect 512288 300150 512316 361791
rect 513024 361622 513052 362879
rect 513012 361616 513064 361622
rect 513012 361558 513064 361564
rect 513194 361312 513250 361321
rect 513194 361247 513250 361256
rect 512920 361004 512972 361010
rect 512920 360946 512972 360952
rect 512366 360768 512422 360777
rect 512366 360703 512368 360712
rect 512420 360703 512422 360712
rect 512368 360674 512420 360680
rect 512932 360233 512960 360946
rect 513208 360602 513236 361247
rect 513196 360596 513248 360602
rect 513196 360538 513248 360544
rect 512918 360224 512974 360233
rect 512918 360159 512974 360168
rect 512734 359680 512790 359689
rect 512734 359615 512790 359624
rect 512748 358834 512776 359615
rect 512736 358828 512788 358834
rect 512736 358770 512788 358776
rect 512366 358592 512422 358601
rect 512366 358527 512422 358536
rect 512380 302938 512408 358527
rect 513286 358048 513342 358057
rect 513286 357983 513342 357992
rect 513300 357882 513328 357983
rect 513288 357876 513340 357882
rect 513288 357818 513340 357824
rect 513286 356960 513342 356969
rect 513286 356895 513342 356904
rect 513300 356114 513328 356895
rect 513288 356108 513340 356114
rect 513288 356050 513340 356056
rect 512458 355328 512514 355337
rect 512458 355263 512514 355272
rect 512368 302932 512420 302938
rect 512368 302874 512420 302880
rect 512472 301578 512500 355263
rect 513288 355020 513340 355026
rect 513288 354962 513340 354968
rect 513300 354793 513328 354962
rect 513286 354784 513342 354793
rect 513286 354719 513342 354728
rect 513484 354674 513512 363582
rect 513656 362364 513708 362370
rect 513656 362306 513708 362312
rect 513484 354646 513604 354674
rect 513286 353696 513342 353705
rect 513286 353631 513342 353640
rect 513300 353530 513328 353631
rect 513288 353524 513340 353530
rect 513288 353466 513340 353472
rect 513286 352064 513342 352073
rect 513286 351999 513342 352008
rect 513300 351966 513328 351999
rect 513288 351960 513340 351966
rect 513288 351902 513340 351908
rect 512642 351520 512698 351529
rect 512642 351455 512698 351464
rect 512550 350976 512606 350985
rect 512656 350946 512684 351455
rect 512550 350911 512606 350920
rect 512644 350940 512696 350946
rect 512564 350674 512592 350911
rect 512644 350882 512696 350888
rect 512552 350668 512604 350674
rect 512552 350610 512604 350616
rect 513286 349888 513342 349897
rect 513286 349823 513342 349832
rect 513300 349586 513328 349823
rect 513288 349580 513340 349586
rect 513288 349522 513340 349528
rect 513286 348800 513342 348809
rect 513286 348735 513342 348744
rect 512918 348256 512974 348265
rect 512918 348191 512974 348200
rect 512932 348090 512960 348191
rect 512920 348084 512972 348090
rect 512920 348026 512972 348032
rect 513300 347818 513328 348735
rect 513288 347812 513340 347818
rect 513288 347754 513340 347760
rect 512550 347712 512606 347721
rect 512550 347647 512606 347656
rect 512564 346594 512592 347647
rect 513286 347168 513342 347177
rect 513286 347103 513342 347112
rect 513300 347002 513328 347103
rect 513288 346996 513340 347002
rect 513288 346938 513340 346944
rect 513286 346624 513342 346633
rect 512552 346588 512604 346594
rect 513286 346559 513342 346568
rect 512552 346530 512604 346536
rect 513300 346526 513328 346559
rect 513288 346520 513340 346526
rect 513288 346462 513340 346468
rect 512550 345536 512606 345545
rect 512550 345471 512606 345480
rect 512460 301572 512512 301578
rect 512460 301514 512512 301520
rect 512564 301510 512592 345471
rect 513010 344992 513066 345001
rect 513010 344927 513066 344936
rect 512826 343904 512882 343913
rect 513024 343874 513052 344927
rect 512826 343839 512882 343848
rect 513012 343868 513064 343874
rect 512840 343806 512868 343839
rect 513012 343810 513064 343816
rect 512828 343800 512880 343806
rect 512828 343742 512880 343748
rect 513010 343360 513066 343369
rect 513010 343295 513066 343304
rect 513024 342378 513052 343295
rect 513012 342372 513064 342378
rect 513012 342314 513064 342320
rect 512826 342272 512882 342281
rect 512826 342207 512882 342216
rect 512642 340640 512698 340649
rect 512642 340575 512698 340584
rect 512656 339794 512684 340575
rect 512644 339788 512696 339794
rect 512644 339730 512696 339736
rect 512642 339552 512698 339561
rect 512642 339487 512644 339496
rect 512696 339487 512698 339496
rect 512644 339458 512696 339464
rect 512734 334656 512790 334665
rect 512734 334591 512790 334600
rect 512642 331392 512698 331401
rect 512642 331327 512644 331336
rect 512696 331327 512698 331336
rect 512644 331298 512696 331304
rect 512642 329216 512698 329225
rect 512642 329151 512698 329160
rect 512656 328642 512684 329151
rect 512644 328636 512696 328642
rect 512644 328578 512696 328584
rect 512644 320816 512696 320822
rect 512644 320758 512696 320764
rect 512552 301504 512604 301510
rect 512552 301446 512604 301452
rect 512656 300286 512684 320758
rect 512748 304298 512776 334591
rect 512840 320822 512868 342207
rect 513286 341728 513342 341737
rect 513286 341663 513342 341672
rect 513300 341426 513328 341663
rect 513288 341420 513340 341426
rect 513288 341362 513340 341368
rect 513286 341184 513342 341193
rect 513286 341119 513288 341128
rect 513340 341119 513342 341128
rect 513288 341090 513340 341096
rect 513010 338464 513066 338473
rect 513010 338399 513012 338408
rect 513064 338399 513066 338408
rect 513012 338370 513064 338376
rect 513286 337376 513342 337385
rect 513196 337340 513248 337346
rect 513286 337311 513342 337320
rect 513196 337282 513248 337288
rect 513208 336841 513236 337282
rect 513300 337210 513328 337311
rect 513288 337204 513340 337210
rect 513288 337146 513340 337152
rect 513194 336832 513250 336841
rect 513194 336767 513250 336776
rect 513010 335200 513066 335209
rect 513010 335135 513066 335144
rect 513024 334762 513052 335135
rect 513288 334892 513340 334898
rect 513288 334834 513340 334840
rect 513012 334756 513064 334762
rect 513012 334698 513064 334704
rect 513300 334121 513328 334834
rect 513286 334112 513342 334121
rect 513286 334047 513342 334056
rect 513194 331936 513250 331945
rect 513194 331871 513250 331880
rect 513208 331214 513236 331871
rect 513208 331186 513420 331214
rect 512918 327040 512974 327049
rect 512918 326975 512974 326984
rect 512828 320816 512880 320822
rect 512828 320758 512880 320764
rect 512932 316034 512960 326975
rect 513392 320754 513420 331186
rect 513470 330848 513526 330857
rect 513470 330783 513526 330792
rect 513380 320748 513432 320754
rect 513380 320690 513432 320696
rect 513484 320686 513512 330783
rect 513472 320680 513524 320686
rect 513472 320622 513524 320628
rect 512840 316006 512960 316034
rect 512736 304292 512788 304298
rect 512736 304234 512788 304240
rect 512840 302841 512868 316006
rect 512826 302832 512882 302841
rect 512826 302767 512882 302776
rect 513576 300558 513604 354646
rect 513668 300694 513696 362306
rect 513748 354000 513800 354006
rect 513748 353942 513800 353948
rect 513760 303074 513788 353942
rect 513840 349308 513892 349314
rect 513840 349250 513892 349256
rect 513748 303068 513800 303074
rect 513748 303010 513800 303016
rect 513852 302977 513880 349250
rect 513932 331356 513984 331362
rect 513932 331298 513984 331304
rect 513838 302968 513894 302977
rect 513838 302903 513894 302912
rect 513656 300688 513708 300694
rect 513656 300630 513708 300636
rect 513564 300552 513616 300558
rect 513564 300494 513616 300500
rect 512644 300280 512696 300286
rect 512644 300222 512696 300228
rect 512276 300144 512328 300150
rect 512276 300086 512328 300092
rect 513944 297634 513972 331298
rect 514036 321162 514064 378150
rect 514760 372700 514812 372706
rect 514760 372642 514812 372648
rect 514116 367124 514168 367130
rect 514116 367066 514168 367072
rect 514024 321156 514076 321162
rect 514024 321098 514076 321104
rect 513932 297628 513984 297634
rect 513932 297570 513984 297576
rect 514128 292194 514156 367066
rect 514208 365900 514260 365906
rect 514208 365842 514260 365848
rect 514220 295322 514248 365842
rect 514208 295316 514260 295322
rect 514208 295258 514260 295264
rect 514772 292330 514800 372642
rect 514852 372632 514904 372638
rect 514852 372574 514904 372580
rect 514864 300422 514892 372574
rect 515036 360732 515088 360738
rect 515036 360674 515088 360680
rect 514944 349444 514996 349450
rect 514944 349386 514996 349392
rect 514852 300416 514904 300422
rect 514852 300358 514904 300364
rect 514760 292324 514812 292330
rect 514760 292266 514812 292272
rect 514116 292188 514168 292194
rect 514116 292130 514168 292136
rect 514956 289066 514984 349386
rect 515048 300626 515076 360674
rect 515128 352436 515180 352442
rect 515128 352378 515180 352384
rect 515140 303006 515168 352378
rect 515220 350668 515272 350674
rect 515220 350610 515272 350616
rect 515232 303210 515260 350610
rect 515312 346588 515364 346594
rect 515312 346530 515364 346536
rect 515220 303204 515272 303210
rect 515220 303146 515272 303152
rect 515324 303142 515352 346530
rect 515416 322658 515444 563042
rect 518164 484424 518216 484430
rect 518164 484366 518216 484372
rect 515496 470620 515548 470626
rect 515496 470562 515548 470568
rect 515404 322652 515456 322658
rect 515404 322594 515456 322600
rect 515508 322590 515536 470562
rect 515588 382492 515640 382498
rect 515588 382434 515640 382440
rect 515600 358494 515628 382434
rect 515680 379772 515732 379778
rect 515680 379714 515732 379720
rect 515692 359854 515720 379714
rect 516232 376780 516284 376786
rect 516232 376722 516284 376728
rect 515680 359848 515732 359854
rect 515680 359790 515732 359796
rect 515588 358488 515640 358494
rect 515588 358430 515640 358436
rect 516140 339788 516192 339794
rect 516140 339730 516192 339736
rect 515588 339516 515640 339522
rect 515588 339458 515640 339464
rect 515496 322584 515548 322590
rect 515496 322526 515548 322532
rect 515312 303136 515364 303142
rect 515312 303078 515364 303084
rect 515128 303000 515180 303006
rect 515128 302942 515180 302948
rect 515036 300620 515088 300626
rect 515036 300562 515088 300568
rect 515600 297566 515628 339458
rect 516152 321026 516180 339730
rect 516140 321020 516192 321026
rect 516140 320962 516192 320968
rect 516244 305726 516272 376722
rect 516324 371952 516376 371958
rect 516324 371894 516376 371900
rect 516232 305720 516284 305726
rect 516232 305662 516284 305668
rect 516336 300354 516364 371894
rect 517612 370388 517664 370394
rect 517612 370330 517664 370336
rect 516876 369980 516928 369986
rect 516876 369922 516928 369928
rect 516416 368620 516468 368626
rect 516416 368562 516468 368568
rect 516428 300490 516456 368562
rect 516508 348084 516560 348090
rect 516508 348026 516560 348032
rect 516416 300484 516468 300490
rect 516416 300426 516468 300432
rect 516324 300348 516376 300354
rect 516324 300290 516376 300296
rect 515588 297560 515640 297566
rect 515588 297502 515640 297508
rect 516520 294710 516548 348026
rect 516692 343868 516744 343874
rect 516692 343810 516744 343816
rect 516600 338428 516652 338434
rect 516600 338370 516652 338376
rect 516508 294704 516560 294710
rect 516508 294646 516560 294652
rect 516612 291922 516640 338370
rect 516704 297702 516732 343810
rect 516784 342372 516836 342378
rect 516784 342314 516836 342320
rect 516692 297696 516744 297702
rect 516692 297638 516744 297644
rect 516796 297430 516824 342314
rect 516784 297424 516836 297430
rect 516784 297366 516836 297372
rect 516888 292262 516916 369922
rect 517520 343800 517572 343806
rect 517520 343742 517572 343748
rect 516968 328636 517020 328642
rect 516968 328578 517020 328584
rect 516980 320793 517008 328578
rect 517532 321094 517560 343742
rect 517520 321088 517572 321094
rect 517520 321030 517572 321036
rect 516966 320784 517022 320793
rect 516966 320719 517022 320728
rect 517624 300218 517652 370330
rect 517980 367260 518032 367266
rect 517980 367202 518032 367208
rect 517704 360596 517756 360602
rect 517704 360538 517756 360544
rect 517612 300212 517664 300218
rect 517612 300154 517664 300160
rect 517716 295118 517744 360538
rect 517888 358828 517940 358834
rect 517888 358770 517940 358776
rect 517796 353524 517848 353530
rect 517796 353466 517848 353472
rect 517704 295112 517756 295118
rect 517704 295054 517756 295060
rect 516876 292256 516928 292262
rect 516876 292198 516928 292204
rect 516600 291916 516652 291922
rect 516600 291858 516652 291864
rect 517808 289678 517836 353466
rect 517900 295050 517928 358770
rect 517992 305697 518020 367202
rect 518072 346520 518124 346526
rect 518072 346462 518124 346468
rect 517978 305688 518034 305697
rect 517978 305623 518034 305632
rect 518084 297770 518112 346462
rect 518176 319734 518204 484366
rect 518256 382628 518308 382634
rect 518256 382570 518308 382576
rect 518268 358698 518296 382570
rect 518900 375964 518952 375970
rect 518900 375906 518952 375912
rect 518348 375420 518400 375426
rect 518348 375362 518400 375368
rect 518256 358692 518308 358698
rect 518256 358634 518308 358640
rect 518256 341148 518308 341154
rect 518256 341090 518308 341096
rect 518164 319728 518216 319734
rect 518164 319670 518216 319676
rect 518268 297974 518296 341090
rect 518256 297968 518308 297974
rect 518256 297910 518308 297916
rect 518072 297764 518124 297770
rect 518072 297706 518124 297712
rect 518360 297498 518388 375362
rect 518348 297492 518400 297498
rect 518348 297434 518400 297440
rect 517888 295044 517940 295050
rect 517888 294986 517940 294992
rect 518912 292398 518940 375906
rect 518992 361004 519044 361010
rect 518992 360946 519044 360952
rect 518900 292392 518952 292398
rect 518900 292334 518952 292340
rect 519004 289746 519032 360946
rect 519084 357876 519136 357882
rect 519084 357818 519136 357824
rect 519096 294914 519124 357818
rect 519176 355020 519228 355026
rect 519176 354962 519228 354968
rect 519084 294908 519136 294914
rect 519084 294850 519136 294856
rect 519188 294846 519216 354962
rect 519360 350940 519412 350946
rect 519360 350882 519412 350888
rect 519268 346996 519320 347002
rect 519268 346938 519320 346944
rect 519176 294840 519228 294846
rect 519176 294782 519228 294788
rect 518992 289740 519044 289746
rect 518992 289682 519044 289688
rect 517796 289672 517848 289678
rect 517796 289614 517848 289620
rect 519280 289474 519308 346938
rect 519372 294778 519400 350882
rect 519452 349580 519504 349586
rect 519452 349522 519504 349528
rect 519360 294772 519412 294778
rect 519360 294714 519412 294720
rect 519464 294642 519492 349522
rect 519556 319802 519584 590650
rect 520292 520946 520320 600086
rect 526732 598262 526760 600100
rect 526720 598256 526772 598262
rect 526720 598198 526772 598204
rect 520280 520940 520332 520946
rect 520280 520882 520332 520888
rect 547878 516760 547934 516769
rect 547878 516695 547934 516704
rect 545120 514072 545172 514078
rect 545120 514014 545172 514020
rect 535460 512644 535512 512650
rect 535460 512586 535512 512592
rect 519636 510672 519688 510678
rect 519636 510614 519688 510620
rect 519648 322726 519676 510614
rect 532700 508564 532752 508570
rect 532700 508506 532752 508512
rect 529940 505776 529992 505782
rect 529940 505718 529992 505724
rect 529952 480254 529980 505718
rect 532712 480254 532740 508506
rect 535472 480254 535500 512586
rect 538220 509924 538272 509930
rect 538220 509866 538272 509872
rect 538232 480254 538260 509866
rect 529952 480226 530256 480254
rect 532712 480226 533200 480254
rect 535472 480226 536144 480254
rect 538232 480226 539088 480254
rect 521750 462904 521806 462913
rect 521750 462839 521806 462848
rect 521764 460972 521792 462839
rect 527640 462460 527692 462466
rect 527640 462402 527692 462408
rect 524696 461100 524748 461106
rect 524696 461042 524748 461048
rect 524708 460972 524736 461042
rect 527652 460972 527680 462402
rect 530228 460986 530256 480226
rect 533172 460986 533200 480226
rect 536116 460986 536144 480226
rect 539060 460986 539088 480226
rect 542360 462392 542412 462398
rect 542360 462334 542412 462340
rect 530228 460958 530610 460986
rect 533172 460958 533554 460986
rect 536116 460958 536498 460986
rect 539060 460958 539442 460986
rect 542372 460972 542400 462334
rect 545132 460986 545160 514014
rect 547892 460986 547920 516695
rect 553860 461032 553912 461038
rect 545132 460958 545330 460986
rect 547892 460958 548274 460986
rect 550928 460970 551218 460986
rect 553912 460980 554162 460986
rect 553860 460974 554162 460980
rect 550916 460964 551218 460970
rect 550968 460958 551218 460964
rect 553872 460958 554162 460974
rect 550916 460906 550968 460912
rect 569224 456816 569276 456822
rect 569224 456758 569276 456764
rect 557538 442912 557594 442921
rect 557538 442847 557594 442856
rect 521212 421598 521240 425068
rect 522304 423496 522356 423502
rect 522304 423438 522356 423444
rect 521200 421592 521252 421598
rect 521200 421534 521252 421540
rect 522316 388822 522344 423438
rect 522500 423434 522528 425068
rect 523788 423570 523816 425068
rect 524708 425054 525090 425082
rect 523776 423564 523828 423570
rect 523776 423506 523828 423512
rect 522488 423428 522540 423434
rect 522488 423370 522540 423376
rect 523684 423428 523736 423434
rect 523684 423370 523736 423376
rect 522304 388816 522356 388822
rect 522304 388758 522356 388764
rect 523696 388754 523724 423370
rect 524708 412634 524736 425054
rect 526364 423366 526392 425068
rect 526352 423360 526404 423366
rect 526352 423302 526404 423308
rect 526444 423360 526496 423366
rect 526444 423302 526496 423308
rect 524432 412606 524736 412634
rect 523684 388748 523736 388754
rect 523684 388690 523736 388696
rect 524432 388618 524460 412606
rect 526456 388890 526484 423302
rect 527652 416090 527680 425068
rect 528940 423298 528968 425068
rect 530228 423638 530256 425068
rect 529204 423632 529256 423638
rect 529204 423574 529256 423580
rect 530216 423632 530268 423638
rect 530216 423574 530268 423580
rect 530584 423632 530636 423638
rect 530584 423574 530636 423580
rect 528928 423292 528980 423298
rect 528928 423234 528980 423240
rect 527640 416084 527692 416090
rect 527640 416026 527692 416032
rect 526444 388884 526496 388890
rect 526444 388826 526496 388832
rect 524420 388612 524472 388618
rect 524420 388554 524472 388560
rect 529216 388482 529244 423574
rect 530596 388550 530624 423574
rect 531516 423230 531544 425068
rect 532804 423638 532832 425068
rect 532792 423632 532844 423638
rect 532792 423574 532844 423580
rect 531504 423224 531556 423230
rect 531504 423166 531556 423172
rect 534092 389842 534120 425068
rect 535012 425054 535394 425082
rect 536300 425054 536682 425082
rect 537588 425054 537970 425082
rect 538876 425054 539258 425082
rect 540164 425054 540546 425082
rect 535012 412634 535040 425054
rect 536300 412634 536328 425054
rect 537588 412634 537616 425054
rect 538876 412634 538904 425054
rect 540164 412634 540192 425054
rect 541820 420238 541848 425068
rect 542740 425054 543122 425082
rect 544028 425054 544410 425082
rect 541808 420232 541860 420238
rect 541808 420174 541860 420180
rect 542740 412634 542768 425054
rect 544028 412634 544056 425054
rect 545684 423162 545712 425068
rect 546604 425054 546986 425082
rect 545672 423156 545724 423162
rect 545672 423098 545724 423104
rect 546604 412634 546632 425054
rect 548260 423094 548288 425068
rect 549548 423502 549576 425068
rect 549536 423496 549588 423502
rect 549536 423438 549588 423444
rect 548248 423088 548300 423094
rect 548248 423030 548300 423036
rect 550836 423026 550864 425068
rect 552124 423434 552152 425068
rect 552112 423428 552164 423434
rect 552112 423370 552164 423376
rect 550824 423020 550876 423026
rect 550824 422962 550876 422968
rect 553412 422958 553440 425068
rect 554700 423366 554728 425068
rect 554688 423360 554740 423366
rect 554688 423302 554740 423308
rect 553400 422952 553452 422958
rect 553400 422894 553452 422900
rect 534184 412606 535040 412634
rect 535472 412606 536328 412634
rect 536852 412606 537616 412634
rect 538232 412606 538904 412634
rect 539612 412606 540192 412634
rect 542372 412606 542768 412634
rect 543752 412606 544056 412634
rect 546512 412606 546632 412634
rect 534184 392630 534212 412606
rect 535472 395350 535500 412606
rect 536852 396778 536880 412606
rect 538232 398138 538260 412606
rect 539612 399498 539640 412606
rect 539600 399492 539652 399498
rect 539600 399434 539652 399440
rect 538220 398132 538272 398138
rect 538220 398074 538272 398080
rect 536840 396772 536892 396778
rect 536840 396714 536892 396720
rect 535460 395344 535512 395350
rect 535460 395286 535512 395292
rect 534172 392624 534224 392630
rect 534172 392566 534224 392572
rect 542372 391338 542400 412606
rect 543752 394058 543780 412606
rect 546512 400926 546540 412606
rect 557552 402286 557580 442847
rect 557540 402280 557592 402286
rect 557540 402222 557592 402228
rect 546500 400920 546552 400926
rect 546500 400862 546552 400868
rect 543740 394052 543792 394058
rect 543740 393994 543792 394000
rect 542360 391332 542412 391338
rect 542360 391274 542412 391280
rect 534080 389836 534132 389842
rect 534080 389778 534132 389784
rect 530584 388544 530636 388550
rect 530584 388486 530636 388492
rect 529204 388476 529256 388482
rect 529204 388418 529256 388424
rect 553952 386640 554004 386646
rect 553952 386582 554004 386588
rect 530584 383784 530636 383790
rect 530584 383726 530636 383732
rect 519728 383036 519780 383042
rect 519728 382978 519780 382984
rect 519740 358630 519768 382978
rect 522304 378344 522356 378350
rect 522304 378286 522356 378292
rect 520280 374060 520332 374066
rect 520280 374002 520332 374008
rect 519728 358624 519780 358630
rect 519728 358566 519780 358572
rect 519728 337340 519780 337346
rect 519728 337282 519780 337288
rect 519636 322720 519688 322726
rect 519636 322662 519688 322668
rect 519544 319796 519596 319802
rect 519544 319738 519596 319744
rect 519452 294636 519504 294642
rect 519452 294578 519504 294584
rect 519740 291854 519768 337282
rect 520292 292058 520320 374002
rect 521660 372768 521712 372774
rect 521660 372710 521712 372716
rect 520372 368552 520424 368558
rect 520372 368494 520424 368500
rect 520280 292052 520332 292058
rect 520280 291994 520332 292000
rect 520384 291990 520412 368494
rect 520464 365220 520516 365226
rect 520464 365162 520516 365168
rect 520476 294982 520504 365162
rect 520556 361616 520608 361622
rect 520556 361558 520608 361564
rect 520568 295254 520596 361558
rect 520648 341420 520700 341426
rect 520648 341362 520700 341368
rect 520556 295248 520608 295254
rect 520556 295190 520608 295196
rect 520464 294976 520516 294982
rect 520464 294918 520516 294924
rect 520372 291984 520424 291990
rect 520372 291926 520424 291932
rect 519728 291848 519780 291854
rect 519728 291790 519780 291796
rect 519268 289468 519320 289474
rect 519268 289410 519320 289416
rect 520660 289134 520688 341362
rect 520924 337204 520976 337210
rect 520924 337146 520976 337152
rect 520740 334892 520792 334898
rect 520740 334834 520792 334840
rect 520648 289128 520700 289134
rect 520648 289070 520700 289076
rect 514944 289060 514996 289066
rect 514944 289002 514996 289008
rect 520752 286482 520780 334834
rect 520832 334756 520884 334762
rect 520832 334698 520884 334704
rect 520844 292466 520872 334698
rect 520936 304434 520964 337146
rect 520924 304428 520976 304434
rect 520924 304370 520976 304376
rect 520832 292460 520884 292466
rect 520832 292402 520884 292408
rect 520740 286476 520792 286482
rect 520740 286418 520792 286424
rect 521672 286414 521700 372710
rect 521752 365764 521804 365770
rect 521752 365706 521804 365712
rect 521764 289202 521792 365706
rect 521844 363044 521896 363050
rect 521844 362986 521896 362992
rect 521856 289610 521884 362986
rect 522316 360058 522344 378286
rect 523040 369912 523092 369918
rect 523040 369854 523092 369860
rect 522304 360052 522356 360058
rect 522304 359994 522356 360000
rect 521936 351960 521988 351966
rect 521936 351902 521988 351908
rect 521844 289604 521896 289610
rect 521844 289546 521896 289552
rect 521948 289270 521976 351902
rect 521936 289264 521988 289270
rect 521936 289206 521988 289212
rect 521752 289196 521804 289202
rect 521752 289138 521804 289144
rect 521660 286408 521712 286414
rect 521660 286350 521712 286356
rect 523052 286346 523080 369854
rect 523132 364404 523184 364410
rect 523132 364346 523184 364352
rect 523144 289338 523172 364346
rect 530596 360126 530624 383726
rect 548524 383716 548576 383722
rect 548524 383658 548576 383664
rect 547144 380928 547196 380934
rect 547144 380870 547196 380876
rect 544384 376032 544436 376038
rect 544384 375974 544436 375980
rect 530584 360120 530636 360126
rect 530584 360062 530636 360068
rect 544396 358562 544424 375974
rect 547156 359922 547184 380870
rect 547236 378276 547288 378282
rect 547236 378218 547288 378224
rect 547248 360194 547276 378218
rect 547236 360188 547288 360194
rect 547236 360130 547288 360136
rect 547144 359916 547196 359922
rect 547144 359858 547196 359864
rect 548536 359786 548564 383658
rect 549904 379568 549956 379574
rect 549904 379510 549956 379516
rect 548616 377460 548668 377466
rect 548616 377402 548668 377408
rect 548524 359780 548576 359786
rect 548524 359722 548576 359728
rect 548628 358766 548656 377402
rect 549916 359990 549944 379510
rect 553964 377890 553992 386582
rect 563428 385144 563480 385150
rect 563428 385086 563480 385092
rect 553964 377862 554438 377890
rect 563440 377876 563468 385086
rect 552032 360194 552322 360210
rect 552020 360188 552322 360194
rect 552072 360182 552322 360188
rect 552020 360130 552072 360136
rect 566740 360120 566792 360126
rect 550652 360058 550850 360074
rect 550640 360052 550850 360058
rect 550692 360046 550850 360052
rect 550640 359994 550692 360000
rect 549904 359984 549956 359990
rect 549904 359926 549956 359932
rect 553780 359854 553808 360060
rect 554976 360046 555266 360074
rect 554976 359990 555004 360046
rect 554964 359984 555016 359990
rect 554964 359926 555016 359932
rect 553768 359848 553820 359854
rect 553768 359790 553820 359796
rect 556724 358766 556752 360060
rect 558196 359922 558224 360060
rect 558184 359916 558236 359922
rect 558184 359858 558236 359864
rect 548616 358760 548668 358766
rect 548616 358702 548668 358708
rect 556712 358760 556764 358766
rect 556712 358702 556764 358708
rect 559668 358562 559696 360060
rect 544384 358556 544436 358562
rect 544384 358498 544436 358504
rect 559656 358556 559708 358562
rect 559656 358498 559708 358504
rect 561140 358494 561168 360060
rect 562612 358698 562640 360060
rect 562600 358692 562652 358698
rect 562600 358634 562652 358640
rect 564084 358630 564112 360060
rect 565280 360046 565570 360074
rect 566792 360068 567042 360074
rect 566740 360062 567042 360068
rect 566752 360046 567042 360062
rect 565280 359990 565308 360046
rect 565268 359984 565320 359990
rect 565268 359926 565320 359932
rect 564072 358624 564124 358630
rect 564072 358566 564124 358572
rect 561128 358488 561180 358494
rect 561128 358430 561180 358436
rect 523224 356108 523276 356114
rect 523224 356050 523276 356056
rect 523236 289542 523264 356050
rect 523316 347812 523368 347818
rect 523316 347754 523368 347760
rect 523224 289536 523276 289542
rect 523224 289478 523276 289484
rect 523328 289406 523356 347754
rect 569236 322862 569264 456758
rect 570616 322930 570644 616830
rect 570604 322924 570656 322930
rect 570604 322866 570656 322872
rect 569224 322856 569276 322862
rect 569224 322798 569276 322804
rect 571996 322794 572024 643078
rect 574744 630692 574796 630698
rect 574744 630634 574796 630640
rect 573364 430636 573416 430642
rect 573364 430578 573416 430584
rect 571984 322788 572036 322794
rect 571984 322730 572036 322736
rect 573376 321298 573404 430578
rect 574756 321366 574784 630634
rect 574744 321360 574796 321366
rect 574744 321302 574796 321308
rect 573364 321292 573416 321298
rect 573364 321234 573416 321240
rect 576136 320074 576164 696934
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579618 591016 579674 591025
rect 579618 590951 579674 590960
rect 579632 590714 579660 590951
rect 579620 590708 579672 590714
rect 579620 590650 579672 590656
rect 579618 577688 579674 577697
rect 579618 577623 579674 577632
rect 579632 576910 579660 577623
rect 579620 576904 579672 576910
rect 579620 576846 579672 576852
rect 579894 564360 579950 564369
rect 579894 564295 579950 564304
rect 579908 563106 579936 564295
rect 579896 563100 579948 563106
rect 579896 563042 579948 563048
rect 579618 511320 579674 511329
rect 579618 511255 579674 511264
rect 579632 510678 579660 511255
rect 579620 510672 579672 510678
rect 579620 510614 579672 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 579618 431624 579674 431633
rect 579618 431559 579674 431568
rect 579632 430642 579660 431559
rect 579620 430636 579672 430642
rect 579620 430578 579672 430584
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 576216 364404 576268 364410
rect 576216 364346 576268 364352
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 576228 321434 576256 364346
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 323678 580212 325207
rect 580172 323672 580224 323678
rect 580172 323614 580224 323620
rect 576216 321428 576268 321434
rect 576216 321370 576268 321376
rect 580276 320958 580304 683839
rect 580354 670712 580410 670721
rect 580354 670647 580410 670656
rect 580264 320952 580316 320958
rect 580264 320894 580316 320900
rect 580368 320890 580396 670647
rect 580446 537840 580502 537849
rect 580446 537775 580502 537784
rect 580356 320884 580408 320890
rect 580356 320826 580408 320832
rect 580460 320142 580488 537775
rect 580538 524512 580594 524521
rect 580538 524447 580594 524456
rect 580552 323610 580580 524447
rect 580630 418296 580686 418305
rect 580630 418231 580686 418240
rect 580644 324970 580672 418231
rect 580722 404968 580778 404977
rect 580722 404903 580778 404912
rect 580632 324964 580684 324970
rect 580632 324906 580684 324912
rect 580540 323604 580592 323610
rect 580540 323546 580592 323552
rect 580736 321502 580764 404903
rect 580814 351928 580870 351937
rect 580814 351863 580870 351872
rect 580828 321570 580856 351863
rect 580816 321564 580868 321570
rect 580816 321506 580868 321512
rect 580724 321496 580776 321502
rect 580724 321438 580776 321444
rect 580448 320136 580500 320142
rect 580448 320078 580500 320084
rect 576124 320068 576176 320074
rect 576124 320010 576176 320016
rect 533344 319592 533396 319598
rect 533344 319534 533396 319540
rect 529940 316804 529992 316810
rect 529940 316746 529992 316752
rect 523316 289400 523368 289406
rect 523316 289342 523368 289348
rect 523132 289332 523184 289338
rect 523132 289274 523184 289280
rect 523040 286340 523092 286346
rect 523040 286282 523092 286288
rect 512000 268388 512052 268394
rect 512000 268330 512052 268336
rect 529952 209273 529980 316746
rect 531412 304564 531464 304570
rect 531412 304506 531464 304512
rect 530032 293344 530084 293350
rect 530032 293286 530084 293292
rect 530044 226250 530072 293286
rect 531320 286612 531372 286618
rect 531320 286554 531372 286560
rect 531332 243681 531360 286554
rect 531424 261089 531452 304506
rect 531410 261080 531466 261089
rect 531410 261015 531466 261024
rect 531318 243672 531374 243681
rect 531318 243607 531374 243616
rect 530122 226264 530178 226273
rect 530044 226222 530122 226250
rect 530122 226199 530178 226208
rect 529938 209264 529994 209273
rect 529938 209199 529994 209208
rect 462320 200728 462372 200734
rect 462320 200670 462372 200676
rect 460768 200110 460980 200138
rect 460388 161492 460440 161498
rect 460388 161434 460440 161440
rect 460400 143546 460428 161434
rect 460388 143540 460440 143546
rect 460388 143482 460440 143488
rect 460848 143540 460900 143546
rect 460848 143482 460900 143488
rect 460860 142322 460888 143482
rect 460848 142316 460900 142322
rect 460848 142258 460900 142264
rect 460860 67697 460888 142258
rect 460386 67688 460442 67697
rect 460386 67623 460442 67632
rect 460846 67688 460902 67697
rect 460846 67623 460902 67632
rect 460296 31748 460348 31754
rect 460296 31690 460348 31696
rect 460400 31686 460428 67623
rect 460388 31680 460440 31686
rect 460388 31622 460440 31628
rect 460952 28490 460980 200110
rect 461584 199436 461636 199442
rect 461584 199378 461636 199384
rect 461596 41410 461624 199378
rect 461584 41404 461636 41410
rect 461584 41346 461636 41352
rect 460940 28484 460992 28490
rect 460940 28426 460992 28432
rect 462332 28286 462360 200670
rect 528560 182844 528612 182850
rect 528560 182786 528612 182792
rect 524420 171828 524472 171834
rect 524420 171770 524472 171776
rect 489920 162240 489972 162246
rect 489920 162182 489972 162188
rect 485780 162172 485832 162178
rect 485780 162114 485832 162120
rect 481916 142316 481968 142322
rect 481916 142258 481968 142264
rect 481928 139890 481956 142258
rect 485792 139890 485820 162114
rect 489932 139890 489960 162182
rect 521660 160744 521712 160750
rect 521660 160686 521712 160692
rect 496820 160472 496872 160478
rect 496820 160414 496872 160420
rect 494060 160336 494112 160342
rect 494060 160278 494112 160284
rect 494072 139890 494100 160278
rect 496832 151814 496860 160414
rect 500960 160404 501012 160410
rect 500960 160346 501012 160352
rect 500972 151814 501000 160346
rect 509240 160268 509292 160274
rect 509240 160210 509292 160216
rect 509252 151814 509280 160210
rect 513380 160200 513432 160206
rect 513380 160142 513432 160148
rect 513392 151814 513420 160142
rect 517520 160132 517572 160138
rect 517520 160074 517572 160080
rect 496832 151786 497688 151814
rect 500972 151786 501644 151814
rect 509252 151786 509556 151814
rect 513392 151786 513512 151814
rect 497660 139890 497688 151786
rect 501616 139890 501644 151786
rect 505652 142248 505704 142254
rect 505652 142190 505704 142196
rect 505664 139890 505692 142190
rect 509528 139890 509556 151786
rect 513484 139890 513512 151786
rect 517532 139890 517560 160074
rect 521672 139890 521700 160686
rect 524432 151814 524460 171770
rect 528572 151814 528600 182786
rect 524432 151786 525380 151814
rect 528572 151786 529336 151814
rect 525352 139890 525380 151786
rect 529308 139890 529336 151786
rect 533356 140078 533384 319534
rect 534724 319524 534776 319530
rect 534724 319466 534776 319472
rect 533436 309800 533488 309806
rect 533436 309742 533488 309748
rect 533448 143546 533476 309742
rect 533436 143540 533488 143546
rect 533436 143482 533488 143488
rect 533988 142180 534040 142186
rect 533988 142122 534040 142128
rect 533344 140072 533396 140078
rect 533344 140014 533396 140020
rect 534000 139890 534028 142122
rect 534736 140146 534764 319466
rect 538864 319456 538916 319462
rect 538864 319398 538916 319404
rect 536104 308440 536156 308446
rect 536104 308382 536156 308388
rect 536116 167006 536144 308382
rect 536104 167000 536156 167006
rect 536104 166942 536156 166948
rect 537300 143540 537352 143546
rect 537300 143482 537352 143488
rect 534724 140140 534776 140146
rect 534724 140082 534776 140088
rect 481928 139862 482264 139890
rect 485792 139862 486220 139890
rect 489932 139862 490176 139890
rect 494072 139862 494132 139890
rect 497660 139862 498088 139890
rect 501616 139862 502044 139890
rect 505664 139862 506000 139890
rect 509528 139862 509956 139890
rect 513484 139862 513912 139890
rect 517532 139862 517868 139890
rect 521672 139862 521824 139890
rect 525352 139862 525780 139890
rect 529308 139862 529736 139890
rect 533692 139862 534028 139890
rect 537312 139890 537340 143482
rect 537312 139862 537648 139890
rect 538876 138650 538904 319398
rect 540980 318164 541032 318170
rect 540980 318106 541032 318112
rect 539692 316940 539744 316946
rect 539692 316882 539744 316888
rect 539600 316872 539652 316878
rect 539600 316814 539652 316820
rect 538956 311228 539008 311234
rect 538956 311170 539008 311176
rect 538864 138644 538916 138650
rect 538864 138586 538916 138592
rect 538968 136610 538996 311170
rect 539048 279472 539100 279478
rect 539048 279414 539100 279420
rect 539060 151814 539088 279414
rect 539060 151786 539364 151814
rect 539336 137737 539364 151786
rect 539322 137728 539378 137737
rect 539322 137663 539378 137672
rect 538956 136604 539008 136610
rect 538956 136546 539008 136552
rect 539508 136604 539560 136610
rect 539508 136546 539560 136552
rect 539520 135969 539548 136546
rect 539506 135960 539562 135969
rect 539506 135895 539562 135904
rect 539612 113257 539640 316814
rect 539704 121417 539732 316882
rect 539784 315444 539836 315450
rect 539784 315386 539836 315392
rect 539690 121408 539746 121417
rect 539690 121343 539746 121352
rect 539796 119649 539824 315386
rect 539876 284980 539928 284986
rect 539876 284922 539928 284928
rect 539782 119640 539838 119649
rect 539782 119575 539838 119584
rect 539598 113248 539654 113257
rect 539598 113183 539654 113192
rect 539888 97209 539916 284922
rect 540244 278044 540296 278050
rect 540244 277986 540296 277992
rect 539968 276684 540020 276690
rect 539968 276626 540020 276632
rect 539980 108769 540008 276626
rect 540152 271244 540204 271250
rect 540152 271186 540204 271192
rect 540060 271176 540112 271182
rect 540060 271118 540112 271124
rect 539966 108760 540022 108769
rect 539966 108695 540022 108704
rect 540072 104689 540100 271118
rect 540164 115025 540192 271186
rect 540256 123185 540284 277986
rect 540336 142248 540388 142254
rect 540336 142190 540388 142196
rect 540242 123176 540298 123185
rect 540242 123111 540298 123120
rect 540150 115016 540206 115025
rect 540150 114951 540206 114960
rect 540058 104680 540114 104689
rect 540058 104615 540114 104624
rect 539874 97200 539930 97209
rect 539874 97135 539930 97144
rect 536840 41404 536892 41410
rect 536840 41346 536892 41352
rect 536852 41041 536880 41346
rect 536838 41032 536894 41041
rect 536838 40967 536894 40976
rect 540348 34241 540376 142190
rect 540992 82385 541020 318106
rect 547144 318096 547196 318102
rect 547144 318038 547196 318044
rect 543004 316736 543056 316742
rect 543004 316678 543056 316684
rect 542728 315376 542780 315382
rect 542728 315318 542780 315324
rect 542452 314016 542504 314022
rect 542452 313958 542504 313964
rect 541072 305788 541124 305794
rect 541072 305730 541124 305736
rect 541084 110945 541112 305730
rect 541256 275324 541308 275330
rect 541256 275266 541308 275272
rect 541164 269884 541216 269890
rect 541164 269826 541216 269832
rect 541070 110936 541126 110945
rect 541070 110871 541126 110880
rect 541176 86465 541204 269826
rect 541268 102785 541296 275266
rect 541348 274032 541400 274038
rect 541348 273974 541400 273980
rect 541360 106865 541388 273974
rect 541440 272536 541492 272542
rect 541440 272478 541492 272484
rect 541452 117065 541480 272478
rect 541438 117056 541494 117065
rect 541438 116991 541494 117000
rect 541346 106856 541402 106865
rect 541346 106791 541402 106800
rect 541254 102776 541310 102785
rect 541254 102711 541310 102720
rect 542464 90545 542492 313958
rect 542544 309868 542596 309874
rect 542544 309810 542596 309816
rect 542556 92585 542584 309810
rect 542636 308508 542688 308514
rect 542636 308450 542688 308456
rect 542648 98705 542676 308450
rect 542740 129305 542768 315318
rect 542820 273964 542872 273970
rect 542820 273906 542872 273912
rect 542726 129296 542782 129305
rect 542726 129231 542782 129240
rect 542634 98696 542690 98705
rect 542634 98631 542690 98640
rect 542832 94625 542860 273906
rect 542912 140140 542964 140146
rect 542912 140082 542964 140088
rect 542924 100745 542952 140082
rect 542910 100736 542966 100745
rect 542910 100671 542966 100680
rect 542818 94616 542874 94625
rect 542818 94551 542874 94560
rect 542542 92576 542598 92585
rect 542542 92511 542598 92520
rect 542450 90536 542506 90545
rect 542450 90471 542506 90480
rect 543016 88505 543044 316678
rect 544384 307148 544436 307154
rect 544384 307090 544436 307096
rect 543740 269952 543792 269958
rect 543740 269894 543792 269900
rect 543188 140072 543240 140078
rect 543188 140014 543240 140020
rect 543096 138644 543148 138650
rect 543096 138586 543148 138592
rect 543108 127265 543136 138586
rect 543200 131345 543228 140014
rect 543278 137864 543334 137873
rect 543278 137799 543334 137808
rect 543186 131336 543242 131345
rect 543186 131271 543242 131280
rect 543094 127256 543150 127265
rect 543094 127191 543150 127200
rect 543292 125225 543320 137799
rect 543278 125216 543334 125225
rect 543278 125151 543334 125160
rect 543002 88496 543058 88505
rect 543002 88431 543058 88440
rect 541162 86456 541218 86465
rect 541162 86391 541218 86400
rect 540978 82376 541034 82385
rect 540978 82311 541034 82320
rect 543752 51134 543780 269894
rect 544396 73166 544424 307090
rect 547156 153202 547184 318038
rect 562324 315308 562376 315314
rect 562324 315250 562376 315256
rect 551284 312588 551336 312594
rect 551284 312530 551336 312536
rect 548524 311160 548576 311166
rect 548524 311102 548576 311108
rect 548536 193186 548564 311102
rect 548524 193180 548576 193186
rect 548524 193122 548576 193128
rect 547144 153196 547196 153202
rect 547144 153138 547196 153144
rect 544384 73160 544436 73166
rect 544384 73102 544436 73108
rect 551296 60722 551324 312530
rect 559564 293276 559616 293282
rect 559564 293218 559616 293224
rect 558184 290488 558236 290494
rect 558184 290430 558236 290436
rect 555424 288924 555476 288930
rect 555424 288866 555476 288872
rect 555436 139398 555464 288866
rect 555424 139392 555476 139398
rect 555424 139334 555476 139340
rect 558196 100706 558224 290430
rect 559576 179382 559604 293218
rect 559656 291712 559708 291718
rect 559656 291654 559708 291660
rect 559668 233238 559696 291654
rect 559656 233232 559708 233238
rect 559656 233174 559708 233180
rect 559564 179376 559616 179382
rect 559564 179318 559616 179324
rect 558184 100700 558236 100706
rect 558184 100642 558236 100648
rect 551284 60716 551336 60722
rect 551284 60658 551336 60664
rect 540612 51128 540664 51134
rect 540612 51070 540664 51076
rect 543740 51128 543792 51134
rect 543740 51070 543792 51076
rect 540624 48929 540652 51070
rect 540610 48920 540666 48929
rect 540610 48855 540666 48864
rect 540334 34232 540390 34241
rect 540334 34167 540390 34176
rect 462320 28280 462372 28286
rect 462320 28222 462372 28228
rect 562336 6866 562364 315250
rect 566464 313948 566516 313954
rect 566464 313890 566516 313896
rect 566476 33114 566504 313890
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 569224 305992 569276 305998
rect 569224 305934 569276 305940
rect 569236 113150 569264 305934
rect 574744 303408 574796 303414
rect 574744 303350 574796 303356
rect 571984 301640 572036 301646
rect 571984 301582 572036 301588
rect 570696 294500 570748 294506
rect 570696 294442 570748 294448
rect 570604 268456 570656 268462
rect 570604 268398 570656 268404
rect 569224 113144 569276 113150
rect 569224 113086 569276 113092
rect 566464 33108 566516 33114
rect 566464 33050 566516 33056
rect 570616 20670 570644 268398
rect 570708 245614 570736 294442
rect 570696 245608 570748 245614
rect 570696 245550 570748 245556
rect 571996 86970 572024 301582
rect 573364 298036 573416 298042
rect 573364 297978 573416 297984
rect 573376 126954 573404 297978
rect 573364 126948 573416 126954
rect 573364 126890 573416 126896
rect 571984 86964 572036 86970
rect 571984 86906 572036 86912
rect 574756 46918 574784 303350
rect 580264 300008 580316 300014
rect 580264 299950 580316 299956
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 576124 295996 576176 296002
rect 576124 295938 576176 295944
rect 576136 206990 576164 295938
rect 579896 273216 579948 273222
rect 579896 273158 579948 273164
rect 579908 272241 579936 273158
rect 579894 272232 579950 272241
rect 579894 272167 579950 272176
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580276 219065 580304 299950
rect 580356 269816 580408 269822
rect 580356 269758 580408 269764
rect 580368 258913 580396 269758
rect 580354 258904 580410 258913
rect 580354 258839 580410 258848
rect 580262 219056 580318 219065
rect 580262 218991 580318 219000
rect 576124 206984 576176 206990
rect 576124 206926 576176 206932
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 574744 46912 574796 46918
rect 574744 46854 574796 46860
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 570604 20664 570656 20670
rect 570604 20606 570656 20612
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 562324 6860 562376 6866
rect 562324 6802 562376 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 460202 3360 460258 3369
rect 460202 3295 460258 3304
rect 360844 3198 360896 3204
rect 365074 3224 365130 3233
rect 365074 3159 365130 3168
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 24306 689288 24362 689344
rect 137834 700440 137890 700496
rect 105450 700304 105506 700360
rect 283838 692008 283894 692064
rect 3146 632032 3202 632088
rect 3238 579944 3294 580000
rect 3330 566888 3386 566944
rect 3514 658144 3570 658200
rect 3422 449520 3478 449576
rect 4066 553832 4122 553888
rect 3974 527856 4030 527912
rect 3882 514800 3938 514856
rect 20902 656240 20958 656296
rect 362222 678952 362278 679008
rect 21454 656240 21510 656296
rect 361762 667956 361818 667992
rect 361762 667936 361764 667956
rect 361764 667936 361816 667956
rect 361816 667936 361818 667956
rect 361762 656940 361818 656976
rect 361762 656920 361764 656940
rect 361764 656920 361816 656940
rect 361816 656920 361818 656940
rect 361762 645924 361818 645960
rect 361762 645904 361764 645924
rect 361764 645904 361816 645924
rect 361816 645904 361818 645924
rect 361578 634888 361634 634944
rect 361578 623872 361634 623928
rect 361578 612876 361634 612912
rect 361578 612856 361580 612876
rect 361580 612856 361632 612876
rect 361632 612856 361634 612876
rect 361762 601840 361818 601896
rect 361578 590844 361634 590880
rect 361578 590824 361580 590844
rect 361580 590824 361632 590844
rect 361632 590824 361634 590844
rect 361762 579808 361818 579864
rect 361578 568812 361634 568848
rect 361578 568792 361580 568812
rect 361580 568792 361632 568812
rect 361632 568792 361634 568812
rect 361670 557776 361726 557832
rect 361762 546760 361818 546816
rect 361762 535744 361818 535800
rect 361762 524728 361818 524784
rect 3790 501744 3846 501800
rect 3698 475632 3754 475688
rect 3606 462576 3662 462632
rect 3514 423544 3570 423600
rect 361762 513712 361818 513768
rect 361762 502696 361818 502752
rect 361762 491680 361818 491736
rect 361762 480664 361818 480720
rect 361762 469648 361818 469704
rect 361762 458632 361818 458688
rect 361762 447616 361818 447672
rect 361762 436600 361818 436656
rect 361762 425584 361818 425640
rect 361578 414568 361634 414624
rect 3974 410488 4030 410544
rect 361578 403552 361634 403608
rect 3790 397432 3846 397488
rect 3422 358400 3478 358456
rect 3606 345344 3662 345400
rect 3422 306176 3478 306232
rect 3330 293120 3386 293176
rect 3330 149776 3386 149832
rect 3238 136720 3294 136776
rect 3146 84632 3202 84688
rect 3146 71576 3202 71632
rect 3514 267144 3570 267200
rect 3422 58520 3478 58576
rect 2870 32408 2926 32464
rect 3606 254088 3662 254144
rect 3698 241032 3754 241088
rect 361578 392536 361634 392592
rect 361578 381520 361634 381576
rect 3882 371320 3938 371376
rect 3790 214920 3846 214976
rect 361578 370504 361634 370560
rect 362222 359488 362278 359544
rect 361762 348472 361818 348528
rect 361762 337456 361818 337512
rect 362222 326440 362278 326496
rect 3974 319232 4030 319288
rect 361762 315424 361818 315480
rect 3882 201864 3938 201920
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3974 188808 4030 188864
rect 4066 162832 4122 162888
rect 19246 49544 19302 49600
rect 20902 59880 20958 59936
rect 21454 59880 21510 59936
rect 359462 46552 359518 46608
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 2870 3576 2926 3632
rect 1674 3440 1730 3496
rect 570 3304 626 3360
rect 8758 3984 8814 4040
rect 9954 3712 10010 3768
rect 13542 3848 13598 3904
rect 17038 3168 17094 3224
rect 361762 304408 361818 304464
rect 362222 302776 362278 302832
rect 361762 293392 361818 293448
rect 361762 282376 361818 282432
rect 361762 271360 361818 271416
rect 361762 260344 361818 260400
rect 361762 249328 361818 249384
rect 361762 238312 361818 238368
rect 361762 227296 361818 227352
rect 361670 216316 361672 216336
rect 361672 216316 361724 216336
rect 361724 216316 361726 216336
rect 361670 216280 361726 216316
rect 361762 205264 361818 205320
rect 361762 194248 361818 194304
rect 361762 183232 361818 183288
rect 361762 172216 361818 172272
rect 361762 161200 361818 161256
rect 361762 150184 361818 150240
rect 361762 139168 361818 139224
rect 361762 128152 361818 128208
rect 361762 117136 361818 117192
rect 361762 106120 361818 106176
rect 361762 95140 361764 95160
rect 361764 95140 361816 95160
rect 361816 95140 361818 95160
rect 361762 95104 361818 95140
rect 361762 84124 361764 84144
rect 361764 84124 361816 84144
rect 361816 84124 361818 84144
rect 361762 84088 361818 84124
rect 361762 73108 361764 73128
rect 361764 73108 361816 73128
rect 361816 73108 361818 73128
rect 361762 73072 361818 73108
rect 361762 62076 361818 62112
rect 361762 62056 361764 62076
rect 361764 62056 361816 62076
rect 361816 62056 361818 62076
rect 361762 51076 361764 51096
rect 361764 51076 361816 51096
rect 361816 51076 361818 51096
rect 361762 51040 361818 51076
rect 362406 297608 362462 297664
rect 362222 3984 362278 4040
rect 365074 297472 365130 297528
rect 365350 297336 365406 297392
rect 370594 305632 370650 305688
rect 371974 294480 372030 294536
rect 378690 302912 378746 302968
rect 379150 303184 379206 303240
rect 379334 303048 379390 303104
rect 381910 306040 381966 306096
rect 381726 305904 381782 305960
rect 381542 305768 381598 305824
rect 380438 291760 380494 291816
rect 371974 3848 372030 3904
rect 381542 3576 381598 3632
rect 382094 306176 382150 306232
rect 385682 306856 385738 306912
rect 384394 46688 384450 46744
rect 384670 46824 384726 46880
rect 381726 3440 381782 3496
rect 427818 336776 427874 336832
rect 420458 334328 420514 334384
rect 424138 334328 424194 334384
rect 421838 162696 421894 162752
rect 425886 162696 425942 162752
rect 428646 162696 428702 162752
rect 432786 332832 432842 332888
rect 432694 329160 432750 329216
rect 432602 325488 432658 325544
rect 432878 321816 432934 321872
rect 432786 318144 432842 318200
rect 432602 314472 432658 314528
rect 432050 310800 432106 310856
rect 432694 307128 432750 307184
rect 445206 320048 445262 320104
rect 445574 683304 445630 683360
rect 446770 683168 446826 683224
rect 446678 322768 446734 322824
rect 446954 682760 447010 682816
rect 446770 319776 446826 319832
rect 447138 383596 447140 383616
rect 447140 383596 447192 383616
rect 447192 383596 447194 383616
rect 447138 383560 447194 383596
rect 447230 382880 447286 382936
rect 447138 382200 447194 382256
rect 447230 381520 447286 381576
rect 447230 380840 447286 380896
rect 447138 380160 447194 380216
rect 447138 378800 447194 378856
rect 447322 378120 447378 378176
rect 447138 377440 447194 377496
rect 447230 376760 447286 376816
rect 447138 376080 447194 376136
rect 447230 375400 447286 375456
rect 447138 374720 447194 374776
rect 447230 374040 447286 374096
rect 447138 373360 447194 373416
rect 447230 372680 447286 372736
rect 447138 372000 447194 372056
rect 447230 371320 447286 371376
rect 447138 370640 447194 370696
rect 447230 369960 447286 370016
rect 447138 369280 447194 369336
rect 447230 368600 447286 368656
rect 447138 367920 447194 367976
rect 447230 367240 447286 367296
rect 447138 366560 447194 366616
rect 447230 365880 447286 365936
rect 447230 365200 447286 365256
rect 447138 364520 447194 364576
rect 447230 363840 447286 363896
rect 447138 363160 447194 363216
rect 447138 362480 447194 362536
rect 447230 361800 447286 361856
rect 447230 361120 447286 361176
rect 447138 360440 447194 360496
rect 447138 359760 447194 359816
rect 447230 359080 447286 359136
rect 447506 379480 447562 379536
rect 447414 354320 447470 354376
rect 447598 353640 447654 353696
rect 447322 351600 447378 351656
rect 447138 350920 447194 350976
rect 447138 347520 447194 347576
rect 447138 342080 447194 342136
rect 447230 341400 447286 341456
rect 447230 340720 447286 340776
rect 447138 340040 447194 340096
rect 447230 339360 447286 339416
rect 447138 338680 447194 338736
rect 447138 337320 447194 337376
rect 447138 336640 447194 336696
rect 447230 335960 447286 336016
rect 447230 335280 447286 335336
rect 447138 334600 447194 334656
rect 447230 333920 447286 333976
rect 447138 333240 447194 333296
rect 447230 330520 447286 330576
rect 447506 338000 447562 338056
rect 447874 355000 447930 355056
rect 447966 352280 448022 352336
rect 447966 345480 448022 345536
rect 447874 344800 447930 344856
rect 447782 331200 447838 331256
rect 447690 330520 447746 330576
rect 447414 329840 447470 329896
rect 448150 352960 448206 353016
rect 448334 349560 448390 349616
rect 448242 348880 448298 348936
rect 449070 386960 449126 387016
rect 449070 357040 449126 357096
rect 448978 346840 449034 346896
rect 448426 343440 448482 343496
rect 448150 332560 448206 332616
rect 448334 331880 448390 331936
rect 448426 331200 448482 331256
rect 543462 700304 543518 700360
rect 527178 699760 527234 699816
rect 559654 699760 559710 699816
rect 580170 697176 580226 697232
rect 457810 667936 457866 667992
rect 457718 652840 457774 652896
rect 457626 650120 457682 650176
rect 457534 645904 457590 645960
rect 457442 643184 457498 643240
rect 457350 640328 457406 640384
rect 457258 637880 457314 637936
rect 450450 516840 450506 516896
rect 450450 514664 450506 514720
rect 458086 662496 458142 662552
rect 457994 659912 458050 659968
rect 457902 657464 457958 657520
rect 458822 635432 458878 635488
rect 458730 611360 458786 611416
rect 459006 633392 459062 633448
rect 458914 623872 458970 623928
rect 459098 630672 459154 630728
rect 458914 599528 458970 599584
rect 459190 628088 459246 628144
rect 459098 589872 459154 589928
rect 459282 625776 459338 625832
rect 459374 621016 459430 621072
rect 460202 618296 460258 618352
rect 459466 615984 459522 616040
rect 460110 613808 460166 613864
rect 460018 608640 460074 608696
rect 459926 606328 459982 606384
rect 459466 603608 459522 603664
rect 460110 601976 460166 602032
rect 458822 518064 458878 518120
rect 450542 512352 450598 512408
rect 450358 510176 450414 510232
rect 449990 507592 450046 507648
rect 449806 503444 449862 503500
rect 449346 348200 449402 348256
rect 449346 344120 449402 344176
rect 449622 357720 449678 357776
rect 449530 356360 449586 356416
rect 449806 358400 449862 358456
rect 449714 355680 449770 355736
rect 449806 350240 449862 350296
rect 449438 342760 449494 342816
rect 450082 505416 450138 505472
rect 450174 503240 450230 503296
rect 450266 337728 450322 337784
rect 449990 334056 450046 334112
rect 449898 328888 449954 328944
rect 449990 326576 450046 326632
rect 450266 336776 450322 336832
rect 450266 327936 450322 327992
rect 450634 505416 450690 505472
rect 450542 337728 450598 337784
rect 463054 517520 463110 517576
rect 463146 501064 463202 501120
rect 482742 517520 482798 517576
rect 492126 512420 492182 512476
rect 473726 462848 473782 462904
rect 489182 496848 489238 496904
rect 476118 428440 476174 428496
rect 472162 389000 472218 389056
rect 473634 389000 473690 389056
rect 472898 388864 472954 388920
rect 479522 389000 479578 389056
rect 494150 508816 494206 508872
rect 500958 516840 501014 516896
rect 502246 516840 502302 516896
rect 494334 515888 494390 515944
rect 507122 516704 507178 516760
rect 494242 505688 494298 505744
rect 495070 505724 495072 505744
rect 495072 505724 495124 505744
rect 495124 505724 495126 505744
rect 495070 505688 495126 505724
rect 494702 501200 494758 501256
rect 493322 395256 493378 395312
rect 509330 365200 509386 365256
rect 450542 334192 450598 334248
rect 450450 328616 450506 328672
rect 450542 327256 450598 327312
rect 510618 359080 510674 359136
rect 509514 357584 509570 357640
rect 509422 356088 509478 356144
rect 450634 325488 450690 325544
rect 450174 325216 450230 325272
rect 450542 324808 450598 324864
rect 450082 324536 450138 324592
rect 450634 324128 450690 324184
rect 509422 324944 509478 325000
rect 509330 322904 509386 322960
rect 458638 322496 458694 322552
rect 462226 322632 462282 322688
rect 461306 322496 461362 322552
rect 451738 158244 451740 158264
rect 451740 158244 451792 158264
rect 451792 158244 451794 158264
rect 451738 158208 451794 158244
rect 451738 156848 451794 156904
rect 451922 155488 451978 155544
rect 451922 154164 451924 154184
rect 451924 154164 451976 154184
rect 451976 154164 451978 154184
rect 451922 154128 451978 154164
rect 452014 151408 452070 151464
rect 451738 147364 451740 147384
rect 451740 147364 451792 147384
rect 451792 147364 451794 147384
rect 451738 147328 451794 147364
rect 451462 144608 451518 144664
rect 452106 132368 452162 132424
rect 451738 125568 451794 125624
rect 452382 152768 452438 152824
rect 452474 150048 452530 150104
rect 452566 148724 452568 148744
rect 452568 148724 452620 148744
rect 452620 148724 452622 148744
rect 452566 148688 452622 148724
rect 452566 146004 452568 146024
rect 452568 146004 452620 146024
rect 452620 146004 452622 146024
rect 452566 145968 452622 146004
rect 452566 143284 452568 143304
rect 452568 143284 452620 143304
rect 452620 143284 452622 143304
rect 452566 143248 452622 143284
rect 452566 141924 452568 141944
rect 452568 141924 452620 141944
rect 452620 141924 452622 141944
rect 452566 141888 452622 141924
rect 452566 140564 452568 140584
rect 452568 140564 452620 140584
rect 452620 140564 452622 140584
rect 452566 140528 452622 140564
rect 452566 139204 452568 139224
rect 452568 139204 452620 139224
rect 452620 139204 452622 139224
rect 452566 139168 452622 139204
rect 452566 137844 452568 137864
rect 452568 137844 452620 137864
rect 452620 137844 452622 137864
rect 452566 137808 452622 137844
rect 452566 136484 452568 136504
rect 452568 136484 452620 136504
rect 452620 136484 452622 136504
rect 452566 136448 452622 136484
rect 452566 135124 452568 135144
rect 452568 135124 452620 135144
rect 452620 135124 452622 135144
rect 452566 135088 452622 135124
rect 452566 133764 452568 133784
rect 452568 133764 452620 133784
rect 452620 133764 452622 133784
rect 452566 133728 452622 133764
rect 452290 131044 452292 131064
rect 452292 131044 452344 131064
rect 452344 131044 452346 131064
rect 452290 131008 452346 131044
rect 452382 129684 452384 129704
rect 452384 129684 452436 129704
rect 452436 129684 452438 129704
rect 452382 129648 452438 129684
rect 452198 128288 452254 128344
rect 452290 126948 452346 126984
rect 452290 126928 452292 126948
rect 452292 126928 452344 126948
rect 452344 126928 452346 126948
rect 452106 124208 452162 124264
rect 451830 122848 451886 122904
rect 456062 321816 456118 321872
rect 451738 121488 451794 121544
rect 456798 262656 456854 262712
rect 456798 248784 456854 248840
rect 456798 234912 456854 234968
rect 460018 321408 460074 321464
rect 460754 321952 460810 322008
rect 460202 319368 460258 319424
rect 457810 234912 457866 234968
rect 457902 221040 457958 221096
rect 460018 207304 460074 207360
rect 385774 3712 385830 3768
rect 462502 321272 462558 321328
rect 461950 321000 462006 321056
rect 480994 322632 481050 322688
rect 473450 322496 473506 322552
rect 473450 322396 473452 322416
rect 473452 322396 473504 322416
rect 473504 322396 473506 322416
rect 473450 322360 473506 322396
rect 480902 322496 480958 322552
rect 481546 322360 481602 322416
rect 470506 321272 470562 321328
rect 471610 319640 471666 319696
rect 472714 319912 472770 319968
rect 472990 319776 473046 319832
rect 482650 321136 482706 321192
rect 483202 320048 483258 320104
rect 496450 318008 496506 318064
rect 501970 319504 502026 319560
rect 503166 313928 503222 313984
rect 507030 320864 507086 320920
rect 507214 320728 507270 320784
rect 509422 322088 509478 322144
rect 509330 319368 509386 319424
rect 509606 343984 509662 344040
rect 509698 335824 509754 335880
rect 509882 333104 509938 333160
rect 510158 328072 510214 328128
rect 509606 303184 509662 303240
rect 510802 355816 510858 355872
rect 510710 353096 510766 353152
rect 510894 346024 510950 346080
rect 510986 342760 511042 342816
rect 511170 340040 511226 340096
rect 511078 337864 511134 337920
rect 512090 377576 512146 377632
rect 513286 384648 513342 384704
rect 512458 384104 512514 384160
rect 512642 383560 512698 383616
rect 513286 383016 513342 383072
rect 512458 382492 512514 382528
rect 512458 382472 512460 382492
rect 512460 382472 512512 382492
rect 512512 382472 512514 382492
rect 513102 381928 513158 381984
rect 512458 381384 512514 381440
rect 512550 379772 512606 379808
rect 512550 379752 512552 379772
rect 512552 379752 512604 379772
rect 512604 379752 512606 379772
rect 512826 379208 512882 379264
rect 512274 378120 512330 378176
rect 512826 377032 512882 377088
rect 512182 376488 512238 376544
rect 513194 380840 513250 380896
rect 513286 380296 513342 380352
rect 513286 378664 513342 378720
rect 513286 375964 513342 376000
rect 513286 375944 513288 375964
rect 513288 375944 513340 375964
rect 513340 375944 513342 375964
rect 513286 375420 513342 375456
rect 513286 375400 513288 375420
rect 513288 375400 513340 375420
rect 513340 375400 513342 375420
rect 511998 374856 512054 374912
rect 512090 374312 512146 374368
rect 511998 373768 512054 373824
rect 512458 373224 512514 373280
rect 512090 372700 512146 372736
rect 512090 372680 512092 372700
rect 512092 372680 512144 372700
rect 512144 372680 512146 372700
rect 512458 372136 512514 372192
rect 512090 371592 512146 371648
rect 511998 367784 512054 367840
rect 511998 366152 512054 366208
rect 511998 362364 512054 362400
rect 511998 362344 512000 362364
rect 512000 362344 512052 362364
rect 512052 362344 512054 362364
rect 511998 354184 512054 354240
rect 511998 352552 512054 352608
rect 511998 350376 512054 350432
rect 511998 349308 512054 349344
rect 511998 349288 512000 349308
rect 512000 349288 512052 349308
rect 512052 349288 512054 349308
rect 511998 338952 512054 339008
rect 511446 335688 511502 335744
rect 511814 327120 511870 327176
rect 511814 320864 511870 320920
rect 510986 306040 511042 306096
rect 510894 303048 510950 303104
rect 512826 371048 512882 371104
rect 512458 370504 512514 370560
rect 513286 369960 513342 370016
rect 513286 369416 513342 369472
rect 512826 368872 512882 368928
rect 512182 368328 512238 368384
rect 513286 367260 513342 367296
rect 513286 367240 513288 367260
rect 513288 367240 513340 367260
rect 513340 367240 513342 367260
rect 513286 366696 513342 366752
rect 513286 365064 513342 365120
rect 512642 364520 512698 364576
rect 513286 363568 513342 363624
rect 512458 363432 512514 363488
rect 513010 362888 513066 362944
rect 512274 361800 512330 361856
rect 513194 361256 513250 361312
rect 512366 360732 512422 360768
rect 512366 360712 512368 360732
rect 512368 360712 512420 360732
rect 512420 360712 512422 360732
rect 512918 360168 512974 360224
rect 512734 359624 512790 359680
rect 512366 358536 512422 358592
rect 513286 357992 513342 358048
rect 513286 356904 513342 356960
rect 512458 355272 512514 355328
rect 513286 354728 513342 354784
rect 513286 353640 513342 353696
rect 513286 352008 513342 352064
rect 512642 351464 512698 351520
rect 512550 350920 512606 350976
rect 513286 349832 513342 349888
rect 513286 348744 513342 348800
rect 512918 348200 512974 348256
rect 512550 347656 512606 347712
rect 513286 347112 513342 347168
rect 513286 346568 513342 346624
rect 512550 345480 512606 345536
rect 513010 344936 513066 344992
rect 512826 343848 512882 343904
rect 513010 343304 513066 343360
rect 512826 342216 512882 342272
rect 512642 340584 512698 340640
rect 512642 339516 512698 339552
rect 512642 339496 512644 339516
rect 512644 339496 512696 339516
rect 512696 339496 512698 339516
rect 512734 334600 512790 334656
rect 512642 331356 512698 331392
rect 512642 331336 512644 331356
rect 512644 331336 512696 331356
rect 512696 331336 512698 331356
rect 512642 329160 512698 329216
rect 513286 341672 513342 341728
rect 513286 341148 513342 341184
rect 513286 341128 513288 341148
rect 513288 341128 513340 341148
rect 513340 341128 513342 341148
rect 513010 338428 513066 338464
rect 513010 338408 513012 338428
rect 513012 338408 513064 338428
rect 513064 338408 513066 338428
rect 513286 337320 513342 337376
rect 513194 336776 513250 336832
rect 513010 335144 513066 335200
rect 513286 334056 513342 334112
rect 513194 331880 513250 331936
rect 512918 326984 512974 327040
rect 513470 330792 513526 330848
rect 512826 302776 512882 302832
rect 513838 302912 513894 302968
rect 516966 320728 517022 320784
rect 517978 305632 518034 305688
rect 547878 516704 547934 516760
rect 521750 462848 521806 462904
rect 557538 442856 557594 442912
rect 580262 683848 580318 683904
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579618 590960 579674 591016
rect 579618 577632 579674 577688
rect 579894 564304 579950 564360
rect 579618 511264 579674 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 579618 431568 579674 431624
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 325216 580226 325272
rect 580354 670656 580410 670712
rect 580446 537784 580502 537840
rect 580538 524456 580594 524512
rect 580630 418240 580686 418296
rect 580722 404912 580778 404968
rect 580814 351872 580870 351928
rect 531410 261024 531466 261080
rect 531318 243616 531374 243672
rect 530122 226208 530178 226264
rect 529938 209208 529994 209264
rect 460386 67632 460442 67688
rect 460846 67632 460902 67688
rect 539322 137672 539378 137728
rect 539506 135904 539562 135960
rect 539690 121352 539746 121408
rect 539782 119584 539838 119640
rect 539598 113192 539654 113248
rect 539966 108704 540022 108760
rect 540242 123120 540298 123176
rect 540150 114960 540206 115016
rect 540058 104624 540114 104680
rect 539874 97144 539930 97200
rect 536838 40976 536894 41032
rect 541070 110880 541126 110936
rect 541438 117000 541494 117056
rect 541346 106800 541402 106856
rect 541254 102720 541310 102776
rect 542726 129240 542782 129296
rect 542634 98640 542690 98696
rect 542910 100680 542966 100736
rect 542818 94560 542874 94616
rect 542542 92520 542598 92576
rect 542450 90480 542506 90536
rect 543278 137808 543334 137864
rect 543186 131280 543242 131336
rect 543094 127200 543150 127256
rect 543278 125160 543334 125216
rect 543002 88440 543058 88496
rect 541162 86400 541218 86456
rect 540978 82320 541034 82376
rect 540610 48864 540666 48920
rect 540334 34176 540390 34232
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 579894 272176 579950 272232
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580170 232328 580226 232384
rect 580354 258848 580410 258904
rect 580262 219000 580318 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
rect 460202 3304 460258 3360
rect 365074 3168 365130 3224
<< metal3 >>
rect 137829 700498 137895 700501
rect 449566 700498 449572 700500
rect 137829 700496 449572 700498
rect 137829 700440 137834 700496
rect 137890 700440 449572 700496
rect 137829 700438 449572 700440
rect 137829 700435 137895 700438
rect 449566 700436 449572 700438
rect 449636 700436 449642 700500
rect 105445 700362 105511 700365
rect 444230 700362 444236 700364
rect 105445 700360 444236 700362
rect 105445 700304 105450 700360
rect 105506 700304 444236 700360
rect 105445 700302 444236 700304
rect 105445 700299 105511 700302
rect 444230 700300 444236 700302
rect 444300 700300 444306 700364
rect 530526 700300 530532 700364
rect 530596 700362 530602 700364
rect 543457 700362 543523 700365
rect 530596 700360 543523 700362
rect 530596 700304 543462 700360
rect 543518 700304 543523 700360
rect 530596 700302 543523 700304
rect 530596 700300 530602 700302
rect 543457 700299 543523 700302
rect 526294 699756 526300 699820
rect 526364 699818 526370 699820
rect 527173 699818 527239 699821
rect 526364 699816 527239 699818
rect 526364 699760 527178 699816
rect 527234 699760 527239 699816
rect 526364 699758 527239 699760
rect 526364 699756 526370 699758
rect 527173 699755 527239 699758
rect 558126 699756 558132 699820
rect 558196 699818 558202 699820
rect 559649 699818 559715 699821
rect 558196 699816 559715 699818
rect 558196 699760 559654 699816
rect 559710 699760 559715 699816
rect 558196 699758 559715 699760
rect 558196 699756 558202 699758
rect 559649 699755 559715 699758
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect 283833 692066 283899 692069
rect 447726 692066 447732 692068
rect 283833 692064 447732 692066
rect 283833 692008 283838 692064
rect 283894 692008 447732 692064
rect 283833 692006 447732 692008
rect 283833 692003 283899 692006
rect 447726 692004 447732 692006
rect 447796 692004 447802 692068
rect 24301 689346 24367 689349
rect 446254 689346 446260 689348
rect 24301 689344 446260 689346
rect 24301 689288 24306 689344
rect 24362 689288 446260 689344
rect 24301 689286 446260 689288
rect 24301 689283 24367 689286
rect 446254 689284 446260 689286
rect 446324 689284 446330 689348
rect -960 684314 480 684404
rect 447910 684314 447916 684316
rect -960 684254 447916 684314
rect -960 684164 480 684254
rect 447910 684252 447916 684254
rect 447980 684252 447986 684316
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect 3550 683300 3556 683364
rect 3620 683362 3626 683364
rect 445569 683362 445635 683365
rect 3620 683360 445635 683362
rect 3620 683304 445574 683360
rect 445630 683304 445635 683360
rect 3620 683302 445635 683304
rect 3620 683300 3626 683302
rect 445569 683299 445635 683302
rect 3734 683164 3740 683228
rect 3804 683226 3810 683228
rect 446765 683226 446831 683229
rect 3804 683224 446831 683226
rect 3804 683168 446770 683224
rect 446826 683168 446831 683224
rect 3804 683166 446831 683168
rect 3804 683164 3810 683166
rect 446765 683163 446831 683166
rect 3366 682756 3372 682820
rect 3436 682818 3442 682820
rect 446949 682818 447015 682821
rect 3436 682816 447015 682818
rect 3436 682760 446954 682816
rect 447010 682760 447015 682816
rect 3436 682758 447015 682760
rect 3436 682756 3442 682758
rect 446949 682755 447015 682758
rect 362217 679010 362283 679013
rect 359812 679008 362283 679010
rect 359812 678952 362222 679008
rect 362278 678952 362283 679008
rect 359812 678950 362283 678952
rect 362217 678947 362283 678950
rect -960 671258 480 671348
rect 3734 671258 3740 671260
rect -960 671198 3740 671258
rect -960 671108 480 671198
rect 3734 671196 3740 671198
rect 3804 671196 3810 671260
rect 580349 670714 580415 670717
rect 583520 670714 584960 670804
rect 580349 670712 584960 670714
rect 580349 670656 580354 670712
rect 580410 670656 584960 670712
rect 580349 670654 584960 670656
rect 580349 670651 580415 670654
rect 583520 670564 584960 670654
rect 361757 667994 361823 667997
rect 359812 667992 361823 667994
rect 359812 667936 361762 667992
rect 361818 667936 361823 667992
rect 359812 667934 361823 667936
rect 361757 667931 361823 667934
rect 457805 667994 457871 667997
rect 457805 667992 460092 667994
rect 457805 667936 457810 667992
rect 457866 667936 460092 667992
rect 457805 667934 460092 667936
rect 457805 667931 457871 667934
rect 458030 665212 458036 665276
rect 458100 665274 458106 665276
rect 460062 665274 460122 665448
rect 458100 665214 460122 665274
rect 458100 665212 458106 665214
rect 458081 662554 458147 662557
rect 460062 662554 460122 663000
rect 458081 662552 460122 662554
rect 458081 662496 458086 662552
rect 458142 662496 460122 662552
rect 458081 662494 460122 662496
rect 458081 662491 458147 662494
rect 457989 659970 458055 659973
rect 460062 659970 460122 660552
rect 457989 659968 460122 659970
rect 457989 659912 457994 659968
rect 458050 659912 460122 659968
rect 457989 659910 460122 659912
rect 457989 659907 458055 659910
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 457897 657522 457963 657525
rect 460062 657522 460122 658104
rect 457897 657520 460122 657522
rect 457897 657464 457902 657520
rect 457958 657464 460122 657520
rect 457897 657462 460122 657464
rect 457897 657459 457963 657462
rect 583520 657236 584960 657476
rect 361757 656978 361823 656981
rect 359812 656976 361823 656978
rect 359812 656920 361762 656976
rect 361818 656920 361823 656976
rect 359812 656918 361823 656920
rect 361757 656915 361823 656918
rect 20897 656298 20963 656301
rect 21449 656298 21515 656301
rect 20897 656296 21515 656298
rect 20897 656240 20902 656296
rect 20958 656240 21454 656296
rect 21510 656240 21515 656296
rect 20897 656238 21515 656240
rect 20897 656235 20963 656238
rect 21449 656235 21515 656238
rect 459134 655692 459140 655756
rect 459204 655754 459210 655756
rect 459204 655694 460092 655754
rect 459204 655692 459210 655694
rect 457713 652898 457779 652901
rect 460062 652898 460122 653208
rect 457713 652896 460122 652898
rect 457713 652840 457718 652896
rect 457774 652840 460122 652896
rect 457713 652838 460122 652840
rect 457713 652835 457779 652838
rect 457621 650178 457687 650181
rect 460062 650178 460122 650760
rect 457621 650176 460122 650178
rect 457621 650120 457626 650176
rect 457682 650120 460122 650176
rect 457621 650118 460122 650120
rect 457621 650115 457687 650118
rect 458950 647668 458956 647732
rect 459020 647730 459026 647732
rect 460062 647730 460122 648312
rect 459020 647670 460122 647730
rect 459020 647668 459026 647670
rect 361757 645962 361823 645965
rect 359812 645960 361823 645962
rect 359812 645904 361762 645960
rect 361818 645904 361823 645960
rect 359812 645902 361823 645904
rect 361757 645899 361823 645902
rect 457529 645962 457595 645965
rect 457529 645960 460092 645962
rect 457529 645904 457534 645960
rect 457590 645904 460092 645960
rect 457529 645902 460092 645904
rect 457529 645899 457595 645902
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect 457437 643242 457503 643245
rect 460062 643242 460122 643416
rect 457437 643240 460122 643242
rect 457437 643184 457442 643240
rect 457498 643184 460122 643240
rect 457437 643182 460122 643184
rect 457437 643179 457503 643182
rect 457345 640386 457411 640389
rect 460062 640386 460122 640968
rect 457345 640384 460122 640386
rect 457345 640328 457350 640384
rect 457406 640328 460122 640384
rect 457345 640326 460122 640328
rect 457345 640323 457411 640326
rect 457253 637938 457319 637941
rect 460062 637938 460122 638520
rect 457253 637936 460122 637938
rect 457253 637880 457258 637936
rect 457314 637880 460122 637936
rect 457253 637878 460122 637880
rect 457253 637875 457319 637878
rect 458817 635490 458883 635493
rect 460062 635490 460122 636072
rect 458817 635488 460122 635490
rect 458817 635432 458822 635488
rect 458878 635432 460122 635488
rect 458817 635430 460122 635432
rect 458817 635427 458883 635430
rect 361573 634946 361639 634949
rect 359812 634944 361639 634946
rect 359812 634888 361578 634944
rect 361634 634888 361639 634944
rect 359812 634886 361639 634888
rect 361573 634883 361639 634886
rect 459001 633450 459067 633453
rect 460062 633450 460122 633624
rect 459001 633448 460122 633450
rect 459001 633392 459006 633448
rect 459062 633392 460122 633448
rect 459001 633390 460122 633392
rect 459001 633387 459067 633390
rect -960 632090 480 632180
rect 3141 632090 3207 632093
rect -960 632088 3207 632090
rect -960 632032 3146 632088
rect 3202 632032 3207 632088
rect -960 632030 3207 632032
rect -960 631940 480 632030
rect 3141 632027 3207 632030
rect 459093 630730 459159 630733
rect 460062 630730 460122 631176
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 459093 630728 460122 630730
rect 459093 630672 459098 630728
rect 459154 630672 460122 630728
rect 583520 630716 584960 630806
rect 459093 630670 460122 630672
rect 459093 630667 459159 630670
rect 459185 628146 459251 628149
rect 460062 628146 460122 628728
rect 459185 628144 460122 628146
rect 459185 628088 459190 628144
rect 459246 628088 460122 628144
rect 459185 628086 460122 628088
rect 459185 628083 459251 628086
rect 459277 625834 459343 625837
rect 460062 625834 460122 626280
rect 459277 625832 460122 625834
rect 459277 625776 459282 625832
rect 459338 625776 460122 625832
rect 459277 625774 460122 625776
rect 459277 625771 459343 625774
rect 361573 623930 361639 623933
rect 359812 623928 361639 623930
rect 359812 623872 361578 623928
rect 361634 623872 361639 623928
rect 359812 623870 361639 623872
rect 361573 623867 361639 623870
rect 458909 623930 458975 623933
rect 458909 623928 460092 623930
rect 458909 623872 458914 623928
rect 458970 623872 460092 623928
rect 458909 623870 460092 623872
rect 458909 623867 458975 623870
rect 459369 621074 459435 621077
rect 460062 621074 460122 621384
rect 459369 621072 460122 621074
rect 459369 621016 459374 621072
rect 459430 621016 460122 621072
rect 459369 621014 460122 621016
rect 459369 621011 459435 621014
rect -960 619170 480 619260
rect 3550 619170 3556 619172
rect -960 619110 3556 619170
rect -960 619020 480 619110
rect 3550 619108 3556 619110
rect 3620 619108 3626 619172
rect 460062 618354 460122 618936
rect 460197 618354 460263 618357
rect 460062 618352 460263 618354
rect 460062 618296 460202 618352
rect 460258 618296 460263 618352
rect 460062 618294 460263 618296
rect 460197 618291 460263 618294
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 459461 616042 459527 616045
rect 460062 616042 460122 616488
rect 459461 616040 460122 616042
rect 459461 615984 459466 616040
rect 459522 615984 460122 616040
rect 459461 615982 460122 615984
rect 459461 615979 459527 615982
rect 460062 613869 460122 614040
rect 460062 613864 460171 613869
rect 460062 613808 460110 613864
rect 460166 613808 460171 613864
rect 460062 613806 460171 613808
rect 460105 613803 460171 613806
rect 361573 612914 361639 612917
rect 359812 612912 361639 612914
rect 359812 612856 361578 612912
rect 361634 612856 361639 612912
rect 359812 612854 361639 612856
rect 361573 612851 361639 612854
rect 458725 611418 458791 611421
rect 460062 611418 460122 611592
rect 458725 611416 460122 611418
rect 458725 611360 458730 611416
rect 458786 611360 460122 611416
rect 458725 611358 460122 611360
rect 458725 611355 458791 611358
rect 460062 608701 460122 609144
rect 460013 608696 460122 608701
rect 460013 608640 460018 608696
rect 460074 608640 460122 608696
rect 460013 608638 460122 608640
rect 460013 608635 460079 608638
rect 459921 606386 459987 606389
rect 460062 606386 460122 606696
rect 459921 606384 460122 606386
rect 459921 606328 459926 606384
rect 459982 606328 460122 606384
rect 459921 606326 460122 606328
rect 459921 606323 459987 606326
rect -960 606114 480 606204
rect 3366 606114 3372 606116
rect -960 606054 3372 606114
rect -960 605964 480 606054
rect 3366 606052 3372 606054
rect 3436 606052 3442 606116
rect 459461 603666 459527 603669
rect 460062 603666 460122 604248
rect 583520 604060 584960 604300
rect 459461 603664 460122 603666
rect 459461 603608 459466 603664
rect 459522 603608 460122 603664
rect 459461 603606 460122 603608
rect 459461 603603 459527 603606
rect 460105 602034 460171 602037
rect 460062 602032 460171 602034
rect 460062 601976 460110 602032
rect 460166 601976 460171 602032
rect 460062 601971 460171 601976
rect 361757 601898 361823 601901
rect 359812 601896 361823 601898
rect 359812 601840 361762 601896
rect 361818 601840 361823 601896
rect 460062 601868 460122 601971
rect 359812 601838 361823 601840
rect 361757 601835 361823 601838
rect 458909 599586 458975 599589
rect 472014 599586 472020 599588
rect 458909 599584 472020 599586
rect 458909 599528 458914 599584
rect 458970 599528 472020 599584
rect 458909 599526 472020 599528
rect 458909 599523 458975 599526
rect 472014 599524 472020 599526
rect 472084 599524 472090 599588
rect 459134 598164 459140 598228
rect 459204 598226 459210 598228
rect 478822 598226 478828 598228
rect 459204 598166 478828 598226
rect 459204 598164 459210 598166
rect 478822 598164 478828 598166
rect 478892 598164 478898 598228
rect -960 592908 480 593148
rect 579613 591018 579679 591021
rect 583520 591018 584960 591108
rect 579613 591016 584960 591018
rect 579613 590960 579618 591016
rect 579674 590960 584960 591016
rect 579613 590958 584960 590960
rect 579613 590955 579679 590958
rect 361573 590882 361639 590885
rect 359812 590880 361639 590882
rect 359812 590824 361578 590880
rect 361634 590824 361639 590880
rect 583520 590868 584960 590958
rect 359812 590822 361639 590824
rect 361573 590819 361639 590822
rect 459093 589930 459159 589933
rect 472198 589930 472204 589932
rect 459093 589928 472204 589930
rect 459093 589872 459098 589928
rect 459154 589872 472204 589928
rect 459093 589870 472204 589872
rect 459093 589867 459159 589870
rect 472198 589868 472204 589870
rect 472268 589868 472274 589932
rect -960 580002 480 580092
rect 3233 580002 3299 580005
rect -960 580000 3299 580002
rect -960 579944 3238 580000
rect 3294 579944 3299 580000
rect -960 579942 3299 579944
rect -960 579852 480 579942
rect 3233 579939 3299 579942
rect 361757 579866 361823 579869
rect 359812 579864 361823 579866
rect 359812 579808 361762 579864
rect 361818 579808 361823 579864
rect 359812 579806 361823 579808
rect 361757 579803 361823 579806
rect 579613 577690 579679 577693
rect 583520 577690 584960 577780
rect 579613 577688 584960 577690
rect 579613 577632 579618 577688
rect 579674 577632 584960 577688
rect 579613 577630 584960 577632
rect 579613 577627 579679 577630
rect 583520 577540 584960 577630
rect 361573 568850 361639 568853
rect 359812 568848 361639 568850
rect 359812 568792 361578 568848
rect 361634 568792 361639 568848
rect 359812 568790 361639 568792
rect 361573 568787 361639 568790
rect -960 566946 480 567036
rect 3325 566946 3391 566949
rect -960 566944 3391 566946
rect -960 566888 3330 566944
rect 3386 566888 3391 566944
rect -960 566886 3391 566888
rect -960 566796 480 566886
rect 3325 566883 3391 566886
rect 579889 564362 579955 564365
rect 583520 564362 584960 564452
rect 579889 564360 584960 564362
rect 579889 564304 579894 564360
rect 579950 564304 584960 564360
rect 579889 564302 584960 564304
rect 579889 564299 579955 564302
rect 583520 564212 584960 564302
rect 361665 557834 361731 557837
rect 359812 557832 361731 557834
rect 359812 557776 361670 557832
rect 361726 557776 361731 557832
rect 359812 557774 361731 557776
rect 361665 557771 361731 557774
rect -960 553890 480 553980
rect 4061 553890 4127 553893
rect -960 553888 4127 553890
rect -960 553832 4066 553888
rect 4122 553832 4127 553888
rect -960 553830 4127 553832
rect -960 553740 480 553830
rect 4061 553827 4127 553830
rect 583520 551020 584960 551260
rect 361757 546818 361823 546821
rect 359812 546816 361823 546818
rect 359812 546760 361762 546816
rect 361818 546760 361823 546816
rect 359812 546758 361823 546760
rect 361757 546755 361823 546758
rect -960 540684 480 540924
rect 580441 537842 580507 537845
rect 583520 537842 584960 537932
rect 580441 537840 584960 537842
rect 580441 537784 580446 537840
rect 580502 537784 584960 537840
rect 580441 537782 584960 537784
rect 580441 537779 580507 537782
rect 583520 537692 584960 537782
rect 361757 535802 361823 535805
rect 359812 535800 361823 535802
rect 359812 535744 361762 535800
rect 361818 535744 361823 535800
rect 359812 535742 361823 535744
rect 361757 535739 361823 535742
rect -960 527914 480 528004
rect 3969 527914 4035 527917
rect -960 527912 4035 527914
rect -960 527856 3974 527912
rect 4030 527856 4035 527912
rect -960 527854 4035 527856
rect -960 527764 480 527854
rect 3969 527851 4035 527854
rect 361757 524786 361823 524789
rect 359812 524784 361823 524786
rect 359812 524728 361762 524784
rect 361818 524728 361823 524784
rect 359812 524726 361823 524728
rect 361757 524723 361823 524726
rect 580533 524514 580599 524517
rect 583520 524514 584960 524604
rect 580533 524512 584960 524514
rect 580533 524456 580538 524512
rect 580594 524456 584960 524512
rect 580533 524454 584960 524456
rect 580533 524451 580599 524454
rect 583520 524364 584960 524454
rect 458817 518122 458883 518125
rect 474406 518122 474412 518124
rect 458817 518120 474412 518122
rect 458817 518064 458822 518120
rect 458878 518064 474412 518120
rect 458817 518062 474412 518064
rect 458817 518059 458883 518062
rect 474406 518060 474412 518062
rect 474476 518060 474482 518124
rect 458030 517516 458036 517580
rect 458100 517578 458106 517580
rect 463049 517578 463115 517581
rect 482737 517580 482803 517581
rect 458100 517576 463115 517578
rect 458100 517520 463054 517576
rect 463110 517520 463115 517576
rect 458100 517518 463115 517520
rect 458100 517516 458106 517518
rect 463049 517515 463115 517518
rect 482686 517516 482692 517580
rect 482756 517578 482803 517580
rect 482756 517576 482848 517578
rect 482798 517520 482848 517576
rect 482756 517518 482848 517520
rect 482756 517516 482803 517518
rect 482737 517515 482803 517516
rect 450445 516898 450511 516901
rect 500953 516898 501019 516901
rect 502241 516898 502307 516901
rect 450445 516896 502307 516898
rect 450445 516840 450450 516896
rect 450506 516840 500958 516896
rect 501014 516840 502246 516896
rect 502302 516840 502307 516896
rect 450445 516838 502307 516840
rect 450445 516835 450511 516838
rect 500953 516835 501019 516838
rect 502241 516835 502307 516838
rect 451038 516762 451044 516764
rect 450678 516702 451044 516762
rect 450678 516528 450738 516702
rect 451038 516700 451044 516702
rect 451108 516762 451114 516764
rect 507117 516762 507183 516765
rect 547873 516762 547939 516765
rect 451108 516760 547939 516762
rect 451108 516704 507122 516760
rect 507178 516704 547878 516760
rect 547934 516704 547939 516760
rect 451108 516702 547939 516704
rect 451108 516700 451114 516702
rect 507117 516699 507183 516702
rect 547873 516699 547939 516702
rect 491894 515946 491954 515984
rect 494329 515946 494395 515949
rect 491894 515944 494395 515946
rect 491894 515888 494334 515944
rect 494390 515888 494395 515944
rect 491894 515886 494395 515888
rect 494329 515883 494395 515886
rect -960 514858 480 514948
rect 3877 514858 3943 514861
rect -960 514856 3943 514858
rect -960 514800 3882 514856
rect 3938 514800 3943 514856
rect -960 514798 3943 514800
rect -960 514708 480 514798
rect 3877 514795 3943 514798
rect 450445 514722 450511 514725
rect 450445 514720 450554 514722
rect 450445 514664 450450 514720
rect 450506 514664 450554 514720
rect 450445 514659 450554 514664
rect 450494 514384 450554 514659
rect 450486 514320 450492 514384
rect 450556 514320 450562 514384
rect 361757 513770 361823 513773
rect 359812 513768 361823 513770
rect 359812 513712 361762 513768
rect 361818 513712 361823 513768
rect 359812 513710 361823 513712
rect 361757 513707 361823 513710
rect 492121 512478 492187 512481
rect 491924 512476 492187 512478
rect 491924 512420 492126 512476
rect 492182 512420 492187 512476
rect 491924 512418 492187 512420
rect 492121 512415 492187 512418
rect 450537 512410 450603 512413
rect 450494 512408 450603 512410
rect 450494 512352 450542 512408
rect 450598 512352 450603 512408
rect 450494 512347 450603 512352
rect 450494 512176 450554 512347
rect 579613 511322 579679 511325
rect 583520 511322 584960 511412
rect 579613 511320 584960 511322
rect 579613 511264 579618 511320
rect 579674 511264 584960 511320
rect 579613 511262 584960 511264
rect 579613 511259 579679 511262
rect 583520 511172 584960 511262
rect 450353 510234 450419 510237
rect 450310 510232 450419 510234
rect 450310 510176 450358 510232
rect 450414 510176 450419 510232
rect 450310 510171 450419 510176
rect 450310 510000 450370 510171
rect 491894 508874 491954 508912
rect 494145 508874 494211 508877
rect 491894 508872 494211 508874
rect 491894 508816 494150 508872
rect 494206 508816 494211 508872
rect 491894 508814 494211 508816
rect 494145 508811 494211 508814
rect 449985 507650 450051 507653
rect 450126 507650 450186 507824
rect 449985 507648 450186 507650
rect 449985 507592 449990 507648
rect 450046 507592 450186 507648
rect 449985 507590 450186 507592
rect 449985 507587 450051 507590
rect 494237 505746 494303 505749
rect 495065 505746 495131 505749
rect 491894 505744 495131 505746
rect 491894 505688 494242 505744
rect 494298 505688 495070 505744
rect 495126 505688 495131 505744
rect 491894 505686 495131 505688
rect 450126 505477 450186 505648
rect 450077 505474 450186 505477
rect 450629 505474 450695 505477
rect 450077 505472 450695 505474
rect 450077 505416 450082 505472
rect 450138 505416 450634 505472
rect 450690 505416 450695 505472
rect 450077 505414 450695 505416
rect 450077 505411 450143 505414
rect 450629 505411 450695 505414
rect 491894 505376 491954 505686
rect 494237 505683 494303 505686
rect 495065 505683 495131 505686
rect 449801 503502 449867 503505
rect 449801 503500 450156 503502
rect 449801 503444 449806 503500
rect 449862 503472 450156 503500
rect 449862 503444 450186 503472
rect 449801 503442 450186 503444
rect 449801 503439 449867 503442
rect 450126 503301 450186 503442
rect 450126 503296 450235 503301
rect 450126 503240 450174 503296
rect 450230 503240 450235 503296
rect 450126 503238 450235 503240
rect 450169 503235 450235 503238
rect 361757 502754 361823 502757
rect 359812 502752 361823 502754
rect 359812 502696 361762 502752
rect 361818 502696 361823 502752
rect 359812 502694 361823 502696
rect 361757 502691 361823 502694
rect -960 501802 480 501892
rect 3785 501802 3851 501805
rect -960 501800 3851 501802
rect -960 501744 3790 501800
rect 3846 501744 3851 501800
rect -960 501742 3851 501744
rect -960 501652 480 501742
rect 3785 501739 3851 501742
rect 491894 501666 491954 501840
rect 470550 501606 491954 501666
rect 450678 501122 450738 501296
rect 463141 501122 463207 501125
rect 470550 501122 470610 501606
rect 491894 501258 491954 501606
rect 494697 501258 494763 501261
rect 491894 501256 494763 501258
rect 491894 501200 494702 501256
rect 494758 501200 494763 501256
rect 491894 501198 494763 501200
rect 494697 501195 494763 501198
rect 450678 501120 470610 501122
rect 450678 501064 463146 501120
rect 463202 501064 470610 501120
rect 450678 501062 470610 501064
rect 463141 501059 463207 501062
rect 583520 497844 584960 498084
rect 489177 496906 489243 496909
rect 489310 496906 489316 496908
rect 489177 496904 489316 496906
rect 489177 496848 489182 496904
rect 489238 496848 489316 496904
rect 489177 496846 489316 496848
rect 489177 496843 489243 496846
rect 489310 496844 489316 496846
rect 489380 496844 489386 496908
rect 361757 491738 361823 491741
rect 359812 491736 361823 491738
rect 359812 491680 361762 491736
rect 361818 491680 361823 491736
rect 359812 491678 361823 491680
rect 361757 491675 361823 491678
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 361757 480722 361823 480725
rect 359812 480720 361823 480722
rect 359812 480664 361762 480720
rect 361818 480664 361823 480720
rect 359812 480662 361823 480664
rect 361757 480659 361823 480662
rect -960 475690 480 475780
rect 3693 475690 3759 475693
rect -960 475688 3759 475690
rect -960 475632 3698 475688
rect 3754 475632 3759 475688
rect -960 475630 3759 475632
rect -960 475540 480 475630
rect 3693 475627 3759 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect 361757 469706 361823 469709
rect 359812 469704 361823 469706
rect 359812 469648 361762 469704
rect 361818 469648 361823 469704
rect 359812 469646 361823 469648
rect 361757 469643 361823 469646
rect 473721 462906 473787 462909
rect 482686 462906 482692 462908
rect 473721 462904 482692 462906
rect 473721 462848 473726 462904
rect 473782 462848 482692 462904
rect 473721 462846 482692 462848
rect 473721 462843 473787 462846
rect 482686 462844 482692 462846
rect 482756 462906 482762 462908
rect 521745 462906 521811 462909
rect 482756 462904 521811 462906
rect 482756 462848 521750 462904
rect 521806 462848 521811 462904
rect 482756 462846 521811 462848
rect 482756 462844 482762 462846
rect 521745 462843 521811 462846
rect -960 462634 480 462724
rect 3601 462634 3667 462637
rect -960 462632 3667 462634
rect -960 462576 3606 462632
rect 3662 462576 3667 462632
rect -960 462574 3667 462576
rect -960 462484 480 462574
rect 3601 462571 3667 462574
rect 361757 458690 361823 458693
rect 359812 458688 361823 458690
rect 359812 458632 361762 458688
rect 361818 458632 361823 458688
rect 359812 458630 361823 458632
rect 361757 458627 361823 458630
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3417 449578 3483 449581
rect -960 449576 3483 449578
rect -960 449520 3422 449576
rect 3478 449520 3483 449576
rect -960 449518 3483 449520
rect -960 449428 480 449518
rect 3417 449515 3483 449518
rect 361757 447674 361823 447677
rect 359812 447672 361823 447674
rect 359812 447616 361762 447672
rect 361818 447616 361823 447672
rect 359812 447614 361823 447616
rect 361757 447611 361823 447614
rect 583520 444668 584960 444908
rect 557533 442914 557599 442917
rect 555956 442912 557599 442914
rect 555956 442856 557538 442912
rect 557594 442856 557599 442912
rect 555956 442854 557599 442856
rect 557533 442851 557599 442854
rect -960 436508 480 436748
rect 361757 436658 361823 436661
rect 359812 436656 361823 436658
rect 359812 436600 361762 436656
rect 361818 436600 361823 436656
rect 359812 436598 361823 436600
rect 361757 436595 361823 436598
rect 579613 431626 579679 431629
rect 583520 431626 584960 431716
rect 579613 431624 584960 431626
rect 579613 431568 579618 431624
rect 579674 431568 584960 431624
rect 579613 431566 584960 431568
rect 579613 431563 579679 431566
rect 583520 431476 584960 431566
rect 458950 428436 458956 428500
rect 459020 428498 459026 428500
rect 476113 428498 476179 428501
rect 459020 428496 476179 428498
rect 459020 428440 476118 428496
rect 476174 428440 476179 428496
rect 459020 428438 476179 428440
rect 459020 428436 459026 428438
rect 476113 428435 476179 428438
rect 361757 425642 361823 425645
rect 359812 425640 361823 425642
rect 359812 425584 361762 425640
rect 361818 425584 361823 425640
rect 359812 425582 361823 425584
rect 361757 425579 361823 425582
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580625 418298 580691 418301
rect 583520 418298 584960 418388
rect 580625 418296 584960 418298
rect 580625 418240 580630 418296
rect 580686 418240 584960 418296
rect 580625 418238 584960 418240
rect 580625 418235 580691 418238
rect 583520 418148 584960 418238
rect 361573 414626 361639 414629
rect 359812 414624 361639 414626
rect 359812 414568 361578 414624
rect 361634 414568 361639 414624
rect 359812 414566 361639 414568
rect 361573 414563 361639 414566
rect -960 410546 480 410636
rect 3969 410546 4035 410549
rect -960 410544 4035 410546
rect -960 410488 3974 410544
rect 4030 410488 4035 410544
rect -960 410486 4035 410488
rect -960 410396 480 410486
rect 3969 410483 4035 410486
rect 580717 404970 580783 404973
rect 583520 404970 584960 405060
rect 580717 404968 584960 404970
rect 580717 404912 580722 404968
rect 580778 404912 584960 404968
rect 580717 404910 584960 404912
rect 580717 404907 580783 404910
rect 583520 404820 584960 404910
rect 361573 403610 361639 403613
rect 359812 403608 361639 403610
rect 359812 403552 361578 403608
rect 361634 403552 361639 403608
rect 359812 403550 361639 403552
rect 361573 403547 361639 403550
rect -960 397490 480 397580
rect 3785 397490 3851 397493
rect -960 397488 3851 397490
rect -960 397432 3790 397488
rect 3846 397432 3851 397488
rect -960 397430 3851 397432
rect -960 397340 480 397430
rect 3785 397427 3851 397430
rect 448278 395252 448284 395316
rect 448348 395314 448354 395316
rect 493317 395314 493383 395317
rect 448348 395312 493383 395314
rect 448348 395256 493322 395312
rect 493378 395256 493383 395312
rect 448348 395254 493383 395256
rect 448348 395252 448354 395254
rect 493317 395251 493383 395254
rect 361573 392594 361639 392597
rect 359812 392592 361639 392594
rect 359812 392536 361578 392592
rect 361634 392536 361639 392592
rect 359812 392534 361639 392536
rect 361573 392531 361639 392534
rect 583520 391628 584960 391868
rect 472157 389060 472223 389061
rect 472157 389058 472204 389060
rect 472112 389056 472204 389058
rect 472112 389000 472162 389056
rect 472112 388998 472204 389000
rect 472157 388996 472204 388998
rect 472268 388996 472274 389060
rect 473629 389058 473695 389061
rect 474406 389058 474412 389060
rect 473629 389056 474412 389058
rect 473629 389000 473634 389056
rect 473690 389000 474412 389056
rect 473629 388998 474412 389000
rect 472157 388995 472223 388996
rect 473629 388995 473695 388998
rect 474406 388996 474412 388998
rect 474476 388996 474482 389060
rect 478822 388996 478828 389060
rect 478892 389058 478898 389060
rect 479517 389058 479583 389061
rect 478892 389056 479583 389058
rect 478892 389000 479522 389056
rect 479578 389000 479583 389056
rect 478892 388998 479583 389000
rect 478892 388996 478898 388998
rect 479517 388995 479583 388998
rect 472014 388860 472020 388924
rect 472084 388922 472090 388924
rect 472893 388922 472959 388925
rect 472084 388920 472959 388922
rect 472084 388864 472898 388920
rect 472954 388864 472959 388920
rect 472084 388862 472959 388864
rect 472084 388860 472090 388862
rect 472893 388859 472959 388862
rect 449065 387018 449131 387021
rect 489310 387018 489316 387020
rect 449065 387016 489316 387018
rect 449065 386960 449070 387016
rect 449126 386960 489316 387016
rect 449065 386958 489316 386960
rect 449065 386955 449131 386958
rect 489310 386956 489316 386958
rect 489380 386956 489386 387020
rect 513281 384706 513347 384709
rect 509956 384704 513347 384706
rect 509956 384648 513286 384704
rect 513342 384648 513347 384704
rect 509956 384646 513347 384648
rect 513281 384643 513347 384646
rect -960 384284 480 384524
rect 512453 384162 512519 384165
rect 509956 384160 512519 384162
rect 509956 384104 512458 384160
rect 512514 384104 512519 384160
rect 509956 384102 512519 384104
rect 512453 384099 512519 384102
rect 447133 383618 447199 383621
rect 512637 383618 512703 383621
rect 447133 383616 450156 383618
rect 447133 383560 447138 383616
rect 447194 383560 450156 383616
rect 447133 383558 450156 383560
rect 509956 383616 512703 383618
rect 509956 383560 512642 383616
rect 512698 383560 512703 383616
rect 509956 383558 512703 383560
rect 447133 383555 447199 383558
rect 512637 383555 512703 383558
rect 513281 383074 513347 383077
rect 509956 383072 513347 383074
rect 509956 383016 513286 383072
rect 513342 383016 513347 383072
rect 509956 383014 513347 383016
rect 513281 383011 513347 383014
rect 447225 382938 447291 382941
rect 447225 382936 450156 382938
rect 447225 382880 447230 382936
rect 447286 382880 450156 382936
rect 447225 382878 450156 382880
rect 447225 382875 447291 382878
rect 512453 382530 512519 382533
rect 509956 382528 512519 382530
rect 509956 382472 512458 382528
rect 512514 382472 512519 382528
rect 509956 382470 512519 382472
rect 512453 382467 512519 382470
rect 447133 382258 447199 382261
rect 447133 382256 450156 382258
rect 447133 382200 447138 382256
rect 447194 382200 450156 382256
rect 447133 382198 450156 382200
rect 447133 382195 447199 382198
rect 513097 381986 513163 381989
rect 509956 381984 513163 381986
rect 509956 381928 513102 381984
rect 513158 381928 513163 381984
rect 509956 381926 513163 381928
rect 513097 381923 513163 381926
rect 361573 381578 361639 381581
rect 359812 381576 361639 381578
rect 359812 381520 361578 381576
rect 361634 381520 361639 381576
rect 359812 381518 361639 381520
rect 361573 381515 361639 381518
rect 447225 381578 447291 381581
rect 447225 381576 450156 381578
rect 447225 381520 447230 381576
rect 447286 381520 450156 381576
rect 447225 381518 450156 381520
rect 447225 381515 447291 381518
rect 512453 381442 512519 381445
rect 509956 381440 512519 381442
rect 509956 381384 512458 381440
rect 512514 381384 512519 381440
rect 509956 381382 512519 381384
rect 512453 381379 512519 381382
rect 447225 380898 447291 380901
rect 513189 380898 513255 380901
rect 447225 380896 450156 380898
rect 447225 380840 447230 380896
rect 447286 380840 450156 380896
rect 447225 380838 450156 380840
rect 509956 380896 513255 380898
rect 509956 380840 513194 380896
rect 513250 380840 513255 380896
rect 509956 380838 513255 380840
rect 447225 380835 447291 380838
rect 513189 380835 513255 380838
rect 513281 380354 513347 380357
rect 509956 380352 513347 380354
rect 509956 380296 513286 380352
rect 513342 380296 513347 380352
rect 509956 380294 513347 380296
rect 513281 380291 513347 380294
rect 447133 380218 447199 380221
rect 447133 380216 450156 380218
rect 447133 380160 447138 380216
rect 447194 380160 450156 380216
rect 447133 380158 450156 380160
rect 447133 380155 447199 380158
rect 512545 379810 512611 379813
rect 509956 379808 512611 379810
rect 509956 379752 512550 379808
rect 512606 379752 512611 379808
rect 509956 379750 512611 379752
rect 512545 379747 512611 379750
rect 447501 379538 447567 379541
rect 447501 379536 450156 379538
rect 447501 379480 447506 379536
rect 447562 379480 450156 379536
rect 447501 379478 450156 379480
rect 447501 379475 447567 379478
rect 512821 379266 512887 379269
rect 509956 379264 512887 379266
rect 509956 379208 512826 379264
rect 512882 379208 512887 379264
rect 509956 379206 512887 379208
rect 512821 379203 512887 379206
rect 447133 378858 447199 378861
rect 447133 378856 450156 378858
rect 447133 378800 447138 378856
rect 447194 378800 450156 378856
rect 447133 378798 450156 378800
rect 447133 378795 447199 378798
rect 513281 378722 513347 378725
rect 509956 378720 513347 378722
rect 509956 378664 513286 378720
rect 513342 378664 513347 378720
rect 509956 378662 513347 378664
rect 513281 378659 513347 378662
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 447317 378178 447383 378181
rect 512269 378178 512335 378181
rect 447317 378176 450156 378178
rect 447317 378120 447322 378176
rect 447378 378120 450156 378176
rect 447317 378118 450156 378120
rect 509956 378176 512335 378178
rect 509956 378120 512274 378176
rect 512330 378120 512335 378176
rect 509956 378118 512335 378120
rect 447317 378115 447383 378118
rect 512269 378115 512335 378118
rect 512085 377634 512151 377637
rect 509956 377632 512151 377634
rect 509956 377576 512090 377632
rect 512146 377576 512151 377632
rect 509956 377574 512151 377576
rect 512085 377571 512151 377574
rect 447133 377498 447199 377501
rect 447133 377496 450156 377498
rect 447133 377440 447138 377496
rect 447194 377440 450156 377496
rect 447133 377438 450156 377440
rect 447133 377435 447199 377438
rect 512821 377090 512887 377093
rect 509956 377088 512887 377090
rect 509956 377032 512826 377088
rect 512882 377032 512887 377088
rect 509956 377030 512887 377032
rect 512821 377027 512887 377030
rect 447225 376818 447291 376821
rect 447225 376816 450156 376818
rect 447225 376760 447230 376816
rect 447286 376760 450156 376816
rect 447225 376758 450156 376760
rect 447225 376755 447291 376758
rect 512177 376546 512243 376549
rect 509956 376544 512243 376546
rect 509956 376488 512182 376544
rect 512238 376488 512243 376544
rect 509956 376486 512243 376488
rect 512177 376483 512243 376486
rect 447133 376138 447199 376141
rect 447133 376136 450156 376138
rect 447133 376080 447138 376136
rect 447194 376080 450156 376136
rect 447133 376078 450156 376080
rect 447133 376075 447199 376078
rect 513281 376002 513347 376005
rect 509956 376000 513347 376002
rect 509956 375944 513286 376000
rect 513342 375944 513347 376000
rect 509956 375942 513347 375944
rect 513281 375939 513347 375942
rect 447225 375458 447291 375461
rect 513281 375458 513347 375461
rect 447225 375456 450156 375458
rect 447225 375400 447230 375456
rect 447286 375400 450156 375456
rect 447225 375398 450156 375400
rect 509956 375456 513347 375458
rect 509956 375400 513286 375456
rect 513342 375400 513347 375456
rect 509956 375398 513347 375400
rect 447225 375395 447291 375398
rect 513281 375395 513347 375398
rect 511993 374914 512059 374917
rect 509956 374912 512059 374914
rect 509956 374856 511998 374912
rect 512054 374856 512059 374912
rect 509956 374854 512059 374856
rect 511993 374851 512059 374854
rect 447133 374778 447199 374781
rect 447133 374776 450156 374778
rect 447133 374720 447138 374776
rect 447194 374720 450156 374776
rect 447133 374718 450156 374720
rect 447133 374715 447199 374718
rect 512085 374370 512151 374373
rect 509956 374368 512151 374370
rect 509956 374312 512090 374368
rect 512146 374312 512151 374368
rect 509956 374310 512151 374312
rect 512085 374307 512151 374310
rect 447225 374098 447291 374101
rect 447225 374096 450156 374098
rect 447225 374040 447230 374096
rect 447286 374040 450156 374096
rect 447225 374038 450156 374040
rect 447225 374035 447291 374038
rect 511993 373826 512059 373829
rect 509956 373824 512059 373826
rect 509956 373768 511998 373824
rect 512054 373768 512059 373824
rect 509956 373766 512059 373768
rect 511993 373763 512059 373766
rect 447133 373418 447199 373421
rect 447133 373416 450156 373418
rect 447133 373360 447138 373416
rect 447194 373360 450156 373416
rect 447133 373358 450156 373360
rect 447133 373355 447199 373358
rect 512453 373282 512519 373285
rect 509956 373280 512519 373282
rect 509956 373224 512458 373280
rect 512514 373224 512519 373280
rect 509956 373222 512519 373224
rect 512453 373219 512519 373222
rect 447225 372738 447291 372741
rect 512085 372738 512151 372741
rect 447225 372736 450156 372738
rect 447225 372680 447230 372736
rect 447286 372680 450156 372736
rect 447225 372678 450156 372680
rect 509956 372736 512151 372738
rect 509956 372680 512090 372736
rect 512146 372680 512151 372736
rect 509956 372678 512151 372680
rect 447225 372675 447291 372678
rect 512085 372675 512151 372678
rect 512453 372194 512519 372197
rect 509956 372192 512519 372194
rect 509956 372136 512458 372192
rect 512514 372136 512519 372192
rect 509956 372134 512519 372136
rect 512453 372131 512519 372134
rect 447133 372058 447199 372061
rect 447133 372056 450156 372058
rect 447133 372000 447138 372056
rect 447194 372000 450156 372056
rect 447133 371998 450156 372000
rect 447133 371995 447199 371998
rect 512085 371650 512151 371653
rect 509956 371648 512151 371650
rect 509956 371592 512090 371648
rect 512146 371592 512151 371648
rect 509956 371590 512151 371592
rect 512085 371587 512151 371590
rect -960 371378 480 371468
rect 3877 371378 3943 371381
rect -960 371376 3943 371378
rect -960 371320 3882 371376
rect 3938 371320 3943 371376
rect -960 371318 3943 371320
rect -960 371228 480 371318
rect 3877 371315 3943 371318
rect 447225 371378 447291 371381
rect 447225 371376 450156 371378
rect 447225 371320 447230 371376
rect 447286 371320 450156 371376
rect 447225 371318 450156 371320
rect 447225 371315 447291 371318
rect 512821 371106 512887 371109
rect 509956 371104 512887 371106
rect 509956 371048 512826 371104
rect 512882 371048 512887 371104
rect 509956 371046 512887 371048
rect 512821 371043 512887 371046
rect 447133 370698 447199 370701
rect 447133 370696 450156 370698
rect 447133 370640 447138 370696
rect 447194 370640 450156 370696
rect 447133 370638 450156 370640
rect 447133 370635 447199 370638
rect 361573 370562 361639 370565
rect 512453 370562 512519 370565
rect 359812 370560 361639 370562
rect 359812 370504 361578 370560
rect 361634 370504 361639 370560
rect 359812 370502 361639 370504
rect 509956 370560 512519 370562
rect 509956 370504 512458 370560
rect 512514 370504 512519 370560
rect 509956 370502 512519 370504
rect 361573 370499 361639 370502
rect 512453 370499 512519 370502
rect 447225 370018 447291 370021
rect 513281 370018 513347 370021
rect 447225 370016 450156 370018
rect 447225 369960 447230 370016
rect 447286 369960 450156 370016
rect 447225 369958 450156 369960
rect 509956 370016 513347 370018
rect 509956 369960 513286 370016
rect 513342 369960 513347 370016
rect 509956 369958 513347 369960
rect 447225 369955 447291 369958
rect 513281 369955 513347 369958
rect 513281 369474 513347 369477
rect 509956 369472 513347 369474
rect 509956 369416 513286 369472
rect 513342 369416 513347 369472
rect 509956 369414 513347 369416
rect 513281 369411 513347 369414
rect 447133 369338 447199 369341
rect 447133 369336 450156 369338
rect 447133 369280 447138 369336
rect 447194 369280 450156 369336
rect 447133 369278 450156 369280
rect 447133 369275 447199 369278
rect 512821 368930 512887 368933
rect 509956 368928 512887 368930
rect 509956 368872 512826 368928
rect 512882 368872 512887 368928
rect 509956 368870 512887 368872
rect 512821 368867 512887 368870
rect 447225 368658 447291 368661
rect 447225 368656 450156 368658
rect 447225 368600 447230 368656
rect 447286 368600 450156 368656
rect 447225 368598 450156 368600
rect 447225 368595 447291 368598
rect 512177 368386 512243 368389
rect 509956 368384 512243 368386
rect 509956 368328 512182 368384
rect 512238 368328 512243 368384
rect 509956 368326 512243 368328
rect 512177 368323 512243 368326
rect 447133 367978 447199 367981
rect 447133 367976 450156 367978
rect 447133 367920 447138 367976
rect 447194 367920 450156 367976
rect 447133 367918 450156 367920
rect 447133 367915 447199 367918
rect 511993 367842 512059 367845
rect 509956 367840 512059 367842
rect 509956 367784 511998 367840
rect 512054 367784 512059 367840
rect 509956 367782 512059 367784
rect 511993 367779 512059 367782
rect 447225 367298 447291 367301
rect 513281 367298 513347 367301
rect 447225 367296 450156 367298
rect 447225 367240 447230 367296
rect 447286 367240 450156 367296
rect 447225 367238 450156 367240
rect 509956 367296 513347 367298
rect 509956 367240 513286 367296
rect 513342 367240 513347 367296
rect 509956 367238 513347 367240
rect 447225 367235 447291 367238
rect 513281 367235 513347 367238
rect 513281 366754 513347 366757
rect 509956 366752 513347 366754
rect 509956 366696 513286 366752
rect 513342 366696 513347 366752
rect 509956 366694 513347 366696
rect 513281 366691 513347 366694
rect 447133 366618 447199 366621
rect 447133 366616 450156 366618
rect 447133 366560 447138 366616
rect 447194 366560 450156 366616
rect 447133 366558 450156 366560
rect 447133 366555 447199 366558
rect 511993 366210 512059 366213
rect 509956 366208 512059 366210
rect 509956 366152 511998 366208
rect 512054 366152 512059 366208
rect 509956 366150 512059 366152
rect 511993 366147 512059 366150
rect 447225 365938 447291 365941
rect 447225 365936 450156 365938
rect 447225 365880 447230 365936
rect 447286 365880 450156 365936
rect 447225 365878 450156 365880
rect 447225 365875 447291 365878
rect 509374 365261 509434 365636
rect 447225 365258 447291 365261
rect 447225 365256 450156 365258
rect 447225 365200 447230 365256
rect 447286 365200 450156 365256
rect 447225 365198 450156 365200
rect 509325 365256 509434 365261
rect 509325 365200 509330 365256
rect 509386 365200 509434 365256
rect 509325 365198 509434 365200
rect 447225 365195 447291 365198
rect 509325 365195 509391 365198
rect 513281 365122 513347 365125
rect 509956 365120 513347 365122
rect 509956 365064 513286 365120
rect 513342 365064 513347 365120
rect 509956 365062 513347 365064
rect 513281 365059 513347 365062
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 447133 364578 447199 364581
rect 512637 364578 512703 364581
rect 447133 364576 450156 364578
rect 447133 364520 447138 364576
rect 447194 364520 450156 364576
rect 447133 364518 450156 364520
rect 509956 364576 512703 364578
rect 509956 364520 512642 364576
rect 512698 364520 512703 364576
rect 509956 364518 512703 364520
rect 447133 364515 447199 364518
rect 512637 364515 512703 364518
rect 447225 363898 447291 363901
rect 447225 363896 450156 363898
rect 447225 363840 447230 363896
rect 447286 363840 450156 363896
rect 447225 363838 450156 363840
rect 447225 363835 447291 363838
rect 509926 363626 509986 364004
rect 513281 363626 513347 363629
rect 509926 363624 513347 363626
rect 509926 363568 513286 363624
rect 513342 363568 513347 363624
rect 509926 363566 513347 363568
rect 513281 363563 513347 363566
rect 512453 363490 512519 363493
rect 509956 363488 512519 363490
rect 509956 363432 512458 363488
rect 512514 363432 512519 363488
rect 509956 363430 512519 363432
rect 512453 363427 512519 363430
rect 447133 363218 447199 363221
rect 447133 363216 450156 363218
rect 447133 363160 447138 363216
rect 447194 363160 450156 363216
rect 447133 363158 450156 363160
rect 447133 363155 447199 363158
rect 513005 362946 513071 362949
rect 509956 362944 513071 362946
rect 509956 362888 513010 362944
rect 513066 362888 513071 362944
rect 509956 362886 513071 362888
rect 513005 362883 513071 362886
rect 447133 362538 447199 362541
rect 447133 362536 450156 362538
rect 447133 362480 447138 362536
rect 447194 362480 450156 362536
rect 447133 362478 450156 362480
rect 447133 362475 447199 362478
rect 511993 362402 512059 362405
rect 509956 362400 512059 362402
rect 509956 362344 511998 362400
rect 512054 362344 512059 362400
rect 509956 362342 512059 362344
rect 511993 362339 512059 362342
rect 447225 361858 447291 361861
rect 512269 361858 512335 361861
rect 447225 361856 450156 361858
rect 447225 361800 447230 361856
rect 447286 361800 450156 361856
rect 447225 361798 450156 361800
rect 509956 361856 512335 361858
rect 509956 361800 512274 361856
rect 512330 361800 512335 361856
rect 509956 361798 512335 361800
rect 447225 361795 447291 361798
rect 512269 361795 512335 361798
rect 513189 361314 513255 361317
rect 509956 361312 513255 361314
rect 509956 361256 513194 361312
rect 513250 361256 513255 361312
rect 509956 361254 513255 361256
rect 513189 361251 513255 361254
rect 447225 361178 447291 361181
rect 447225 361176 450156 361178
rect 447225 361120 447230 361176
rect 447286 361120 450156 361176
rect 447225 361118 450156 361120
rect 447225 361115 447291 361118
rect 512361 360770 512427 360773
rect 509956 360768 512427 360770
rect 509956 360712 512366 360768
rect 512422 360712 512427 360768
rect 509956 360710 512427 360712
rect 512361 360707 512427 360710
rect 447133 360498 447199 360501
rect 447133 360496 450156 360498
rect 447133 360440 447138 360496
rect 447194 360440 450156 360496
rect 447133 360438 450156 360440
rect 447133 360435 447199 360438
rect 512913 360226 512979 360229
rect 509956 360224 512979 360226
rect 509956 360168 512918 360224
rect 512974 360168 512979 360224
rect 509956 360166 512979 360168
rect 512913 360163 512979 360166
rect 447133 359818 447199 359821
rect 447133 359816 450156 359818
rect 447133 359760 447138 359816
rect 447194 359760 450156 359816
rect 447133 359758 450156 359760
rect 447133 359755 447199 359758
rect 512729 359682 512795 359685
rect 509956 359680 512795 359682
rect 509956 359624 512734 359680
rect 512790 359624 512795 359680
rect 509956 359622 512795 359624
rect 512729 359619 512795 359622
rect 362217 359546 362283 359549
rect 359812 359544 362283 359546
rect 359812 359488 362222 359544
rect 362278 359488 362283 359544
rect 359812 359486 362283 359488
rect 362217 359483 362283 359486
rect 447225 359138 447291 359141
rect 510613 359138 510679 359141
rect 447225 359136 450156 359138
rect 447225 359080 447230 359136
rect 447286 359080 450156 359136
rect 447225 359078 450156 359080
rect 509956 359136 510679 359138
rect 509956 359080 510618 359136
rect 510674 359080 510679 359136
rect 509956 359078 510679 359080
rect 447225 359075 447291 359078
rect 510613 359075 510679 359078
rect 512361 358594 512427 358597
rect 509956 358592 512427 358594
rect -960 358458 480 358548
rect 509956 358536 512366 358592
rect 512422 358536 512427 358592
rect 509956 358534 512427 358536
rect 512361 358531 512427 358534
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect -960 358398 3483 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 449801 358458 449867 358461
rect 449801 358456 450156 358458
rect 449801 358400 449806 358456
rect 449862 358400 450156 358456
rect 449801 358398 450156 358400
rect 449801 358395 449867 358398
rect 513281 358050 513347 358053
rect 509956 358048 513347 358050
rect 509956 357992 513286 358048
rect 513342 357992 513347 358048
rect 509956 357990 513347 357992
rect 513281 357987 513347 357990
rect 449617 357778 449683 357781
rect 449617 357776 450156 357778
rect 449617 357720 449622 357776
rect 449678 357720 450156 357776
rect 449617 357718 450156 357720
rect 449617 357715 449683 357718
rect 509509 357642 509575 357645
rect 509509 357640 509618 357642
rect 509509 357584 509514 357640
rect 509570 357584 509618 357640
rect 509509 357579 509618 357584
rect 509558 357476 509618 357579
rect 449065 357098 449131 357101
rect 449065 357096 450156 357098
rect 449065 357040 449070 357096
rect 449126 357040 450156 357096
rect 449065 357038 450156 357040
rect 449065 357035 449131 357038
rect 513281 356962 513347 356965
rect 509956 356960 513347 356962
rect 509956 356904 513286 356960
rect 513342 356904 513347 356960
rect 509956 356902 513347 356904
rect 513281 356899 513347 356902
rect 449525 356418 449591 356421
rect 449525 356416 450156 356418
rect 449525 356360 449530 356416
rect 449586 356360 450156 356416
rect 449525 356358 450156 356360
rect 449525 356355 449591 356358
rect 509374 356149 509434 356388
rect 509374 356144 509483 356149
rect 509374 356088 509422 356144
rect 509478 356088 509483 356144
rect 509374 356086 509483 356088
rect 509417 356083 509483 356086
rect 510797 355874 510863 355877
rect 509956 355872 510863 355874
rect 509956 355816 510802 355872
rect 510858 355816 510863 355872
rect 509956 355814 510863 355816
rect 510797 355811 510863 355814
rect 449709 355738 449775 355741
rect 449709 355736 450156 355738
rect 449709 355680 449714 355736
rect 449770 355680 450156 355736
rect 449709 355678 450156 355680
rect 449709 355675 449775 355678
rect 512453 355330 512519 355333
rect 509956 355328 512519 355330
rect 509956 355272 512458 355328
rect 512514 355272 512519 355328
rect 509956 355270 512519 355272
rect 512453 355267 512519 355270
rect 447869 355058 447935 355061
rect 447869 355056 450156 355058
rect 447869 355000 447874 355056
rect 447930 355000 450156 355056
rect 447869 354998 450156 355000
rect 447869 354995 447935 354998
rect 513281 354786 513347 354789
rect 509956 354784 513347 354786
rect 509956 354728 513286 354784
rect 513342 354728 513347 354784
rect 509956 354726 513347 354728
rect 513281 354723 513347 354726
rect 447409 354378 447475 354381
rect 447409 354376 450156 354378
rect 447409 354320 447414 354376
rect 447470 354320 450156 354376
rect 447409 354318 450156 354320
rect 447409 354315 447475 354318
rect 511993 354242 512059 354245
rect 509956 354240 512059 354242
rect 509956 354184 511998 354240
rect 512054 354184 512059 354240
rect 509956 354182 512059 354184
rect 511993 354179 512059 354182
rect 447593 353698 447659 353701
rect 513281 353698 513347 353701
rect 447593 353696 450156 353698
rect 447593 353640 447598 353696
rect 447654 353640 450156 353696
rect 447593 353638 450156 353640
rect 509956 353696 513347 353698
rect 509956 353640 513286 353696
rect 513342 353640 513347 353696
rect 509956 353638 513347 353640
rect 447593 353635 447659 353638
rect 513281 353635 513347 353638
rect 510705 353154 510771 353157
rect 509956 353152 510771 353154
rect 509956 353096 510710 353152
rect 510766 353096 510771 353152
rect 509956 353094 510771 353096
rect 510705 353091 510771 353094
rect 448145 353018 448211 353021
rect 448145 353016 450156 353018
rect 448145 352960 448150 353016
rect 448206 352960 450156 353016
rect 448145 352958 450156 352960
rect 448145 352955 448211 352958
rect 511993 352610 512059 352613
rect 509956 352608 512059 352610
rect 509956 352552 511998 352608
rect 512054 352552 512059 352608
rect 509956 352550 512059 352552
rect 511993 352547 512059 352550
rect 447961 352338 448027 352341
rect 447961 352336 450156 352338
rect 447961 352280 447966 352336
rect 448022 352280 450156 352336
rect 447961 352278 450156 352280
rect 447961 352275 448027 352278
rect 513281 352066 513347 352069
rect 509956 352064 513347 352066
rect 509956 352008 513286 352064
rect 513342 352008 513347 352064
rect 509956 352006 513347 352008
rect 513281 352003 513347 352006
rect 580809 351930 580875 351933
rect 583520 351930 584960 352020
rect 580809 351928 584960 351930
rect 580809 351872 580814 351928
rect 580870 351872 584960 351928
rect 580809 351870 584960 351872
rect 580809 351867 580875 351870
rect 583520 351780 584960 351870
rect 447317 351658 447383 351661
rect 447317 351656 450156 351658
rect 447317 351600 447322 351656
rect 447378 351600 450156 351656
rect 447317 351598 450156 351600
rect 447317 351595 447383 351598
rect 512637 351522 512703 351525
rect 509956 351520 512703 351522
rect 509956 351464 512642 351520
rect 512698 351464 512703 351520
rect 509956 351462 512703 351464
rect 512637 351459 512703 351462
rect 447133 350978 447199 350981
rect 512545 350978 512611 350981
rect 447133 350976 450156 350978
rect 447133 350920 447138 350976
rect 447194 350920 450156 350976
rect 447133 350918 450156 350920
rect 509956 350976 512611 350978
rect 509956 350920 512550 350976
rect 512606 350920 512611 350976
rect 509956 350918 512611 350920
rect 447133 350915 447199 350918
rect 512545 350915 512611 350918
rect 511993 350434 512059 350437
rect 509956 350432 512059 350434
rect 509956 350376 511998 350432
rect 512054 350376 512059 350432
rect 509956 350374 512059 350376
rect 511993 350371 512059 350374
rect 449801 350298 449867 350301
rect 449801 350296 450156 350298
rect 449801 350240 449806 350296
rect 449862 350240 450156 350296
rect 449801 350238 450156 350240
rect 449801 350235 449867 350238
rect 513281 349890 513347 349893
rect 509956 349888 513347 349890
rect 509956 349832 513286 349888
rect 513342 349832 513347 349888
rect 509956 349830 513347 349832
rect 513281 349827 513347 349830
rect 448329 349618 448395 349621
rect 448329 349616 450156 349618
rect 448329 349560 448334 349616
rect 448390 349560 450156 349616
rect 448329 349558 450156 349560
rect 448329 349555 448395 349558
rect 511993 349346 512059 349349
rect 509956 349344 512059 349346
rect 509956 349288 511998 349344
rect 512054 349288 512059 349344
rect 509956 349286 512059 349288
rect 511993 349283 512059 349286
rect 448237 348938 448303 348941
rect 448237 348936 450156 348938
rect 448237 348880 448242 348936
rect 448298 348880 450156 348936
rect 448237 348878 450156 348880
rect 448237 348875 448303 348878
rect 513281 348802 513347 348805
rect 509956 348800 513347 348802
rect 509956 348744 513286 348800
rect 513342 348744 513347 348800
rect 509956 348742 513347 348744
rect 513281 348739 513347 348742
rect 361757 348530 361823 348533
rect 359812 348528 361823 348530
rect 359812 348472 361762 348528
rect 361818 348472 361823 348528
rect 359812 348470 361823 348472
rect 361757 348467 361823 348470
rect 449341 348258 449407 348261
rect 512913 348258 512979 348261
rect 449341 348256 450156 348258
rect 449341 348200 449346 348256
rect 449402 348200 450156 348256
rect 449341 348198 450156 348200
rect 509956 348256 512979 348258
rect 509956 348200 512918 348256
rect 512974 348200 512979 348256
rect 509956 348198 512979 348200
rect 449341 348195 449407 348198
rect 512913 348195 512979 348198
rect 512545 347714 512611 347717
rect 509956 347712 512611 347714
rect 509956 347656 512550 347712
rect 512606 347656 512611 347712
rect 509956 347654 512611 347656
rect 512545 347651 512611 347654
rect 447133 347578 447199 347581
rect 447133 347576 450156 347578
rect 447133 347520 447138 347576
rect 447194 347520 450156 347576
rect 447133 347518 450156 347520
rect 447133 347515 447199 347518
rect 513281 347170 513347 347173
rect 509956 347168 513347 347170
rect 509956 347112 513286 347168
rect 513342 347112 513347 347168
rect 509956 347110 513347 347112
rect 513281 347107 513347 347110
rect 448973 346898 449039 346901
rect 448973 346896 450156 346898
rect 448973 346840 448978 346896
rect 449034 346840 450156 346896
rect 448973 346838 450156 346840
rect 448973 346835 449039 346838
rect 513281 346626 513347 346629
rect 509956 346624 513347 346626
rect 509956 346568 513286 346624
rect 513342 346568 513347 346624
rect 509956 346566 513347 346568
rect 513281 346563 513347 346566
rect 448278 346156 448284 346220
rect 448348 346218 448354 346220
rect 448348 346158 450156 346218
rect 448348 346156 448354 346158
rect 510889 346082 510955 346085
rect 509956 346080 510955 346082
rect 509956 346024 510894 346080
rect 510950 346024 510955 346080
rect 509956 346022 510955 346024
rect 510889 346019 510955 346022
rect 447961 345538 448027 345541
rect 512545 345538 512611 345541
rect 447961 345536 450156 345538
rect -960 345402 480 345492
rect 447961 345480 447966 345536
rect 448022 345480 450156 345536
rect 447961 345478 450156 345480
rect 509956 345536 512611 345538
rect 509956 345480 512550 345536
rect 512606 345480 512611 345536
rect 509956 345478 512611 345480
rect 447961 345475 448027 345478
rect 512545 345475 512611 345478
rect 3601 345402 3667 345405
rect -960 345400 3667 345402
rect -960 345344 3606 345400
rect 3662 345344 3667 345400
rect -960 345342 3667 345344
rect -960 345252 480 345342
rect 3601 345339 3667 345342
rect 513005 344994 513071 344997
rect 509956 344992 513071 344994
rect 509956 344936 513010 344992
rect 513066 344936 513071 344992
rect 509956 344934 513071 344936
rect 513005 344931 513071 344934
rect 447869 344858 447935 344861
rect 447869 344856 450156 344858
rect 447869 344800 447874 344856
rect 447930 344800 450156 344856
rect 447869 344798 450156 344800
rect 447869 344795 447935 344798
rect 449341 344178 449407 344181
rect 449341 344176 450156 344178
rect 449341 344120 449346 344176
rect 449402 344120 450156 344176
rect 449341 344118 450156 344120
rect 449341 344115 449407 344118
rect 509558 344045 509618 344420
rect 509558 344040 509667 344045
rect 509558 343984 509606 344040
rect 509662 343984 509667 344040
rect 509558 343982 509667 343984
rect 509601 343979 509667 343982
rect 512821 343906 512887 343909
rect 509956 343904 512887 343906
rect 509956 343848 512826 343904
rect 512882 343848 512887 343904
rect 509956 343846 512887 343848
rect 512821 343843 512887 343846
rect 448421 343498 448487 343501
rect 448421 343496 450156 343498
rect 448421 343440 448426 343496
rect 448482 343440 450156 343496
rect 448421 343438 450156 343440
rect 448421 343435 448487 343438
rect 513005 343362 513071 343365
rect 509956 343360 513071 343362
rect 509956 343304 513010 343360
rect 513066 343304 513071 343360
rect 509956 343302 513071 343304
rect 513005 343299 513071 343302
rect 449433 342818 449499 342821
rect 510981 342818 511047 342821
rect 449433 342816 450156 342818
rect 449433 342760 449438 342816
rect 449494 342760 450156 342816
rect 449433 342758 450156 342760
rect 509956 342816 511047 342818
rect 509956 342760 510986 342816
rect 511042 342760 511047 342816
rect 509956 342758 511047 342760
rect 449433 342755 449499 342758
rect 510981 342755 511047 342758
rect 512821 342274 512887 342277
rect 509956 342272 512887 342274
rect 509956 342216 512826 342272
rect 512882 342216 512887 342272
rect 509956 342214 512887 342216
rect 512821 342211 512887 342214
rect 447133 342138 447199 342141
rect 447133 342136 450156 342138
rect 447133 342080 447138 342136
rect 447194 342080 450156 342136
rect 447133 342078 450156 342080
rect 447133 342075 447199 342078
rect 513281 341730 513347 341733
rect 509956 341728 513347 341730
rect 509956 341672 513286 341728
rect 513342 341672 513347 341728
rect 509956 341670 513347 341672
rect 513281 341667 513347 341670
rect 447225 341458 447291 341461
rect 447225 341456 450156 341458
rect 447225 341400 447230 341456
rect 447286 341400 450156 341456
rect 447225 341398 450156 341400
rect 447225 341395 447291 341398
rect 513281 341186 513347 341189
rect 509956 341184 513347 341186
rect 509956 341128 513286 341184
rect 513342 341128 513347 341184
rect 509956 341126 513347 341128
rect 513281 341123 513347 341126
rect 447225 340778 447291 340781
rect 447225 340776 450156 340778
rect 447225 340720 447230 340776
rect 447286 340720 450156 340776
rect 447225 340718 450156 340720
rect 447225 340715 447291 340718
rect 512637 340642 512703 340645
rect 509956 340640 512703 340642
rect 509956 340584 512642 340640
rect 512698 340584 512703 340640
rect 509956 340582 512703 340584
rect 512637 340579 512703 340582
rect 447133 340098 447199 340101
rect 511165 340098 511231 340101
rect 447133 340096 450156 340098
rect 447133 340040 447138 340096
rect 447194 340040 450156 340096
rect 447133 340038 450156 340040
rect 509956 340096 511231 340098
rect 509956 340040 511170 340096
rect 511226 340040 511231 340096
rect 509956 340038 511231 340040
rect 447133 340035 447199 340038
rect 511165 340035 511231 340038
rect 512637 339554 512703 339557
rect 509956 339552 512703 339554
rect 509956 339496 512642 339552
rect 512698 339496 512703 339552
rect 509956 339494 512703 339496
rect 512637 339491 512703 339494
rect 447225 339418 447291 339421
rect 447225 339416 450156 339418
rect 447225 339360 447230 339416
rect 447286 339360 450156 339416
rect 447225 339358 450156 339360
rect 447225 339355 447291 339358
rect 511993 339010 512059 339013
rect 509956 339008 512059 339010
rect 509956 338952 511998 339008
rect 512054 338952 512059 339008
rect 509956 338950 512059 338952
rect 511993 338947 512059 338950
rect 447133 338738 447199 338741
rect 447133 338736 450156 338738
rect 447133 338680 447138 338736
rect 447194 338680 450156 338736
rect 447133 338678 450156 338680
rect 447133 338675 447199 338678
rect 513005 338466 513071 338469
rect 509956 338464 513071 338466
rect 509956 338408 513010 338464
rect 513066 338408 513071 338464
rect 583520 338452 584960 338692
rect 509956 338406 513071 338408
rect 513005 338403 513071 338406
rect 447501 338058 447567 338061
rect 447501 338056 450156 338058
rect 447501 338000 447506 338056
rect 447562 338000 450156 338056
rect 447501 337998 450156 338000
rect 447501 337995 447567 337998
rect 511073 337922 511139 337925
rect 509956 337920 511139 337922
rect 509956 337864 511078 337920
rect 511134 337864 511139 337920
rect 509956 337862 511139 337864
rect 511073 337859 511139 337862
rect 450261 337786 450327 337789
rect 450537 337786 450603 337789
rect 450261 337784 450603 337786
rect 450261 337728 450266 337784
rect 450322 337728 450542 337784
rect 450598 337728 450603 337784
rect 450261 337726 450603 337728
rect 450261 337723 450327 337726
rect 450537 337723 450603 337726
rect 361757 337514 361823 337517
rect 359812 337512 361823 337514
rect 359812 337456 361762 337512
rect 361818 337456 361823 337512
rect 359812 337454 361823 337456
rect 361757 337451 361823 337454
rect 447133 337378 447199 337381
rect 513281 337378 513347 337381
rect 447133 337376 450156 337378
rect 447133 337320 447138 337376
rect 447194 337320 450156 337376
rect 447133 337318 450156 337320
rect 509956 337376 513347 337378
rect 509956 337320 513286 337376
rect 513342 337320 513347 337376
rect 509956 337318 513347 337320
rect 447133 337315 447199 337318
rect 513281 337315 513347 337318
rect 427813 336834 427879 336837
rect 428406 336834 428412 336836
rect 427813 336832 428412 336834
rect 427813 336776 427818 336832
rect 427874 336776 428412 336832
rect 427813 336774 428412 336776
rect 427813 336771 427879 336774
rect 428406 336772 428412 336774
rect 428476 336834 428482 336836
rect 450261 336834 450327 336837
rect 513189 336834 513255 336837
rect 428476 336832 450327 336834
rect 428476 336776 450266 336832
rect 450322 336776 450327 336832
rect 428476 336774 450327 336776
rect 509956 336832 513255 336834
rect 509956 336776 513194 336832
rect 513250 336776 513255 336832
rect 509956 336774 513255 336776
rect 428476 336772 428482 336774
rect 450261 336771 450327 336774
rect 513189 336771 513255 336774
rect 447133 336698 447199 336701
rect 447133 336696 450156 336698
rect 447133 336640 447138 336696
rect 447194 336640 450156 336696
rect 447133 336638 450156 336640
rect 447133 336635 447199 336638
rect 447225 336018 447291 336021
rect 447225 336016 450156 336018
rect 447225 335960 447230 336016
rect 447286 335960 450156 336016
rect 447225 335958 450156 335960
rect 447225 335955 447291 335958
rect 509742 335885 509802 336260
rect 509693 335880 509802 335885
rect 509693 335824 509698 335880
rect 509754 335824 509802 335880
rect 509693 335822 509802 335824
rect 509693 335819 509759 335822
rect 511441 335746 511507 335749
rect 509956 335744 511507 335746
rect 509956 335688 511446 335744
rect 511502 335688 511507 335744
rect 509956 335686 511507 335688
rect 511441 335683 511507 335686
rect 447225 335338 447291 335341
rect 447225 335336 450156 335338
rect 447225 335280 447230 335336
rect 447286 335280 450156 335336
rect 447225 335278 450156 335280
rect 447225 335275 447291 335278
rect 513005 335202 513071 335205
rect 509956 335200 513071 335202
rect 509956 335144 513010 335200
rect 513066 335144 513071 335200
rect 509956 335142 513071 335144
rect 513005 335139 513071 335142
rect 447133 334658 447199 334661
rect 512729 334658 512795 334661
rect 447133 334656 450156 334658
rect 447133 334600 447138 334656
rect 447194 334600 450156 334656
rect 447133 334598 450156 334600
rect 509956 334656 512795 334658
rect 509956 334600 512734 334656
rect 512790 334600 512795 334656
rect 509956 334598 512795 334600
rect 447133 334595 447199 334598
rect 512729 334595 512795 334598
rect 420453 334386 420519 334389
rect 424133 334386 424199 334389
rect 425830 334386 425836 334388
rect 420453 334384 421482 334386
rect 420453 334328 420458 334384
rect 420514 334328 421482 334384
rect 420453 334326 421482 334328
rect 420453 334323 420519 334326
rect 421422 334116 421482 334326
rect 424133 334384 425836 334386
rect 424133 334328 424138 334384
rect 424194 334328 425836 334384
rect 424133 334326 425836 334328
rect 424133 334323 424199 334326
rect 425830 334324 425836 334326
rect 425900 334386 425906 334388
rect 425900 334326 431970 334386
rect 425900 334324 425906 334326
rect 431910 334250 431970 334326
rect 450537 334250 450603 334253
rect 431910 334248 450603 334250
rect 431910 334192 450542 334248
rect 450598 334192 450603 334248
rect 431910 334190 450603 334192
rect 450537 334187 450603 334190
rect 421414 334052 421420 334116
rect 421484 334114 421490 334116
rect 449985 334114 450051 334117
rect 513281 334114 513347 334117
rect 421484 334112 450051 334114
rect 421484 334056 449990 334112
rect 450046 334056 450051 334112
rect 421484 334054 450051 334056
rect 509956 334112 513347 334114
rect 509956 334056 513286 334112
rect 513342 334056 513347 334112
rect 509956 334054 513347 334056
rect 421484 334052 421490 334054
rect 449985 334051 450051 334054
rect 513281 334051 513347 334054
rect 447225 333978 447291 333981
rect 447225 333976 450156 333978
rect 447225 333920 447230 333976
rect 447286 333920 450156 333976
rect 447225 333918 450156 333920
rect 447225 333915 447291 333918
rect 447133 333298 447199 333301
rect 447133 333296 450156 333298
rect 447133 333240 447138 333296
rect 447194 333240 450156 333296
rect 447133 333238 450156 333240
rect 447133 333235 447199 333238
rect 509926 333165 509986 333540
rect 509877 333160 509986 333165
rect 509877 333104 509882 333160
rect 509938 333104 509986 333160
rect 509877 333102 509986 333104
rect 509877 333099 509943 333102
rect 510654 333026 510660 333028
rect 509956 332966 510660 333026
rect 510654 332964 510660 332966
rect 510724 332964 510730 333028
rect 432781 332890 432847 332893
rect 429916 332888 432847 332890
rect 429916 332832 432786 332888
rect 432842 332832 432847 332888
rect 429916 332830 432847 332832
rect 432781 332827 432847 332830
rect 448145 332618 448211 332621
rect 448145 332616 450156 332618
rect 448145 332560 448150 332616
rect 448206 332560 450156 332616
rect 448145 332558 450156 332560
rect 448145 332555 448211 332558
rect 518014 332482 518020 332484
rect -960 332196 480 332436
rect 509956 332422 518020 332482
rect 518014 332420 518020 332422
rect 518084 332420 518090 332484
rect 448329 331938 448395 331941
rect 513189 331938 513255 331941
rect 448329 331936 450156 331938
rect 448329 331880 448334 331936
rect 448390 331880 450156 331936
rect 448329 331878 450156 331880
rect 509956 331936 513255 331938
rect 509956 331880 513194 331936
rect 513250 331880 513255 331936
rect 509956 331878 513255 331880
rect 448329 331875 448395 331878
rect 513189 331875 513255 331878
rect 512637 331394 512703 331397
rect 509956 331392 512703 331394
rect 509956 331336 512642 331392
rect 512698 331336 512703 331392
rect 509956 331334 512703 331336
rect 512637 331331 512703 331334
rect 447777 331258 447843 331261
rect 448421 331258 448487 331261
rect 447777 331256 450156 331258
rect 447777 331200 447782 331256
rect 447838 331200 448426 331256
rect 448482 331200 450156 331256
rect 447777 331198 450156 331200
rect 447777 331195 447843 331198
rect 448421 331195 448487 331198
rect 513465 330850 513531 330853
rect 509956 330848 513531 330850
rect 509956 330792 513470 330848
rect 513526 330792 513531 330848
rect 509956 330790 513531 330792
rect 513465 330787 513531 330790
rect 447225 330578 447291 330581
rect 447685 330578 447751 330581
rect 447225 330576 450156 330578
rect 447225 330520 447230 330576
rect 447286 330520 447690 330576
rect 447746 330520 450156 330576
rect 447225 330518 450156 330520
rect 447225 330515 447291 330518
rect 447685 330515 447751 330518
rect 515070 330306 515076 330308
rect 509956 330246 515076 330306
rect 515070 330244 515076 330246
rect 515140 330244 515146 330308
rect 447409 329898 447475 329901
rect 447409 329896 450156 329898
rect 447409 329840 447414 329896
rect 447470 329840 450156 329896
rect 447409 329838 450156 329840
rect 447409 329835 447475 329838
rect 514886 329762 514892 329764
rect 509956 329702 514892 329762
rect 514886 329700 514892 329702
rect 514956 329700 514962 329764
rect 432689 329218 432755 329221
rect 429916 329216 432755 329218
rect 429916 329160 432694 329216
rect 432750 329160 432755 329216
rect 429916 329158 432755 329160
rect 432689 329155 432755 329158
rect 450126 329082 450186 329188
rect 450670 329156 450676 329220
rect 450740 329156 450746 329220
rect 512637 329218 512703 329221
rect 509956 329216 512703 329218
rect 509956 329160 512642 329216
rect 512698 329160 512703 329216
rect 509956 329158 512703 329160
rect 450678 329082 450738 329156
rect 512637 329155 512703 329158
rect 450126 329022 450738 329082
rect 449893 328946 449959 328949
rect 450126 328946 450186 329022
rect 449893 328944 450186 328946
rect 449893 328888 449898 328944
rect 449954 328888 450186 328944
rect 449893 328886 450186 328888
rect 449893 328883 449959 328886
rect 450445 328676 450511 328677
rect 450445 328674 450492 328676
rect 450404 328672 450492 328674
rect 450404 328616 450450 328672
rect 450404 328614 450492 328616
rect 450445 328612 450492 328614
rect 450556 328612 450562 328676
rect 514150 328674 514156 328676
rect 509956 328614 514156 328674
rect 514150 328612 514156 328614
rect 514220 328612 514226 328676
rect 450445 328611 450554 328612
rect 450494 328508 450554 328611
rect 510153 328130 510219 328133
rect 509956 328128 510219 328130
rect 509956 328072 510158 328128
rect 510214 328072 510219 328128
rect 509956 328070 510219 328072
rect 510153 328067 510219 328070
rect 450261 327994 450327 327997
rect 450261 327992 450370 327994
rect 450261 327936 450266 327992
rect 450322 327936 450370 327992
rect 450261 327931 450370 327936
rect 450310 327828 450370 327931
rect 450537 327314 450603 327317
rect 450494 327312 450603 327314
rect 450494 327256 450542 327312
rect 450598 327256 450603 327312
rect 450494 327251 450603 327256
rect 450494 327148 450554 327251
rect 509926 327178 509986 327556
rect 511809 327178 511875 327181
rect 509926 327176 511875 327178
rect 509926 327120 511814 327176
rect 511870 327120 511875 327176
rect 509926 327118 511875 327120
rect 511809 327115 511875 327118
rect 512913 327042 512979 327045
rect 509956 327040 512979 327042
rect 509956 326984 512918 327040
rect 512974 326984 512979 327040
rect 509956 326982 512979 326984
rect 512913 326979 512979 326982
rect 449985 326634 450051 326637
rect 449985 326632 450186 326634
rect 449985 326576 449990 326632
rect 450046 326576 450186 326632
rect 449985 326574 450186 326576
rect 449985 326571 450051 326574
rect 362217 326498 362283 326501
rect 359812 326496 362283 326498
rect 359812 326440 362222 326496
rect 362278 326440 362283 326496
rect 450126 326468 450186 326574
rect 510286 326498 510292 326500
rect 359812 326438 362283 326440
rect 509956 326438 510292 326498
rect 362217 326435 362283 326438
rect 510286 326436 510292 326438
rect 510356 326436 510362 326500
rect 510838 325954 510844 325956
rect 509956 325894 510844 325954
rect 510838 325892 510844 325894
rect 510908 325892 510914 325956
rect 450678 325549 450738 325788
rect 432597 325546 432663 325549
rect 429916 325544 432663 325546
rect 429916 325488 432602 325544
rect 432658 325488 432663 325544
rect 429916 325486 432663 325488
rect 432597 325483 432663 325486
rect 450629 325544 450738 325549
rect 450629 325488 450634 325544
rect 450690 325488 450738 325544
rect 450629 325486 450738 325488
rect 450629 325483 450695 325486
rect 450169 325274 450235 325277
rect 450169 325272 450554 325274
rect 450169 325216 450174 325272
rect 450230 325216 450554 325272
rect 450169 325214 450554 325216
rect 450169 325211 450235 325214
rect 450494 324869 450554 325214
rect 509374 325005 509434 325380
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 509374 325000 509483 325005
rect 509374 324944 509422 325000
rect 509478 324944 509483 325000
rect 509374 324942 509483 324944
rect 509417 324939 509483 324942
rect 450494 324864 450603 324869
rect 517830 324866 517836 324868
rect 450494 324808 450542 324864
rect 450598 324808 450603 324864
rect 450494 324806 450603 324808
rect 509956 324806 517836 324866
rect 450537 324803 450603 324806
rect 517830 324804 517836 324806
rect 517900 324804 517906 324868
rect 450077 324594 450143 324597
rect 450077 324592 450738 324594
rect 450077 324536 450082 324592
rect 450138 324536 450738 324592
rect 450077 324534 450738 324536
rect 450077 324531 450143 324534
rect 450678 324189 450738 324534
rect 511206 324322 511212 324324
rect 509956 324262 511212 324322
rect 511206 324260 511212 324262
rect 511276 324260 511282 324324
rect 450629 324184 450738 324189
rect 450629 324128 450634 324184
rect 450690 324128 450738 324184
rect 450629 324126 450738 324128
rect 450629 324123 450695 324126
rect 511022 323778 511028 323780
rect 509956 323718 511028 323778
rect 511022 323716 511028 323718
rect 511092 323716 511098 323780
rect 509374 322965 509434 323204
rect 509325 322960 509434 322965
rect 509325 322904 509330 322960
rect 509386 322904 509434 322960
rect 509325 322902 509434 322904
rect 509325 322899 509391 322902
rect 446673 322826 446739 322829
rect 526294 322826 526300 322828
rect 446673 322824 451290 322826
rect 446673 322768 446678 322824
rect 446734 322768 451290 322824
rect 446673 322766 451290 322768
rect 446673 322763 446739 322766
rect 451230 322690 451290 322766
rect 485730 322766 526300 322826
rect 462221 322690 462287 322693
rect 451230 322688 462287 322690
rect 451230 322632 462226 322688
rect 462282 322632 462287 322688
rect 451230 322630 462287 322632
rect 462221 322627 462287 322630
rect 480989 322690 481055 322693
rect 485730 322690 485790 322766
rect 526294 322764 526300 322766
rect 526364 322764 526370 322828
rect 480989 322688 485790 322690
rect 480989 322632 480994 322688
rect 481050 322632 485790 322688
rect 480989 322630 485790 322632
rect 480989 322627 481055 322630
rect 509182 322628 509188 322692
rect 509252 322690 509258 322692
rect 510286 322690 510292 322692
rect 509252 322630 510292 322690
rect 509252 322628 509258 322630
rect 510286 322628 510292 322630
rect 510356 322628 510362 322692
rect 458633 322554 458699 322557
rect 461301 322554 461367 322557
rect 458633 322552 461367 322554
rect 458633 322496 458638 322552
rect 458694 322496 461306 322552
rect 461362 322496 461367 322552
rect 458633 322494 461367 322496
rect 458633 322491 458699 322494
rect 461301 322491 461367 322494
rect 473445 322554 473511 322557
rect 480897 322554 480963 322557
rect 473445 322552 480963 322554
rect 473445 322496 473450 322552
rect 473506 322496 480902 322552
rect 480958 322496 480963 322552
rect 473445 322494 480963 322496
rect 473445 322491 473511 322494
rect 480897 322491 480963 322494
rect 473445 322418 473511 322421
rect 481541 322418 481607 322421
rect 473445 322416 481607 322418
rect 473445 322360 473450 322416
rect 473506 322360 481546 322416
rect 481602 322360 481607 322416
rect 473445 322358 481607 322360
rect 473445 322355 473511 322358
rect 481541 322355 481607 322358
rect 510838 322282 510844 322284
rect 466410 322222 510844 322282
rect 460749 322010 460815 322013
rect 466410 322010 466470 322222
rect 510838 322220 510844 322222
rect 510908 322220 510914 322284
rect 509417 322146 509483 322149
rect 460749 322008 466470 322010
rect 460749 321952 460754 322008
rect 460810 321952 466470 322008
rect 460749 321950 466470 321952
rect 476070 322144 509483 322146
rect 476070 322088 509422 322144
rect 509478 322088 509483 322144
rect 476070 322086 509483 322088
rect 460749 321947 460815 321950
rect 432873 321874 432939 321877
rect 429916 321872 432939 321874
rect 429916 321816 432878 321872
rect 432934 321816 432939 321872
rect 429916 321814 432939 321816
rect 432873 321811 432939 321814
rect 456057 321874 456123 321877
rect 476070 321874 476130 322086
rect 509417 322083 509483 322086
rect 456057 321872 476130 321874
rect 456057 321816 456062 321872
rect 456118 321816 476130 321872
rect 456057 321814 476130 321816
rect 456057 321811 456123 321814
rect 460013 321466 460079 321469
rect 558126 321466 558132 321468
rect 460013 321464 558132 321466
rect 460013 321408 460018 321464
rect 460074 321408 558132 321464
rect 460013 321406 558132 321408
rect 460013 321403 460079 321406
rect 558126 321404 558132 321406
rect 558196 321404 558202 321468
rect 447910 321268 447916 321332
rect 447980 321330 447986 321332
rect 462497 321330 462563 321333
rect 447980 321328 462563 321330
rect 447980 321272 462502 321328
rect 462558 321272 462563 321328
rect 447980 321270 462563 321272
rect 447980 321268 447986 321270
rect 462497 321267 462563 321270
rect 470501 321330 470567 321333
rect 530526 321330 530532 321332
rect 470501 321328 530532 321330
rect 470501 321272 470506 321328
rect 470562 321272 530532 321328
rect 470501 321270 530532 321272
rect 470501 321267 470567 321270
rect 530526 321268 530532 321270
rect 530596 321268 530602 321332
rect 449566 321132 449572 321196
rect 449636 321194 449642 321196
rect 482645 321194 482711 321197
rect 449636 321192 482711 321194
rect 449636 321136 482650 321192
rect 482706 321136 482711 321192
rect 449636 321134 482711 321136
rect 449636 321132 449642 321134
rect 482645 321131 482711 321134
rect 444230 320996 444236 321060
rect 444300 321058 444306 321060
rect 461945 321058 462011 321061
rect 444300 321056 462011 321058
rect 444300 321000 461950 321056
rect 462006 321000 462011 321056
rect 444300 320998 462011 321000
rect 444300 320996 444306 320998
rect 461945 320995 462011 320998
rect 507025 320922 507091 320925
rect 511809 320922 511875 320925
rect 507025 320920 511875 320922
rect 507025 320864 507030 320920
rect 507086 320864 511814 320920
rect 511870 320864 511875 320920
rect 507025 320862 511875 320864
rect 507025 320859 507091 320862
rect 511809 320859 511875 320862
rect 507209 320786 507275 320789
rect 516961 320786 517027 320789
rect 507209 320784 517027 320786
rect 507209 320728 507214 320784
rect 507270 320728 516966 320784
rect 517022 320728 517027 320784
rect 507209 320726 517027 320728
rect 507209 320723 507275 320726
rect 516961 320723 517027 320726
rect 445201 320106 445267 320109
rect 483197 320106 483263 320109
rect 445201 320104 483263 320106
rect 445201 320048 445206 320104
rect 445262 320048 483202 320104
rect 483258 320048 483263 320104
rect 445201 320046 483263 320048
rect 445201 320043 445267 320046
rect 483197 320043 483263 320046
rect 446254 319908 446260 319972
rect 446324 319970 446330 319972
rect 472709 319970 472775 319973
rect 446324 319968 472775 319970
rect 446324 319912 472714 319968
rect 472770 319912 472775 319968
rect 446324 319910 472775 319912
rect 446324 319908 446330 319910
rect 472709 319907 472775 319910
rect 446765 319834 446831 319837
rect 472985 319834 473051 319837
rect 446765 319832 473051 319834
rect 446765 319776 446770 319832
rect 446826 319776 472990 319832
rect 473046 319776 473051 319832
rect 446765 319774 473051 319776
rect 446765 319771 446831 319774
rect 472985 319771 473051 319774
rect 447726 319636 447732 319700
rect 447796 319698 447802 319700
rect 471605 319698 471671 319701
rect 447796 319696 471671 319698
rect 447796 319640 471610 319696
rect 471666 319640 471671 319696
rect 447796 319638 471671 319640
rect 447796 319636 447802 319638
rect 471605 319635 471671 319638
rect 501965 319562 502031 319565
rect 538806 319562 538812 319564
rect 501965 319560 538812 319562
rect 501965 319504 501970 319560
rect 502026 319504 538812 319560
rect 501965 319502 538812 319504
rect 501965 319499 502031 319502
rect 538806 319500 538812 319502
rect 538876 319500 538882 319564
rect 460197 319426 460263 319429
rect 509325 319426 509391 319429
rect 460197 319424 509391 319426
rect -960 319290 480 319380
rect 460197 319368 460202 319424
rect 460258 319368 509330 319424
rect 509386 319368 509391 319424
rect 460197 319366 509391 319368
rect 460197 319363 460263 319366
rect 509325 319363 509391 319366
rect 3969 319290 4035 319293
rect -960 319288 4035 319290
rect -960 319232 3974 319288
rect 4030 319232 4035 319288
rect -960 319230 4035 319232
rect -960 319140 480 319230
rect 3969 319227 4035 319230
rect 432781 318202 432847 318205
rect 429916 318200 432847 318202
rect 429916 318144 432786 318200
rect 432842 318144 432847 318200
rect 429916 318142 432847 318144
rect 432781 318139 432847 318142
rect 496445 318066 496511 318069
rect 542670 318066 542676 318068
rect 496445 318064 542676 318066
rect 496445 318008 496450 318064
rect 496506 318008 542676 318064
rect 496445 318006 542676 318008
rect 496445 318003 496511 318006
rect 542670 318004 542676 318006
rect 542740 318004 542746 318068
rect 361757 315482 361823 315485
rect 359812 315480 361823 315482
rect 359812 315424 361762 315480
rect 361818 315424 361823 315480
rect 359812 315422 361823 315424
rect 361757 315419 361823 315422
rect 432597 314530 432663 314533
rect 429916 314528 432663 314530
rect 429916 314472 432602 314528
rect 432658 314472 432663 314528
rect 429916 314470 432663 314472
rect 432597 314467 432663 314470
rect 503161 313986 503227 313989
rect 538254 313986 538260 313988
rect 503161 313984 538260 313986
rect 503161 313928 503166 313984
rect 503222 313928 538260 313984
rect 503161 313926 538260 313928
rect 503161 313923 503227 313926
rect 538254 313924 538260 313926
rect 538324 313924 538330 313988
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 432045 310858 432111 310861
rect 429916 310856 432111 310858
rect 429916 310800 432050 310856
rect 432106 310800 432111 310856
rect 429916 310798 432111 310800
rect 432045 310795 432111 310798
rect 432689 307186 432755 307189
rect 429916 307184 432755 307186
rect 429916 307128 432694 307184
rect 432750 307128 432755 307184
rect 429916 307126 432755 307128
rect 432689 307123 432755 307126
rect 385677 306914 385743 306917
rect 518014 306914 518020 306916
rect 385677 306912 518020 306914
rect 385677 306856 385682 306912
rect 385738 306856 518020 306912
rect 385677 306854 518020 306856
rect 385677 306851 385743 306854
rect 518014 306852 518020 306854
rect 518084 306852 518090 306916
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 382089 306234 382155 306237
rect 508998 306234 509004 306236
rect 382089 306232 509004 306234
rect 382089 306176 382094 306232
rect 382150 306176 509004 306232
rect 382089 306174 509004 306176
rect 382089 306171 382155 306174
rect 508998 306172 509004 306174
rect 509068 306172 509074 306236
rect 381905 306098 381971 306101
rect 510981 306098 511047 306101
rect 381905 306096 511047 306098
rect 381905 306040 381910 306096
rect 381966 306040 510986 306096
rect 511042 306040 511047 306096
rect 381905 306038 511047 306040
rect 381905 306035 381971 306038
rect 510981 306035 511047 306038
rect 381721 305962 381787 305965
rect 510838 305962 510844 305964
rect 381721 305960 510844 305962
rect 381721 305904 381726 305960
rect 381782 305904 510844 305960
rect 381721 305902 510844 305904
rect 381721 305899 381787 305902
rect 510838 305900 510844 305902
rect 510908 305900 510914 305964
rect 381537 305826 381603 305829
rect 511022 305826 511028 305828
rect 381537 305824 511028 305826
rect 381537 305768 381542 305824
rect 381598 305768 511028 305824
rect 381537 305766 511028 305768
rect 381537 305763 381603 305766
rect 511022 305764 511028 305766
rect 511092 305764 511098 305828
rect 370589 305690 370655 305693
rect 517973 305690 518039 305693
rect 370589 305688 518039 305690
rect 370589 305632 370594 305688
rect 370650 305632 517978 305688
rect 518034 305632 518039 305688
rect 370589 305630 518039 305632
rect 370589 305627 370655 305630
rect 517973 305627 518039 305630
rect 361757 304466 361823 304469
rect 359812 304464 361823 304466
rect 359812 304408 361762 304464
rect 361818 304408 361823 304464
rect 359812 304406 361823 304408
rect 361757 304403 361823 304406
rect 379145 303242 379211 303245
rect 509601 303242 509667 303245
rect 379145 303240 509667 303242
rect 379145 303184 379150 303240
rect 379206 303184 509606 303240
rect 509662 303184 509667 303240
rect 379145 303182 509667 303184
rect 379145 303179 379211 303182
rect 509601 303179 509667 303182
rect 379329 303106 379395 303109
rect 510889 303106 510955 303109
rect 379329 303104 510955 303106
rect 379329 303048 379334 303104
rect 379390 303048 510894 303104
rect 510950 303048 510955 303104
rect 379329 303046 510955 303048
rect 379329 303043 379395 303046
rect 510889 303043 510955 303046
rect 378685 302970 378751 302973
rect 513833 302970 513899 302973
rect 378685 302968 513899 302970
rect 378685 302912 378690 302968
rect 378746 302912 513838 302968
rect 513894 302912 513899 302968
rect 378685 302910 513899 302912
rect 378685 302907 378751 302910
rect 513833 302907 513899 302910
rect 362217 302834 362283 302837
rect 512821 302834 512887 302837
rect 362217 302832 512887 302834
rect 362217 302776 362222 302832
rect 362278 302776 512826 302832
rect 512882 302776 512887 302832
rect 362217 302774 512887 302776
rect 362217 302771 362283 302774
rect 512821 302771 512887 302774
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 362401 297666 362467 297669
rect 510654 297666 510660 297668
rect 362401 297664 510660 297666
rect 362401 297608 362406 297664
rect 362462 297608 510660 297664
rect 362401 297606 510660 297608
rect 362401 297603 362467 297606
rect 510654 297604 510660 297606
rect 510724 297604 510730 297668
rect 365069 297530 365135 297533
rect 514886 297530 514892 297532
rect 365069 297528 514892 297530
rect 365069 297472 365074 297528
rect 365130 297472 514892 297528
rect 365069 297470 514892 297472
rect 365069 297467 365135 297470
rect 514886 297468 514892 297470
rect 514956 297468 514962 297532
rect 365345 297394 365411 297397
rect 517830 297394 517836 297396
rect 365345 297392 517836 297394
rect 365345 297336 365350 297392
rect 365406 297336 517836 297392
rect 365345 297334 517836 297336
rect 365345 297331 365411 297334
rect 517830 297332 517836 297334
rect 517900 297332 517906 297396
rect 371969 294538 372035 294541
rect 514150 294538 514156 294540
rect 371969 294536 514156 294538
rect 371969 294480 371974 294536
rect 372030 294480 514156 294536
rect 371969 294478 514156 294480
rect 371969 294475 372035 294478
rect 514150 294476 514156 294478
rect 514220 294476 514226 294540
rect 361757 293450 361823 293453
rect 359812 293448 361823 293450
rect 359812 293392 361762 293448
rect 361818 293392 361823 293448
rect 359812 293390 361823 293392
rect 361757 293387 361823 293390
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 380433 291818 380499 291821
rect 515070 291818 515076 291820
rect 380433 291816 515076 291818
rect 380433 291760 380438 291816
rect 380494 291760 515076 291816
rect 380433 291758 515076 291760
rect 380433 291755 380499 291758
rect 515070 291756 515076 291758
rect 515140 291756 515146 291820
rect 583520 285276 584960 285516
rect 361757 282434 361823 282437
rect 359812 282432 361823 282434
rect 359812 282376 361762 282432
rect 361818 282376 361823 282432
rect 359812 282374 361823 282376
rect 361757 282371 361823 282374
rect -960 279972 480 280212
rect 579889 272234 579955 272237
rect 583520 272234 584960 272324
rect 579889 272232 584960 272234
rect 579889 272176 579894 272232
rect 579950 272176 584960 272232
rect 579889 272174 584960 272176
rect 579889 272171 579955 272174
rect 583520 272084 584960 272174
rect 361757 271418 361823 271421
rect 359812 271416 361823 271418
rect 359812 271360 361762 271416
rect 361818 271360 361823 271416
rect 359812 271358 361823 271360
rect 361757 271355 361823 271358
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 456793 262714 456859 262717
rect 456793 262712 460092 262714
rect 456793 262656 456798 262712
rect 456854 262656 460092 262712
rect 456793 262654 460092 262656
rect 456793 262651 456859 262654
rect 531405 261082 531471 261085
rect 529828 261080 531471 261082
rect 529828 261024 531410 261080
rect 531466 261024 531471 261080
rect 529828 261022 531471 261024
rect 531405 261019 531471 261022
rect 361757 260402 361823 260405
rect 359812 260400 361823 260402
rect 359812 260344 361762 260400
rect 361818 260344 361823 260400
rect 359812 260342 361823 260344
rect 361757 260339 361823 260342
rect 580349 258906 580415 258909
rect 583520 258906 584960 258996
rect 580349 258904 584960 258906
rect 580349 258848 580354 258904
rect 580410 258848 584960 258904
rect 580349 258846 584960 258848
rect 580349 258843 580415 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3601 254146 3667 254149
rect -960 254144 3667 254146
rect -960 254088 3606 254144
rect 3662 254088 3667 254144
rect -960 254086 3667 254088
rect -960 253996 480 254086
rect 3601 254083 3667 254086
rect 361757 249386 361823 249389
rect 359812 249384 361823 249386
rect 359812 249328 361762 249384
rect 361818 249328 361823 249384
rect 359812 249326 361823 249328
rect 361757 249323 361823 249326
rect 456793 248842 456859 248845
rect 456793 248840 460092 248842
rect 456793 248784 456798 248840
rect 456854 248784 460092 248840
rect 456793 248782 460092 248784
rect 456793 248779 456859 248782
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 531313 243674 531379 243677
rect 529828 243672 531379 243674
rect 529828 243616 531318 243672
rect 531374 243616 531379 243672
rect 529828 243614 531379 243616
rect 531313 243611 531379 243614
rect -960 241090 480 241180
rect 3693 241090 3759 241093
rect -960 241088 3759 241090
rect -960 241032 3698 241088
rect 3754 241032 3759 241088
rect -960 241030 3759 241032
rect -960 240940 480 241030
rect 3693 241027 3759 241030
rect 361757 238370 361823 238373
rect 359812 238368 361823 238370
rect 359812 238312 361762 238368
rect 361818 238312 361823 238368
rect 359812 238310 361823 238312
rect 361757 238307 361823 238310
rect 456793 234970 456859 234973
rect 457805 234970 457871 234973
rect 456793 234968 460092 234970
rect 456793 234912 456798 234968
rect 456854 234912 457810 234968
rect 457866 234912 460092 234968
rect 456793 234910 460092 234912
rect 456793 234907 456859 234910
rect 457805 234907 457871 234910
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 361757 227354 361823 227357
rect 359812 227352 361823 227354
rect 359812 227296 361762 227352
rect 361818 227296 361823 227352
rect 359812 227294 361823 227296
rect 361757 227291 361823 227294
rect 530117 226266 530183 226269
rect 529828 226264 530183 226266
rect 529828 226208 530122 226264
rect 530178 226208 530183 226264
rect 529828 226206 530183 226208
rect 530117 226203 530183 226206
rect 457897 221098 457963 221101
rect 457897 221096 460092 221098
rect 457897 221040 457902 221096
rect 457958 221040 460092 221096
rect 457897 221038 460092 221040
rect 457897 221035 457963 221038
rect 580257 219058 580323 219061
rect 583520 219058 584960 219148
rect 580257 219056 584960 219058
rect 580257 219000 580262 219056
rect 580318 219000 584960 219056
rect 580257 218998 584960 219000
rect 580257 218995 580323 218998
rect 583520 218908 584960 218998
rect 361665 216338 361731 216341
rect 359812 216336 361731 216338
rect 359812 216280 361670 216336
rect 361726 216280 361731 216336
rect 359812 216278 361731 216280
rect 361665 216275 361731 216278
rect -960 214978 480 215068
rect 3785 214978 3851 214981
rect -960 214976 3851 214978
rect -960 214920 3790 214976
rect 3846 214920 3851 214976
rect -960 214918 3851 214920
rect -960 214828 480 214918
rect 3785 214915 3851 214918
rect 529933 209266 529999 209269
rect 529798 209264 529999 209266
rect 529798 209208 529938 209264
rect 529994 209208 529999 209264
rect 529798 209206 529999 209208
rect 529798 208828 529858 209206
rect 529933 209203 529999 209206
rect 460013 207362 460079 207365
rect 460013 207360 460122 207362
rect 460013 207304 460018 207360
rect 460074 207304 460122 207360
rect 460013 207299 460122 207304
rect 460062 207196 460122 207299
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect 361757 205322 361823 205325
rect 359812 205320 361823 205322
rect 359812 205264 361762 205320
rect 361818 205264 361823 205320
rect 359812 205262 361823 205264
rect 361757 205259 361823 205262
rect -960 201922 480 202012
rect 3877 201922 3943 201925
rect -960 201920 3943 201922
rect -960 201864 3882 201920
rect 3938 201864 3943 201920
rect -960 201862 3943 201864
rect -960 201772 480 201862
rect 3877 201859 3943 201862
rect 361757 194306 361823 194309
rect 359812 194304 361823 194306
rect 359812 194248 361762 194304
rect 361818 194248 361823 194304
rect 359812 194246 361823 194248
rect 361757 194243 361823 194246
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3969 188866 4035 188869
rect -960 188864 4035 188866
rect -960 188808 3974 188864
rect 4030 188808 4035 188864
rect -960 188806 4035 188808
rect -960 188716 480 188806
rect 3969 188803 4035 188806
rect 361757 183290 361823 183293
rect 359812 183288 361823 183290
rect 359812 183232 361762 183288
rect 361818 183232 361823 183288
rect 359812 183230 361823 183232
rect 361757 183227 361823 183230
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 361757 172274 361823 172277
rect 359812 172272 361823 172274
rect 359812 172216 361762 172272
rect 361818 172216 361823 172272
rect 359812 172214 361823 172216
rect 361757 172211 361823 172214
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 4061 162890 4127 162893
rect -960 162888 4127 162890
rect -960 162832 4066 162888
rect 4122 162832 4127 162888
rect -960 162830 4127 162832
rect -960 162740 480 162830
rect 4061 162827 4127 162830
rect 421414 162692 421420 162756
rect 421484 162754 421490 162756
rect 421833 162754 421899 162757
rect 425881 162756 425947 162757
rect 425830 162754 425836 162756
rect 421484 162752 421899 162754
rect 421484 162696 421838 162752
rect 421894 162696 421899 162752
rect 421484 162694 421899 162696
rect 425790 162694 425836 162754
rect 425900 162752 425947 162756
rect 425942 162696 425947 162752
rect 421484 162692 421490 162694
rect 421833 162691 421899 162694
rect 425830 162692 425836 162694
rect 425900 162692 425947 162696
rect 428406 162692 428412 162756
rect 428476 162754 428482 162756
rect 428641 162754 428707 162757
rect 428476 162752 428707 162754
rect 428476 162696 428646 162752
rect 428702 162696 428707 162752
rect 428476 162694 428707 162696
rect 428476 162692 428482 162694
rect 425881 162691 425947 162692
rect 428641 162691 428707 162694
rect 361757 161258 361823 161261
rect 359812 161256 361823 161258
rect 359812 161200 361762 161256
rect 361818 161200 361823 161256
rect 359812 161198 361823 161200
rect 361757 161195 361823 161198
rect 451733 158266 451799 158269
rect 449788 158264 451799 158266
rect 449788 158208 451738 158264
rect 451794 158208 451799 158264
rect 449788 158206 451799 158208
rect 451733 158203 451799 158206
rect 451733 156906 451799 156909
rect 449788 156904 451799 156906
rect 449788 156848 451738 156904
rect 451794 156848 451799 156904
rect 449788 156846 451799 156848
rect 451733 156843 451799 156846
rect 451917 155546 451983 155549
rect 449788 155544 451983 155546
rect 449788 155488 451922 155544
rect 451978 155488 451983 155544
rect 449788 155486 451983 155488
rect 451917 155483 451983 155486
rect 451917 154186 451983 154189
rect 449788 154184 451983 154186
rect 449788 154128 451922 154184
rect 451978 154128 451983 154184
rect 449788 154126 451983 154128
rect 451917 154123 451983 154126
rect 452377 152826 452443 152829
rect 449788 152824 452443 152826
rect 449788 152768 452382 152824
rect 452438 152768 452443 152824
rect 449788 152766 452443 152768
rect 452377 152763 452443 152766
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect 452009 151466 452075 151469
rect 449788 151464 452075 151466
rect 449788 151408 452014 151464
rect 452070 151408 452075 151464
rect 449788 151406 452075 151408
rect 452009 151403 452075 151406
rect 361757 150242 361823 150245
rect 359812 150240 361823 150242
rect 359812 150184 361762 150240
rect 361818 150184 361823 150240
rect 359812 150182 361823 150184
rect 361757 150179 361823 150182
rect 452469 150106 452535 150109
rect 449788 150104 452535 150106
rect 449788 150048 452474 150104
rect 452530 150048 452535 150104
rect 449788 150046 452535 150048
rect 452469 150043 452535 150046
rect -960 149834 480 149924
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 452561 148746 452627 148749
rect 449788 148744 452627 148746
rect 449788 148688 452566 148744
rect 452622 148688 452627 148744
rect 449788 148686 452627 148688
rect 452561 148683 452627 148686
rect 451733 147386 451799 147389
rect 449788 147384 451799 147386
rect 449788 147328 451738 147384
rect 451794 147328 451799 147384
rect 449788 147326 451799 147328
rect 451733 147323 451799 147326
rect 452561 146026 452627 146029
rect 449788 146024 452627 146026
rect 449788 145968 452566 146024
rect 452622 145968 452627 146024
rect 449788 145966 452627 145968
rect 452561 145963 452627 145966
rect 451457 144666 451523 144669
rect 449788 144664 451523 144666
rect 449788 144608 451462 144664
rect 451518 144608 451523 144664
rect 449788 144606 451523 144608
rect 451457 144603 451523 144606
rect 452561 143306 452627 143309
rect 449788 143304 452627 143306
rect 449788 143248 452566 143304
rect 452622 143248 452627 143304
rect 449788 143246 452627 143248
rect 452561 143243 452627 143246
rect 452561 141946 452627 141949
rect 449788 141944 452627 141946
rect 449788 141888 452566 141944
rect 452622 141888 452627 141944
rect 449788 141886 452627 141888
rect 452561 141883 452627 141886
rect 452561 140586 452627 140589
rect 449788 140584 452627 140586
rect 449788 140528 452566 140584
rect 452622 140528 452627 140584
rect 449788 140526 452627 140528
rect 452561 140523 452627 140526
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 361757 139226 361823 139229
rect 452561 139226 452627 139229
rect 359812 139224 361823 139226
rect 359812 139168 361762 139224
rect 361818 139168 361823 139224
rect 359812 139166 361823 139168
rect 449788 139224 452627 139226
rect 449788 139168 452566 139224
rect 452622 139168 452627 139224
rect 583520 139212 584960 139302
rect 449788 139166 452627 139168
rect 361757 139163 361823 139166
rect 452561 139163 452627 139166
rect 452561 137866 452627 137869
rect 449788 137864 452627 137866
rect 449788 137808 452566 137864
rect 452622 137808 452627 137864
rect 449788 137806 452627 137808
rect 452561 137803 452627 137806
rect 538806 137804 538812 137868
rect 538876 137866 538882 137868
rect 543273 137866 543339 137869
rect 538876 137864 543339 137866
rect 538876 137808 543278 137864
rect 543334 137808 543339 137864
rect 538876 137806 543339 137808
rect 538876 137804 538882 137806
rect 543273 137803 543339 137806
rect 539317 137730 539383 137733
rect 539317 137728 539426 137730
rect 539317 137672 539322 137728
rect 539378 137672 539426 137728
rect 539317 137667 539426 137672
rect 539366 137428 539426 137667
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 452561 136506 452627 136509
rect 449788 136504 452627 136506
rect 449788 136448 452566 136504
rect 452622 136448 452627 136504
rect 449788 136446 452627 136448
rect 452561 136443 452627 136446
rect 539501 135962 539567 135965
rect 539501 135960 539610 135962
rect 539501 135904 539506 135960
rect 539562 135904 539610 135960
rect 539501 135899 539610 135904
rect 539550 135388 539610 135899
rect 452561 135146 452627 135149
rect 449788 135144 452627 135146
rect 449788 135088 452566 135144
rect 452622 135088 452627 135144
rect 449788 135086 452627 135088
rect 452561 135083 452627 135086
rect 452561 133786 452627 133789
rect 449788 133784 452627 133786
rect 449788 133728 452566 133784
rect 452622 133728 452627 133784
rect 449788 133726 452627 133728
rect 452561 133723 452627 133726
rect 539358 133316 539364 133380
rect 539428 133316 539434 133380
rect 452101 132426 452167 132429
rect 449788 132424 452167 132426
rect 449788 132368 452106 132424
rect 452162 132368 452167 132424
rect 449788 132366 452167 132368
rect 452101 132363 452167 132366
rect 543181 131338 543247 131341
rect 539948 131336 543247 131338
rect 539948 131280 543186 131336
rect 543242 131280 543247 131336
rect 539948 131278 543247 131280
rect 543181 131275 543247 131278
rect 452285 131066 452351 131069
rect 449788 131064 452351 131066
rect 449788 131008 452290 131064
rect 452346 131008 452351 131064
rect 449788 131006 452351 131008
rect 452285 131003 452351 131006
rect 452377 129706 452443 129709
rect 449788 129704 452443 129706
rect 449788 129648 452382 129704
rect 452438 129648 452443 129704
rect 449788 129646 452443 129648
rect 452377 129643 452443 129646
rect 542721 129298 542787 129301
rect 539948 129296 542787 129298
rect 539948 129240 542726 129296
rect 542782 129240 542787 129296
rect 539948 129238 542787 129240
rect 542721 129235 542787 129238
rect 452193 128346 452259 128349
rect 449788 128344 452259 128346
rect 449788 128288 452198 128344
rect 452254 128288 452259 128344
rect 449788 128286 452259 128288
rect 452193 128283 452259 128286
rect 361757 128210 361823 128213
rect 359812 128208 361823 128210
rect 359812 128152 361762 128208
rect 361818 128152 361823 128208
rect 359812 128150 361823 128152
rect 361757 128147 361823 128150
rect 543089 127258 543155 127261
rect 539948 127256 543155 127258
rect 539948 127200 543094 127256
rect 543150 127200 543155 127256
rect 539948 127198 543155 127200
rect 543089 127195 543155 127198
rect 452285 126986 452351 126989
rect 449788 126984 452351 126986
rect 449788 126928 452290 126984
rect 452346 126928 452351 126984
rect 449788 126926 452351 126928
rect 452285 126923 452351 126926
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 451733 125626 451799 125629
rect 449788 125624 451799 125626
rect 449788 125568 451738 125624
rect 451794 125568 451799 125624
rect 449788 125566 451799 125568
rect 451733 125563 451799 125566
rect 543273 125218 543339 125221
rect 539948 125216 543339 125218
rect 539948 125160 543278 125216
rect 543334 125160 543339 125216
rect 539948 125158 543339 125160
rect 543273 125155 543339 125158
rect 452101 124266 452167 124269
rect 449788 124264 452167 124266
rect 449788 124208 452106 124264
rect 452162 124208 452167 124264
rect 449788 124206 452167 124208
rect 452101 124203 452167 124206
rect -960 123572 480 123812
rect 540237 123178 540303 123181
rect 539948 123176 540303 123178
rect 539948 123120 540242 123176
rect 540298 123120 540303 123176
rect 539948 123118 540303 123120
rect 540237 123115 540303 123118
rect 451825 122906 451891 122909
rect 449788 122904 451891 122906
rect 449788 122848 451830 122904
rect 451886 122848 451891 122904
rect 449788 122846 451891 122848
rect 451825 122843 451891 122846
rect 451733 121546 451799 121549
rect 449788 121544 451799 121546
rect 449788 121488 451738 121544
rect 451794 121488 451799 121544
rect 449788 121486 451799 121488
rect 451733 121483 451799 121486
rect 539685 121410 539751 121413
rect 539685 121408 539794 121410
rect 539685 121352 539690 121408
rect 539746 121352 539794 121408
rect 539685 121347 539794 121352
rect 539734 121108 539794 121347
rect 539777 119642 539843 119645
rect 539734 119640 539843 119642
rect 539734 119584 539782 119640
rect 539838 119584 539843 119640
rect 539734 119579 539843 119584
rect 539734 119068 539794 119579
rect 361757 117194 361823 117197
rect 359812 117192 361823 117194
rect 359812 117136 361762 117192
rect 361818 117136 361823 117192
rect 359812 117134 361823 117136
rect 361757 117131 361823 117134
rect 541433 117058 541499 117061
rect 539948 117056 541499 117058
rect 539948 117000 541438 117056
rect 541494 117000 541499 117056
rect 539948 116998 541499 117000
rect 541433 116995 541499 116998
rect 540145 115018 540211 115021
rect 539948 115016 540211 115018
rect 539948 114960 540150 115016
rect 540206 114960 540211 115016
rect 539948 114958 540211 114960
rect 540145 114955 540211 114958
rect 539593 113250 539659 113253
rect 539550 113248 539659 113250
rect 539550 113192 539598 113248
rect 539654 113192 539659 113248
rect 539550 113187 539659 113192
rect 539550 112948 539610 113187
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect 541065 110938 541131 110941
rect 539948 110936 541131 110938
rect 539948 110880 541070 110936
rect 541126 110880 541131 110936
rect 539948 110878 541131 110880
rect 541065 110875 541131 110878
rect -960 110666 480 110756
rect 3366 110666 3372 110668
rect -960 110606 3372 110666
rect -960 110516 480 110606
rect 3366 110604 3372 110606
rect 3436 110604 3442 110668
rect 539918 108765 539978 108868
rect 539918 108760 540027 108765
rect 539918 108704 539966 108760
rect 540022 108704 540027 108760
rect 539918 108702 540027 108704
rect 539961 108699 540027 108702
rect 541341 106858 541407 106861
rect 539948 106856 541407 106858
rect 539948 106800 541346 106856
rect 541402 106800 541407 106856
rect 539948 106798 541407 106800
rect 541341 106795 541407 106798
rect 361757 106178 361823 106181
rect 359812 106176 361823 106178
rect 359812 106120 361762 106176
rect 361818 106120 361823 106176
rect 359812 106118 361823 106120
rect 361757 106115 361823 106118
rect 539918 104682 539978 104788
rect 540053 104682 540119 104685
rect 539918 104680 540119 104682
rect 539918 104624 540058 104680
rect 540114 104624 540119 104680
rect 539918 104622 540119 104624
rect 540053 104619 540119 104622
rect 541249 102778 541315 102781
rect 539948 102776 541315 102778
rect 539948 102720 541254 102776
rect 541310 102720 541315 102776
rect 539948 102718 541315 102720
rect 541249 102715 541315 102718
rect 542905 100738 542971 100741
rect 539948 100736 542971 100738
rect 539948 100680 542910 100736
rect 542966 100680 542971 100736
rect 539948 100678 542971 100680
rect 542905 100675 542971 100678
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 542629 98698 542695 98701
rect 539948 98696 542695 98698
rect 539948 98640 542634 98696
rect 542690 98640 542695 98696
rect 539948 98638 542695 98640
rect 542629 98635 542695 98638
rect -960 97610 480 97700
rect 3550 97610 3556 97612
rect -960 97550 3556 97610
rect -960 97460 480 97550
rect 3550 97548 3556 97550
rect 3620 97548 3626 97612
rect 539869 97202 539935 97205
rect 539869 97200 539978 97202
rect 539869 97144 539874 97200
rect 539930 97144 539978 97200
rect 539869 97139 539978 97144
rect 539918 96628 539978 97139
rect 361757 95162 361823 95165
rect 359812 95160 361823 95162
rect 359812 95104 361762 95160
rect 361818 95104 361823 95160
rect 359812 95102 361823 95104
rect 361757 95099 361823 95102
rect 542813 94618 542879 94621
rect 539948 94616 542879 94618
rect 539948 94560 542818 94616
rect 542874 94560 542879 94616
rect 539948 94558 542879 94560
rect 542813 94555 542879 94558
rect 542537 92578 542603 92581
rect 539948 92576 542603 92578
rect 539948 92520 542542 92576
rect 542598 92520 542603 92576
rect 539948 92518 542603 92520
rect 542537 92515 542603 92518
rect 542445 90538 542511 90541
rect 539948 90536 542511 90538
rect 539948 90480 542450 90536
rect 542506 90480 542511 90536
rect 539948 90478 542511 90480
rect 542445 90475 542511 90478
rect 542997 88498 543063 88501
rect 539948 88496 543063 88498
rect 539948 88440 543002 88496
rect 543058 88440 543063 88496
rect 539948 88438 543063 88440
rect 542997 88435 543063 88438
rect 541157 86458 541223 86461
rect 539948 86456 541223 86458
rect 539948 86400 541162 86456
rect 541218 86400 541223 86456
rect 539948 86398 541223 86400
rect 541157 86395 541223 86398
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 542670 84418 542676 84420
rect 539948 84358 542676 84418
rect 542670 84356 542676 84358
rect 542740 84356 542746 84420
rect 361757 84146 361823 84149
rect 359812 84144 361823 84146
rect 359812 84088 361762 84144
rect 361818 84088 361823 84144
rect 359812 84086 361823 84088
rect 361757 84083 361823 84086
rect 540973 82378 541039 82381
rect 539948 82376 541039 82378
rect 539948 82320 540978 82376
rect 541034 82320 541039 82376
rect 539948 82318 541039 82320
rect 540973 82315 541039 82318
rect 361757 73130 361823 73133
rect 359812 73128 361823 73130
rect 359812 73072 361762 73128
rect 361818 73072 361823 73128
rect 359812 73070 361823 73072
rect 361757 73067 361823 73070
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3141 71634 3207 71637
rect -960 71632 3207 71634
rect -960 71576 3146 71632
rect 3202 71576 3207 71632
rect -960 71574 3207 71576
rect -960 71484 480 71574
rect 3141 71571 3207 71574
rect 460381 67690 460447 67693
rect 460841 67690 460907 67693
rect 460381 67688 460907 67690
rect 460381 67632 460386 67688
rect 460442 67632 460846 67688
rect 460902 67632 460907 67688
rect 460381 67630 460907 67632
rect 460381 67627 460447 67630
rect 460798 67627 460907 67630
rect 460798 67524 460858 67627
rect 361757 62114 361823 62117
rect 359812 62112 361823 62114
rect 359812 62056 361762 62112
rect 361818 62056 361823 62112
rect 359812 62054 361823 62056
rect 361757 62051 361823 62054
rect 20897 59938 20963 59941
rect 21449 59938 21515 59941
rect 20897 59936 21515 59938
rect 20897 59880 20902 59936
rect 20958 59880 21454 59936
rect 21510 59880 21515 59936
rect 20897 59878 21515 59880
rect 20897 59875 20963 59878
rect 21449 59875 21515 59878
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3417 58578 3483 58581
rect -960 58576 3483 58578
rect -960 58520 3422 58576
rect 3478 58520 3483 58576
rect -960 58518 3483 58520
rect -960 58428 480 58518
rect 3417 58515 3483 58518
rect 361757 51098 361823 51101
rect 359812 51096 361823 51098
rect 359812 51040 361762 51096
rect 361818 51040 361823 51096
rect 359812 51038 361823 51040
rect 361757 51035 361823 51038
rect 19241 49602 19307 49605
rect 22134 49602 22140 49604
rect 19241 49600 22140 49602
rect 19241 49544 19246 49600
rect 19302 49544 22140 49600
rect 19241 49542 22140 49544
rect 19241 49539 19307 49542
rect 22134 49540 22140 49542
rect 22204 49540 22210 49604
rect 540605 48922 540671 48925
rect 540605 48920 540714 48922
rect 540605 48864 540610 48920
rect 540666 48864 540714 48920
rect 540605 48859 540714 48864
rect 540654 48348 540714 48859
rect 3550 46820 3556 46884
rect 3620 46882 3626 46884
rect 384665 46882 384731 46885
rect 3620 46880 384731 46882
rect 3620 46824 384670 46880
rect 384726 46824 384731 46880
rect 3620 46822 384731 46824
rect 3620 46820 3626 46822
rect 384665 46819 384731 46822
rect 3366 46684 3372 46748
rect 3436 46746 3442 46748
rect 384389 46746 384455 46749
rect 3436 46744 384455 46746
rect 3436 46688 384394 46744
rect 384450 46688 384455 46744
rect 3436 46686 384455 46688
rect 3436 46684 3442 46686
rect 384389 46683 384455 46686
rect 22134 46548 22140 46612
rect 22204 46610 22210 46612
rect 359457 46610 359523 46613
rect 22204 46608 359523 46610
rect 22204 46552 359462 46608
rect 359518 46552 359523 46608
rect 22204 46550 359523 46552
rect 22204 46548 22210 46550
rect 359457 46547 359523 46550
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 536833 41034 536899 41037
rect 536833 41032 540132 41034
rect 536833 40976 536838 41032
rect 536894 40976 540132 41032
rect 536833 40974 540132 40976
rect 536833 40971 536899 40974
rect 540329 34234 540395 34237
rect 540286 34232 540395 34234
rect 540286 34176 540334 34232
rect 540390 34176 540395 34232
rect 540286 34171 540395 34176
rect 540286 33660 540346 34171
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 8753 4042 8819 4045
rect 362217 4042 362283 4045
rect 8753 4040 362283 4042
rect 8753 3984 8758 4040
rect 8814 3984 362222 4040
rect 362278 3984 362283 4040
rect 8753 3982 362283 3984
rect 8753 3979 8819 3982
rect 362217 3979 362283 3982
rect 13537 3906 13603 3909
rect 371969 3906 372035 3909
rect 13537 3904 372035 3906
rect 13537 3848 13542 3904
rect 13598 3848 371974 3904
rect 372030 3848 372035 3904
rect 13537 3846 372035 3848
rect 13537 3843 13603 3846
rect 371969 3843 372035 3846
rect 9949 3770 10015 3773
rect 385769 3770 385835 3773
rect 9949 3768 385835 3770
rect 9949 3712 9954 3768
rect 10010 3712 385774 3768
rect 385830 3712 385835 3768
rect 9949 3710 385835 3712
rect 9949 3707 10015 3710
rect 385769 3707 385835 3710
rect 2865 3634 2931 3637
rect 381537 3634 381603 3637
rect 2865 3632 381603 3634
rect 2865 3576 2870 3632
rect 2926 3576 381542 3632
rect 381598 3576 381603 3632
rect 2865 3574 381603 3576
rect 2865 3571 2931 3574
rect 381537 3571 381603 3574
rect 1669 3498 1735 3501
rect 381721 3498 381787 3501
rect 1669 3496 381787 3498
rect 1669 3440 1674 3496
rect 1730 3440 381726 3496
rect 381782 3440 381787 3496
rect 1669 3438 381787 3440
rect 1669 3435 1735 3438
rect 381721 3435 381787 3438
rect 565 3362 631 3365
rect 460197 3362 460263 3365
rect 565 3360 460263 3362
rect 565 3304 570 3360
rect 626 3304 460202 3360
rect 460258 3304 460263 3360
rect 565 3302 460263 3304
rect 565 3299 631 3302
rect 460197 3299 460263 3302
rect 17033 3226 17099 3229
rect 365069 3226 365135 3229
rect 17033 3224 365135 3226
rect 17033 3168 17038 3224
rect 17094 3168 365074 3224
rect 365130 3168 365135 3224
rect 17033 3166 365135 3168
rect 17033 3163 17099 3166
rect 365069 3163 365135 3166
<< via3 >>
rect 449572 700436 449636 700500
rect 444236 700300 444300 700364
rect 530532 700300 530596 700364
rect 526300 699756 526364 699820
rect 558132 699756 558196 699820
rect 447732 692004 447796 692068
rect 446260 689284 446324 689348
rect 447916 684252 447980 684316
rect 3556 683300 3620 683364
rect 3740 683164 3804 683228
rect 3372 682756 3436 682820
rect 3740 671196 3804 671260
rect 458036 665212 458100 665276
rect 459140 655692 459204 655756
rect 458956 647668 459020 647732
rect 3556 619108 3620 619172
rect 3372 606052 3436 606116
rect 472020 599524 472084 599588
rect 459140 598164 459204 598228
rect 478828 598164 478892 598228
rect 472204 589868 472268 589932
rect 474412 518060 474476 518124
rect 458036 517516 458100 517580
rect 482692 517576 482756 517580
rect 482692 517520 482742 517576
rect 482742 517520 482756 517576
rect 482692 517516 482756 517520
rect 451044 516700 451108 516764
rect 450492 514320 450556 514384
rect 489316 496844 489380 496908
rect 482692 462844 482756 462908
rect 458956 428436 459020 428500
rect 448284 395252 448348 395316
rect 472204 389056 472268 389060
rect 472204 389000 472218 389056
rect 472218 389000 472268 389056
rect 472204 388996 472268 389000
rect 474412 388996 474476 389060
rect 478828 388996 478892 389060
rect 472020 388860 472084 388924
rect 489316 386956 489380 387020
rect 448284 346156 448348 346220
rect 428412 336772 428476 336836
rect 425836 334324 425900 334388
rect 421420 334052 421484 334116
rect 510660 332964 510724 333028
rect 518020 332420 518084 332484
rect 515076 330244 515140 330308
rect 514892 329700 514956 329764
rect 450676 329156 450740 329220
rect 450492 328672 450556 328676
rect 450492 328616 450506 328672
rect 450506 328616 450556 328672
rect 450492 328612 450556 328616
rect 514156 328612 514220 328676
rect 510292 326436 510356 326500
rect 510844 325892 510908 325956
rect 517836 324804 517900 324868
rect 511212 324260 511276 324324
rect 511028 323716 511092 323780
rect 526300 322764 526364 322828
rect 509188 322628 509252 322692
rect 510292 322628 510356 322692
rect 510844 322220 510908 322284
rect 558132 321404 558196 321468
rect 447916 321268 447980 321332
rect 530532 321268 530596 321332
rect 449572 321132 449636 321196
rect 444236 320996 444300 321060
rect 446260 319908 446324 319972
rect 447732 319636 447796 319700
rect 538812 319500 538876 319564
rect 542676 318004 542740 318068
rect 538260 313924 538324 313988
rect 518020 306852 518084 306916
rect 509004 306172 509068 306236
rect 510844 305900 510908 305964
rect 511028 305764 511092 305828
rect 510660 297604 510724 297668
rect 514892 297468 514956 297532
rect 517836 297332 517900 297396
rect 514156 294476 514220 294540
rect 515076 291756 515140 291820
rect 421420 162692 421484 162756
rect 425836 162752 425900 162756
rect 425836 162696 425886 162752
rect 425886 162696 425900 162752
rect 425836 162692 425900 162696
rect 428412 162692 428476 162756
rect 538812 137804 538876 137868
rect 539364 133316 539428 133380
rect 3372 110604 3436 110668
rect 3556 97548 3620 97612
rect 542676 84356 542740 84420
rect 22140 49540 22204 49604
rect 3556 46820 3620 46884
rect 3372 46684 3436 46748
rect 22140 46548 22204 46612
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 3555 683364 3621 683365
rect 3555 683300 3556 683364
rect 3620 683300 3621 683364
rect 3555 683299 3621 683300
rect 3371 682820 3437 682821
rect 3371 682756 3372 682820
rect 3436 682756 3437 682820
rect 3371 682755 3437 682756
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 3374 606117 3434 682755
rect 3558 619173 3618 683299
rect 3739 683228 3805 683229
rect 3739 683164 3740 683228
rect 3804 683164 3805 683228
rect 3739 683163 3805 683164
rect 3742 671261 3802 683163
rect 3739 671260 3805 671261
rect 3739 671196 3740 671260
rect 3804 671196 3805 671260
rect 3739 671195 3805 671196
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 3555 619172 3621 619173
rect 3555 619108 3556 619172
rect 3620 619108 3621 619172
rect 3555 619107 3621 619108
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 3371 606116 3437 606117
rect 3371 606052 3372 606116
rect 3436 606052 3437 606116
rect 3371 606051 3437 606052
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 3371 110668 3437 110669
rect 3371 110604 3372 110668
rect 3436 110604 3437 110668
rect 3371 110603 3437 110604
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 3374 46749 3434 110603
rect 3555 97612 3621 97613
rect 3555 97548 3556 97612
rect 3620 97548 3621 97612
rect 3555 97547 3621 97548
rect 3558 46885 3618 97547
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 3555 46884 3621 46885
rect 3555 46820 3556 46884
rect 3620 46820 3621 46884
rect 3555 46819 3621 46820
rect 3371 46748 3437 46749
rect 3371 46684 3372 46748
rect 3436 46684 3437 46748
rect 3371 46683 3437 46684
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 16674 630334 17294 665778
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 594334 17294 629778
rect 16674 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 17294 594334
rect 16674 594014 17294 594098
rect 16674 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 17294 594014
rect 16674 558334 17294 593778
rect 16674 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 17294 558334
rect 16674 558014 17294 558098
rect 16674 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 17294 558014
rect 16674 522334 17294 557778
rect 16674 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 17294 522334
rect 16674 522014 17294 522098
rect 16674 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 17294 522014
rect 16674 486334 17294 521778
rect 16674 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 17294 486334
rect 16674 486014 17294 486098
rect 16674 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 17294 486014
rect 16674 450334 17294 485778
rect 16674 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 17294 450334
rect 16674 450014 17294 450098
rect 16674 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 17294 450014
rect 16674 414334 17294 449778
rect 16674 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 17294 414334
rect 16674 414014 17294 414098
rect 16674 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 17294 414014
rect 16674 378334 17294 413778
rect 16674 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 17294 378334
rect 16674 378014 17294 378098
rect 16674 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 17294 378014
rect 16674 342334 17294 377778
rect 16674 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 17294 342334
rect 16674 342014 17294 342098
rect 16674 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 17294 342014
rect 16674 306334 17294 341778
rect 16674 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 17294 306334
rect 16674 306014 17294 306098
rect 16674 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 17294 306014
rect 16674 270334 17294 305778
rect 16674 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 17294 270334
rect 16674 270014 17294 270098
rect 16674 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 17294 270014
rect 16674 234334 17294 269778
rect 16674 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 17294 234334
rect 16674 234014 17294 234098
rect 16674 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 17294 234014
rect 16674 198334 17294 233778
rect 16674 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 17294 198334
rect 16674 198014 17294 198098
rect 16674 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 17294 198014
rect 16674 162334 17294 197778
rect 16674 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 17294 162334
rect 16674 162014 17294 162098
rect 16674 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 17294 162014
rect 16674 126334 17294 161778
rect 16674 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 17294 126334
rect 16674 126014 17294 126098
rect 16674 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 17294 126014
rect 16674 90334 17294 125778
rect 16674 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 17294 90334
rect 16674 90014 17294 90098
rect 16674 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 17294 90014
rect 16674 54334 17294 89778
rect 16674 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 17294 54334
rect 16674 54014 17294 54098
rect 16674 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 17294 54014
rect 16674 18334 17294 53778
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 -4186 17294 17778
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 670054 21014 709082
rect 20394 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 21014 670054
rect 20394 669734 21014 669818
rect 20394 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 21014 669734
rect 20394 634054 21014 669498
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 27834 677494 28454 711002
rect 27834 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 28454 677494
rect 27834 677174 28454 677258
rect 27834 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 28454 677174
rect 24208 651454 24528 651486
rect 24208 651218 24250 651454
rect 24486 651218 24528 651454
rect 24208 651134 24528 651218
rect 24208 650898 24250 651134
rect 24486 650898 24528 651134
rect 24208 650866 24528 650898
rect 20394 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 21014 634054
rect 20394 633734 21014 633818
rect 20394 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 21014 633734
rect 20394 598054 21014 633498
rect 27834 641494 28454 676938
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 674393 38414 686898
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 674393 42134 690618
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 674393 45854 694338
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 674393 49574 698058
rect 63834 711558 64454 711590
rect 63834 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 64454 711558
rect 63834 711238 64454 711322
rect 63834 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 64454 711238
rect 63834 677494 64454 711002
rect 63834 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 64454 677494
rect 63834 677174 64454 677258
rect 63834 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 64454 677174
rect 63834 674393 64454 676938
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 674393 74414 686898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 674393 78134 690618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 674393 81854 694338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 674393 85574 698058
rect 99834 711558 100454 711590
rect 99834 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 100454 711558
rect 99834 711238 100454 711322
rect 99834 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 100454 711238
rect 99834 677494 100454 711002
rect 99834 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 100454 677494
rect 99834 677174 100454 677258
rect 99834 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 100454 677174
rect 99834 674393 100454 676938
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 674393 110414 686898
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 674393 114134 690618
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 674393 117854 694338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 674393 121574 698058
rect 135834 711558 136454 711590
rect 135834 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 136454 711558
rect 135834 711238 136454 711322
rect 135834 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 136454 711238
rect 135834 677494 136454 711002
rect 135834 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 136454 677494
rect 135834 677174 136454 677258
rect 135834 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 136454 677174
rect 135834 674393 136454 676938
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 674393 146414 686898
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 674393 150134 690618
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 674393 153854 694338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 674393 157574 698058
rect 171834 711558 172454 711590
rect 171834 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 172454 711558
rect 171834 711238 172454 711322
rect 171834 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 172454 711238
rect 171834 677494 172454 711002
rect 171834 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 172454 677494
rect 171834 677174 172454 677258
rect 171834 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 172454 677174
rect 171834 674393 172454 676938
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 674393 182414 686898
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 674393 186134 690618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 674393 189854 694338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 684676 193574 698058
rect 207834 711558 208454 711590
rect 207834 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 208454 711558
rect 207834 711238 208454 711322
rect 207834 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 208454 711238
rect 207834 677494 208454 711002
rect 207834 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 208454 677494
rect 207834 677174 208454 677258
rect 207834 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 208454 677174
rect 207834 674393 208454 676938
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 674393 218414 686898
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 674393 222134 690618
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 674393 225854 694338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 674393 229574 698058
rect 243834 711558 244454 711590
rect 243834 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 244454 711558
rect 243834 711238 244454 711322
rect 243834 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 244454 711238
rect 243834 677494 244454 711002
rect 243834 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 244454 677494
rect 243834 677174 244454 677258
rect 243834 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 244454 677174
rect 243834 674393 244454 676938
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 674393 254414 686898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 674393 258134 690618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 674393 261854 694338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 674393 265574 698058
rect 279834 711558 280454 711590
rect 279834 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 280454 711558
rect 279834 711238 280454 711322
rect 279834 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 280454 711238
rect 279834 677494 280454 711002
rect 279834 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 280454 677494
rect 279834 677174 280454 677258
rect 279834 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 280454 677174
rect 279834 674393 280454 676938
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 674393 290414 686898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 674393 294134 690618
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 674393 297854 694338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 684676 301574 698058
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 674393 326414 686898
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 674393 330134 690618
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 674393 333854 694338
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 674393 337574 698058
rect 351834 711558 352454 711590
rect 351834 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 352454 711558
rect 351834 711238 352454 711322
rect 351834 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 352454 711238
rect 351834 677494 352454 711002
rect 351834 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 352454 677494
rect 351834 677174 352454 677258
rect 351834 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 352454 677174
rect 351834 674393 352454 676938
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 39568 655174 39888 655206
rect 39568 654938 39610 655174
rect 39846 654938 39888 655174
rect 39568 654854 39888 654938
rect 39568 654618 39610 654854
rect 39846 654618 39888 654854
rect 39568 654586 39888 654618
rect 70288 655174 70608 655206
rect 70288 654938 70330 655174
rect 70566 654938 70608 655174
rect 70288 654854 70608 654938
rect 70288 654618 70330 654854
rect 70566 654618 70608 654854
rect 70288 654586 70608 654618
rect 101008 655174 101328 655206
rect 101008 654938 101050 655174
rect 101286 654938 101328 655174
rect 101008 654854 101328 654938
rect 101008 654618 101050 654854
rect 101286 654618 101328 654854
rect 101008 654586 101328 654618
rect 131728 655174 132048 655206
rect 131728 654938 131770 655174
rect 132006 654938 132048 655174
rect 131728 654854 132048 654938
rect 131728 654618 131770 654854
rect 132006 654618 132048 654854
rect 131728 654586 132048 654618
rect 162448 655174 162768 655206
rect 162448 654938 162490 655174
rect 162726 654938 162768 655174
rect 162448 654854 162768 654938
rect 162448 654618 162490 654854
rect 162726 654618 162768 654854
rect 162448 654586 162768 654618
rect 193168 655174 193488 655206
rect 193168 654938 193210 655174
rect 193446 654938 193488 655174
rect 193168 654854 193488 654938
rect 193168 654618 193210 654854
rect 193446 654618 193488 654854
rect 193168 654586 193488 654618
rect 223888 655174 224208 655206
rect 223888 654938 223930 655174
rect 224166 654938 224208 655174
rect 223888 654854 224208 654938
rect 223888 654618 223930 654854
rect 224166 654618 224208 654854
rect 223888 654586 224208 654618
rect 254608 655174 254928 655206
rect 254608 654938 254650 655174
rect 254886 654938 254928 655174
rect 254608 654854 254928 654938
rect 254608 654618 254650 654854
rect 254886 654618 254928 654854
rect 254608 654586 254928 654618
rect 285328 655174 285648 655206
rect 285328 654938 285370 655174
rect 285606 654938 285648 655174
rect 285328 654854 285648 654938
rect 285328 654618 285370 654854
rect 285606 654618 285648 654854
rect 285328 654586 285648 654618
rect 316048 655174 316368 655206
rect 316048 654938 316090 655174
rect 316326 654938 316368 655174
rect 316048 654854 316368 654938
rect 316048 654618 316090 654854
rect 316326 654618 316368 654854
rect 316048 654586 316368 654618
rect 346768 655174 347088 655206
rect 346768 654938 346810 655174
rect 347046 654938 347088 655174
rect 346768 654854 347088 654938
rect 346768 654618 346810 654854
rect 347046 654618 347088 654854
rect 346768 654586 347088 654618
rect 54928 651454 55248 651486
rect 54928 651218 54970 651454
rect 55206 651218 55248 651454
rect 54928 651134 55248 651218
rect 54928 650898 54970 651134
rect 55206 650898 55248 651134
rect 54928 650866 55248 650898
rect 85648 651454 85968 651486
rect 85648 651218 85690 651454
rect 85926 651218 85968 651454
rect 85648 651134 85968 651218
rect 85648 650898 85690 651134
rect 85926 650898 85968 651134
rect 85648 650866 85968 650898
rect 116368 651454 116688 651486
rect 116368 651218 116410 651454
rect 116646 651218 116688 651454
rect 116368 651134 116688 651218
rect 116368 650898 116410 651134
rect 116646 650898 116688 651134
rect 116368 650866 116688 650898
rect 147088 651454 147408 651486
rect 147088 651218 147130 651454
rect 147366 651218 147408 651454
rect 147088 651134 147408 651218
rect 147088 650898 147130 651134
rect 147366 650898 147408 651134
rect 147088 650866 147408 650898
rect 177808 651454 178128 651486
rect 177808 651218 177850 651454
rect 178086 651218 178128 651454
rect 177808 651134 178128 651218
rect 177808 650898 177850 651134
rect 178086 650898 178128 651134
rect 177808 650866 178128 650898
rect 208528 651454 208848 651486
rect 208528 651218 208570 651454
rect 208806 651218 208848 651454
rect 208528 651134 208848 651218
rect 208528 650898 208570 651134
rect 208806 650898 208848 651134
rect 208528 650866 208848 650898
rect 239248 651454 239568 651486
rect 239248 651218 239290 651454
rect 239526 651218 239568 651454
rect 239248 651134 239568 651218
rect 239248 650898 239290 651134
rect 239526 650898 239568 651134
rect 239248 650866 239568 650898
rect 269968 651454 270288 651486
rect 269968 651218 270010 651454
rect 270246 651218 270288 651454
rect 269968 651134 270288 651218
rect 269968 650898 270010 651134
rect 270246 650898 270288 651134
rect 269968 650866 270288 650898
rect 300688 651454 301008 651486
rect 300688 651218 300730 651454
rect 300966 651218 301008 651454
rect 300688 651134 301008 651218
rect 300688 650898 300730 651134
rect 300966 650898 301008 651134
rect 300688 650866 301008 650898
rect 331408 651454 331728 651486
rect 331408 651218 331450 651454
rect 331686 651218 331728 651454
rect 331408 651134 331728 651218
rect 331408 650898 331450 651134
rect 331686 650898 331728 651134
rect 331408 650866 331728 650898
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 27834 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 28454 641494
rect 27834 641174 28454 641258
rect 27834 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 28454 641174
rect 24208 615454 24528 615486
rect 24208 615218 24250 615454
rect 24486 615218 24528 615454
rect 24208 615134 24528 615218
rect 24208 614898 24250 615134
rect 24486 614898 24528 615134
rect 24208 614866 24528 614898
rect 20394 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 21014 598054
rect 20394 597734 21014 597818
rect 20394 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 21014 597734
rect 20394 562054 21014 597498
rect 27834 605494 28454 640938
rect 39568 619174 39888 619206
rect 39568 618938 39610 619174
rect 39846 618938 39888 619174
rect 39568 618854 39888 618938
rect 39568 618618 39610 618854
rect 39846 618618 39888 618854
rect 39568 618586 39888 618618
rect 70288 619174 70608 619206
rect 70288 618938 70330 619174
rect 70566 618938 70608 619174
rect 70288 618854 70608 618938
rect 70288 618618 70330 618854
rect 70566 618618 70608 618854
rect 70288 618586 70608 618618
rect 101008 619174 101328 619206
rect 101008 618938 101050 619174
rect 101286 618938 101328 619174
rect 101008 618854 101328 618938
rect 101008 618618 101050 618854
rect 101286 618618 101328 618854
rect 101008 618586 101328 618618
rect 131728 619174 132048 619206
rect 131728 618938 131770 619174
rect 132006 618938 132048 619174
rect 131728 618854 132048 618938
rect 131728 618618 131770 618854
rect 132006 618618 132048 618854
rect 131728 618586 132048 618618
rect 162448 619174 162768 619206
rect 162448 618938 162490 619174
rect 162726 618938 162768 619174
rect 162448 618854 162768 618938
rect 162448 618618 162490 618854
rect 162726 618618 162768 618854
rect 162448 618586 162768 618618
rect 193168 619174 193488 619206
rect 193168 618938 193210 619174
rect 193446 618938 193488 619174
rect 193168 618854 193488 618938
rect 193168 618618 193210 618854
rect 193446 618618 193488 618854
rect 193168 618586 193488 618618
rect 223888 619174 224208 619206
rect 223888 618938 223930 619174
rect 224166 618938 224208 619174
rect 223888 618854 224208 618938
rect 223888 618618 223930 618854
rect 224166 618618 224208 618854
rect 223888 618586 224208 618618
rect 254608 619174 254928 619206
rect 254608 618938 254650 619174
rect 254886 618938 254928 619174
rect 254608 618854 254928 618938
rect 254608 618618 254650 618854
rect 254886 618618 254928 618854
rect 254608 618586 254928 618618
rect 285328 619174 285648 619206
rect 285328 618938 285370 619174
rect 285606 618938 285648 619174
rect 285328 618854 285648 618938
rect 285328 618618 285370 618854
rect 285606 618618 285648 618854
rect 285328 618586 285648 618618
rect 316048 619174 316368 619206
rect 316048 618938 316090 619174
rect 316326 618938 316368 619174
rect 316048 618854 316368 618938
rect 316048 618618 316090 618854
rect 316326 618618 316368 618854
rect 316048 618586 316368 618618
rect 346768 619174 347088 619206
rect 346768 618938 346810 619174
rect 347046 618938 347088 619174
rect 346768 618854 347088 618938
rect 346768 618618 346810 618854
rect 347046 618618 347088 618854
rect 346768 618586 347088 618618
rect 54928 615454 55248 615486
rect 54928 615218 54970 615454
rect 55206 615218 55248 615454
rect 54928 615134 55248 615218
rect 54928 614898 54970 615134
rect 55206 614898 55248 615134
rect 54928 614866 55248 614898
rect 85648 615454 85968 615486
rect 85648 615218 85690 615454
rect 85926 615218 85968 615454
rect 85648 615134 85968 615218
rect 85648 614898 85690 615134
rect 85926 614898 85968 615134
rect 85648 614866 85968 614898
rect 116368 615454 116688 615486
rect 116368 615218 116410 615454
rect 116646 615218 116688 615454
rect 116368 615134 116688 615218
rect 116368 614898 116410 615134
rect 116646 614898 116688 615134
rect 116368 614866 116688 614898
rect 147088 615454 147408 615486
rect 147088 615218 147130 615454
rect 147366 615218 147408 615454
rect 147088 615134 147408 615218
rect 147088 614898 147130 615134
rect 147366 614898 147408 615134
rect 147088 614866 147408 614898
rect 177808 615454 178128 615486
rect 177808 615218 177850 615454
rect 178086 615218 178128 615454
rect 177808 615134 178128 615218
rect 177808 614898 177850 615134
rect 178086 614898 178128 615134
rect 177808 614866 178128 614898
rect 208528 615454 208848 615486
rect 208528 615218 208570 615454
rect 208806 615218 208848 615454
rect 208528 615134 208848 615218
rect 208528 614898 208570 615134
rect 208806 614898 208848 615134
rect 208528 614866 208848 614898
rect 239248 615454 239568 615486
rect 239248 615218 239290 615454
rect 239526 615218 239568 615454
rect 239248 615134 239568 615218
rect 239248 614898 239290 615134
rect 239526 614898 239568 615134
rect 239248 614866 239568 614898
rect 269968 615454 270288 615486
rect 269968 615218 270010 615454
rect 270246 615218 270288 615454
rect 269968 615134 270288 615218
rect 269968 614898 270010 615134
rect 270246 614898 270288 615134
rect 269968 614866 270288 614898
rect 300688 615454 301008 615486
rect 300688 615218 300730 615454
rect 300966 615218 301008 615454
rect 300688 615134 301008 615218
rect 300688 614898 300730 615134
rect 300966 614898 301008 615134
rect 300688 614866 301008 614898
rect 331408 615454 331728 615486
rect 331408 615218 331450 615454
rect 331686 615218 331728 615454
rect 331408 615134 331728 615218
rect 331408 614898 331450 615134
rect 331686 614898 331728 615134
rect 331408 614866 331728 614898
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 27834 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 28454 605494
rect 27834 605174 28454 605258
rect 27834 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 28454 605174
rect 24208 579454 24528 579486
rect 24208 579218 24250 579454
rect 24486 579218 24528 579454
rect 24208 579134 24528 579218
rect 24208 578898 24250 579134
rect 24486 578898 24528 579134
rect 24208 578866 24528 578898
rect 20394 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 21014 562054
rect 20394 561734 21014 561818
rect 20394 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 21014 561734
rect 20394 526054 21014 561498
rect 27834 569494 28454 604938
rect 39568 583174 39888 583206
rect 39568 582938 39610 583174
rect 39846 582938 39888 583174
rect 39568 582854 39888 582938
rect 39568 582618 39610 582854
rect 39846 582618 39888 582854
rect 39568 582586 39888 582618
rect 70288 583174 70608 583206
rect 70288 582938 70330 583174
rect 70566 582938 70608 583174
rect 70288 582854 70608 582938
rect 70288 582618 70330 582854
rect 70566 582618 70608 582854
rect 70288 582586 70608 582618
rect 101008 583174 101328 583206
rect 101008 582938 101050 583174
rect 101286 582938 101328 583174
rect 101008 582854 101328 582938
rect 101008 582618 101050 582854
rect 101286 582618 101328 582854
rect 101008 582586 101328 582618
rect 131728 583174 132048 583206
rect 131728 582938 131770 583174
rect 132006 582938 132048 583174
rect 131728 582854 132048 582938
rect 131728 582618 131770 582854
rect 132006 582618 132048 582854
rect 131728 582586 132048 582618
rect 162448 583174 162768 583206
rect 162448 582938 162490 583174
rect 162726 582938 162768 583174
rect 162448 582854 162768 582938
rect 162448 582618 162490 582854
rect 162726 582618 162768 582854
rect 162448 582586 162768 582618
rect 193168 583174 193488 583206
rect 193168 582938 193210 583174
rect 193446 582938 193488 583174
rect 193168 582854 193488 582938
rect 193168 582618 193210 582854
rect 193446 582618 193488 582854
rect 193168 582586 193488 582618
rect 223888 583174 224208 583206
rect 223888 582938 223930 583174
rect 224166 582938 224208 583174
rect 223888 582854 224208 582938
rect 223888 582618 223930 582854
rect 224166 582618 224208 582854
rect 223888 582586 224208 582618
rect 254608 583174 254928 583206
rect 254608 582938 254650 583174
rect 254886 582938 254928 583174
rect 254608 582854 254928 582938
rect 254608 582618 254650 582854
rect 254886 582618 254928 582854
rect 254608 582586 254928 582618
rect 285328 583174 285648 583206
rect 285328 582938 285370 583174
rect 285606 582938 285648 583174
rect 285328 582854 285648 582938
rect 285328 582618 285370 582854
rect 285606 582618 285648 582854
rect 285328 582586 285648 582618
rect 316048 583174 316368 583206
rect 316048 582938 316090 583174
rect 316326 582938 316368 583174
rect 316048 582854 316368 582938
rect 316048 582618 316090 582854
rect 316326 582618 316368 582854
rect 316048 582586 316368 582618
rect 346768 583174 347088 583206
rect 346768 582938 346810 583174
rect 347046 582938 347088 583174
rect 346768 582854 347088 582938
rect 346768 582618 346810 582854
rect 347046 582618 347088 582854
rect 346768 582586 347088 582618
rect 54928 579454 55248 579486
rect 54928 579218 54970 579454
rect 55206 579218 55248 579454
rect 54928 579134 55248 579218
rect 54928 578898 54970 579134
rect 55206 578898 55248 579134
rect 54928 578866 55248 578898
rect 85648 579454 85968 579486
rect 85648 579218 85690 579454
rect 85926 579218 85968 579454
rect 85648 579134 85968 579218
rect 85648 578898 85690 579134
rect 85926 578898 85968 579134
rect 85648 578866 85968 578898
rect 116368 579454 116688 579486
rect 116368 579218 116410 579454
rect 116646 579218 116688 579454
rect 116368 579134 116688 579218
rect 116368 578898 116410 579134
rect 116646 578898 116688 579134
rect 116368 578866 116688 578898
rect 147088 579454 147408 579486
rect 147088 579218 147130 579454
rect 147366 579218 147408 579454
rect 147088 579134 147408 579218
rect 147088 578898 147130 579134
rect 147366 578898 147408 579134
rect 147088 578866 147408 578898
rect 177808 579454 178128 579486
rect 177808 579218 177850 579454
rect 178086 579218 178128 579454
rect 177808 579134 178128 579218
rect 177808 578898 177850 579134
rect 178086 578898 178128 579134
rect 177808 578866 178128 578898
rect 208528 579454 208848 579486
rect 208528 579218 208570 579454
rect 208806 579218 208848 579454
rect 208528 579134 208848 579218
rect 208528 578898 208570 579134
rect 208806 578898 208848 579134
rect 208528 578866 208848 578898
rect 239248 579454 239568 579486
rect 239248 579218 239290 579454
rect 239526 579218 239568 579454
rect 239248 579134 239568 579218
rect 239248 578898 239290 579134
rect 239526 578898 239568 579134
rect 239248 578866 239568 578898
rect 269968 579454 270288 579486
rect 269968 579218 270010 579454
rect 270246 579218 270288 579454
rect 269968 579134 270288 579218
rect 269968 578898 270010 579134
rect 270246 578898 270288 579134
rect 269968 578866 270288 578898
rect 300688 579454 301008 579486
rect 300688 579218 300730 579454
rect 300966 579218 301008 579454
rect 300688 579134 301008 579218
rect 300688 578898 300730 579134
rect 300966 578898 301008 579134
rect 300688 578866 301008 578898
rect 331408 579454 331728 579486
rect 331408 579218 331450 579454
rect 331686 579218 331728 579454
rect 331408 579134 331728 579218
rect 331408 578898 331450 579134
rect 331686 578898 331728 579134
rect 331408 578866 331728 578898
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 27834 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 28454 569494
rect 27834 569174 28454 569258
rect 27834 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 28454 569174
rect 24208 543454 24528 543486
rect 24208 543218 24250 543454
rect 24486 543218 24528 543454
rect 24208 543134 24528 543218
rect 24208 542898 24250 543134
rect 24486 542898 24528 543134
rect 24208 542866 24528 542898
rect 20394 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 21014 526054
rect 20394 525734 21014 525818
rect 20394 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 21014 525734
rect 20394 490054 21014 525498
rect 27834 533494 28454 568938
rect 39568 547174 39888 547206
rect 39568 546938 39610 547174
rect 39846 546938 39888 547174
rect 39568 546854 39888 546938
rect 39568 546618 39610 546854
rect 39846 546618 39888 546854
rect 39568 546586 39888 546618
rect 70288 547174 70608 547206
rect 70288 546938 70330 547174
rect 70566 546938 70608 547174
rect 70288 546854 70608 546938
rect 70288 546618 70330 546854
rect 70566 546618 70608 546854
rect 70288 546586 70608 546618
rect 101008 547174 101328 547206
rect 101008 546938 101050 547174
rect 101286 546938 101328 547174
rect 101008 546854 101328 546938
rect 101008 546618 101050 546854
rect 101286 546618 101328 546854
rect 101008 546586 101328 546618
rect 131728 547174 132048 547206
rect 131728 546938 131770 547174
rect 132006 546938 132048 547174
rect 131728 546854 132048 546938
rect 131728 546618 131770 546854
rect 132006 546618 132048 546854
rect 131728 546586 132048 546618
rect 162448 547174 162768 547206
rect 162448 546938 162490 547174
rect 162726 546938 162768 547174
rect 162448 546854 162768 546938
rect 162448 546618 162490 546854
rect 162726 546618 162768 546854
rect 162448 546586 162768 546618
rect 193168 547174 193488 547206
rect 193168 546938 193210 547174
rect 193446 546938 193488 547174
rect 193168 546854 193488 546938
rect 193168 546618 193210 546854
rect 193446 546618 193488 546854
rect 193168 546586 193488 546618
rect 223888 547174 224208 547206
rect 223888 546938 223930 547174
rect 224166 546938 224208 547174
rect 223888 546854 224208 546938
rect 223888 546618 223930 546854
rect 224166 546618 224208 546854
rect 223888 546586 224208 546618
rect 254608 547174 254928 547206
rect 254608 546938 254650 547174
rect 254886 546938 254928 547174
rect 254608 546854 254928 546938
rect 254608 546618 254650 546854
rect 254886 546618 254928 546854
rect 254608 546586 254928 546618
rect 285328 547174 285648 547206
rect 285328 546938 285370 547174
rect 285606 546938 285648 547174
rect 285328 546854 285648 546938
rect 285328 546618 285370 546854
rect 285606 546618 285648 546854
rect 285328 546586 285648 546618
rect 316048 547174 316368 547206
rect 316048 546938 316090 547174
rect 316326 546938 316368 547174
rect 316048 546854 316368 546938
rect 316048 546618 316090 546854
rect 316326 546618 316368 546854
rect 316048 546586 316368 546618
rect 346768 547174 347088 547206
rect 346768 546938 346810 547174
rect 347046 546938 347088 547174
rect 346768 546854 347088 546938
rect 346768 546618 346810 546854
rect 347046 546618 347088 546854
rect 346768 546586 347088 546618
rect 54928 543454 55248 543486
rect 54928 543218 54970 543454
rect 55206 543218 55248 543454
rect 54928 543134 55248 543218
rect 54928 542898 54970 543134
rect 55206 542898 55248 543134
rect 54928 542866 55248 542898
rect 85648 543454 85968 543486
rect 85648 543218 85690 543454
rect 85926 543218 85968 543454
rect 85648 543134 85968 543218
rect 85648 542898 85690 543134
rect 85926 542898 85968 543134
rect 85648 542866 85968 542898
rect 116368 543454 116688 543486
rect 116368 543218 116410 543454
rect 116646 543218 116688 543454
rect 116368 543134 116688 543218
rect 116368 542898 116410 543134
rect 116646 542898 116688 543134
rect 116368 542866 116688 542898
rect 147088 543454 147408 543486
rect 147088 543218 147130 543454
rect 147366 543218 147408 543454
rect 147088 543134 147408 543218
rect 147088 542898 147130 543134
rect 147366 542898 147408 543134
rect 147088 542866 147408 542898
rect 177808 543454 178128 543486
rect 177808 543218 177850 543454
rect 178086 543218 178128 543454
rect 177808 543134 178128 543218
rect 177808 542898 177850 543134
rect 178086 542898 178128 543134
rect 177808 542866 178128 542898
rect 208528 543454 208848 543486
rect 208528 543218 208570 543454
rect 208806 543218 208848 543454
rect 208528 543134 208848 543218
rect 208528 542898 208570 543134
rect 208806 542898 208848 543134
rect 208528 542866 208848 542898
rect 239248 543454 239568 543486
rect 239248 543218 239290 543454
rect 239526 543218 239568 543454
rect 239248 543134 239568 543218
rect 239248 542898 239290 543134
rect 239526 542898 239568 543134
rect 239248 542866 239568 542898
rect 269968 543454 270288 543486
rect 269968 543218 270010 543454
rect 270246 543218 270288 543454
rect 269968 543134 270288 543218
rect 269968 542898 270010 543134
rect 270246 542898 270288 543134
rect 269968 542866 270288 542898
rect 300688 543454 301008 543486
rect 300688 543218 300730 543454
rect 300966 543218 301008 543454
rect 300688 543134 301008 543218
rect 300688 542898 300730 543134
rect 300966 542898 301008 543134
rect 300688 542866 301008 542898
rect 331408 543454 331728 543486
rect 331408 543218 331450 543454
rect 331686 543218 331728 543454
rect 331408 543134 331728 543218
rect 331408 542898 331450 543134
rect 331686 542898 331728 543134
rect 331408 542866 331728 542898
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 27834 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 28454 533494
rect 27834 533174 28454 533258
rect 27834 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 28454 533174
rect 24208 507454 24528 507486
rect 24208 507218 24250 507454
rect 24486 507218 24528 507454
rect 24208 507134 24528 507218
rect 24208 506898 24250 507134
rect 24486 506898 24528 507134
rect 24208 506866 24528 506898
rect 20394 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 21014 490054
rect 20394 489734 21014 489818
rect 20394 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 21014 489734
rect 20394 454054 21014 489498
rect 27834 497494 28454 532938
rect 39568 511174 39888 511206
rect 39568 510938 39610 511174
rect 39846 510938 39888 511174
rect 39568 510854 39888 510938
rect 39568 510618 39610 510854
rect 39846 510618 39888 510854
rect 39568 510586 39888 510618
rect 70288 511174 70608 511206
rect 70288 510938 70330 511174
rect 70566 510938 70608 511174
rect 70288 510854 70608 510938
rect 70288 510618 70330 510854
rect 70566 510618 70608 510854
rect 70288 510586 70608 510618
rect 101008 511174 101328 511206
rect 101008 510938 101050 511174
rect 101286 510938 101328 511174
rect 101008 510854 101328 510938
rect 101008 510618 101050 510854
rect 101286 510618 101328 510854
rect 101008 510586 101328 510618
rect 131728 511174 132048 511206
rect 131728 510938 131770 511174
rect 132006 510938 132048 511174
rect 131728 510854 132048 510938
rect 131728 510618 131770 510854
rect 132006 510618 132048 510854
rect 131728 510586 132048 510618
rect 162448 511174 162768 511206
rect 162448 510938 162490 511174
rect 162726 510938 162768 511174
rect 162448 510854 162768 510938
rect 162448 510618 162490 510854
rect 162726 510618 162768 510854
rect 162448 510586 162768 510618
rect 193168 511174 193488 511206
rect 193168 510938 193210 511174
rect 193446 510938 193488 511174
rect 193168 510854 193488 510938
rect 193168 510618 193210 510854
rect 193446 510618 193488 510854
rect 193168 510586 193488 510618
rect 223888 511174 224208 511206
rect 223888 510938 223930 511174
rect 224166 510938 224208 511174
rect 223888 510854 224208 510938
rect 223888 510618 223930 510854
rect 224166 510618 224208 510854
rect 223888 510586 224208 510618
rect 254608 511174 254928 511206
rect 254608 510938 254650 511174
rect 254886 510938 254928 511174
rect 254608 510854 254928 510938
rect 254608 510618 254650 510854
rect 254886 510618 254928 510854
rect 254608 510586 254928 510618
rect 285328 511174 285648 511206
rect 285328 510938 285370 511174
rect 285606 510938 285648 511174
rect 285328 510854 285648 510938
rect 285328 510618 285370 510854
rect 285606 510618 285648 510854
rect 285328 510586 285648 510618
rect 316048 511174 316368 511206
rect 316048 510938 316090 511174
rect 316326 510938 316368 511174
rect 316048 510854 316368 510938
rect 316048 510618 316090 510854
rect 316326 510618 316368 510854
rect 316048 510586 316368 510618
rect 346768 511174 347088 511206
rect 346768 510938 346810 511174
rect 347046 510938 347088 511174
rect 346768 510854 347088 510938
rect 346768 510618 346810 510854
rect 347046 510618 347088 510854
rect 346768 510586 347088 510618
rect 54928 507454 55248 507486
rect 54928 507218 54970 507454
rect 55206 507218 55248 507454
rect 54928 507134 55248 507218
rect 54928 506898 54970 507134
rect 55206 506898 55248 507134
rect 54928 506866 55248 506898
rect 85648 507454 85968 507486
rect 85648 507218 85690 507454
rect 85926 507218 85968 507454
rect 85648 507134 85968 507218
rect 85648 506898 85690 507134
rect 85926 506898 85968 507134
rect 85648 506866 85968 506898
rect 116368 507454 116688 507486
rect 116368 507218 116410 507454
rect 116646 507218 116688 507454
rect 116368 507134 116688 507218
rect 116368 506898 116410 507134
rect 116646 506898 116688 507134
rect 116368 506866 116688 506898
rect 147088 507454 147408 507486
rect 147088 507218 147130 507454
rect 147366 507218 147408 507454
rect 147088 507134 147408 507218
rect 147088 506898 147130 507134
rect 147366 506898 147408 507134
rect 147088 506866 147408 506898
rect 177808 507454 178128 507486
rect 177808 507218 177850 507454
rect 178086 507218 178128 507454
rect 177808 507134 178128 507218
rect 177808 506898 177850 507134
rect 178086 506898 178128 507134
rect 177808 506866 178128 506898
rect 208528 507454 208848 507486
rect 208528 507218 208570 507454
rect 208806 507218 208848 507454
rect 208528 507134 208848 507218
rect 208528 506898 208570 507134
rect 208806 506898 208848 507134
rect 208528 506866 208848 506898
rect 239248 507454 239568 507486
rect 239248 507218 239290 507454
rect 239526 507218 239568 507454
rect 239248 507134 239568 507218
rect 239248 506898 239290 507134
rect 239526 506898 239568 507134
rect 239248 506866 239568 506898
rect 269968 507454 270288 507486
rect 269968 507218 270010 507454
rect 270246 507218 270288 507454
rect 269968 507134 270288 507218
rect 269968 506898 270010 507134
rect 270246 506898 270288 507134
rect 269968 506866 270288 506898
rect 300688 507454 301008 507486
rect 300688 507218 300730 507454
rect 300966 507218 301008 507454
rect 300688 507134 301008 507218
rect 300688 506898 300730 507134
rect 300966 506898 301008 507134
rect 300688 506866 301008 506898
rect 331408 507454 331728 507486
rect 331408 507218 331450 507454
rect 331686 507218 331728 507454
rect 331408 507134 331728 507218
rect 331408 506898 331450 507134
rect 331686 506898 331728 507134
rect 331408 506866 331728 506898
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 27834 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 28454 497494
rect 27834 497174 28454 497258
rect 27834 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 28454 497174
rect 24208 471454 24528 471486
rect 24208 471218 24250 471454
rect 24486 471218 24528 471454
rect 24208 471134 24528 471218
rect 24208 470898 24250 471134
rect 24486 470898 24528 471134
rect 24208 470866 24528 470898
rect 20394 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 21014 454054
rect 20394 453734 21014 453818
rect 20394 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 21014 453734
rect 20394 418054 21014 453498
rect 27834 461494 28454 496938
rect 39568 475174 39888 475206
rect 39568 474938 39610 475174
rect 39846 474938 39888 475174
rect 39568 474854 39888 474938
rect 39568 474618 39610 474854
rect 39846 474618 39888 474854
rect 39568 474586 39888 474618
rect 70288 475174 70608 475206
rect 70288 474938 70330 475174
rect 70566 474938 70608 475174
rect 70288 474854 70608 474938
rect 70288 474618 70330 474854
rect 70566 474618 70608 474854
rect 70288 474586 70608 474618
rect 101008 475174 101328 475206
rect 101008 474938 101050 475174
rect 101286 474938 101328 475174
rect 101008 474854 101328 474938
rect 101008 474618 101050 474854
rect 101286 474618 101328 474854
rect 101008 474586 101328 474618
rect 131728 475174 132048 475206
rect 131728 474938 131770 475174
rect 132006 474938 132048 475174
rect 131728 474854 132048 474938
rect 131728 474618 131770 474854
rect 132006 474618 132048 474854
rect 131728 474586 132048 474618
rect 162448 475174 162768 475206
rect 162448 474938 162490 475174
rect 162726 474938 162768 475174
rect 162448 474854 162768 474938
rect 162448 474618 162490 474854
rect 162726 474618 162768 474854
rect 162448 474586 162768 474618
rect 193168 475174 193488 475206
rect 193168 474938 193210 475174
rect 193446 474938 193488 475174
rect 193168 474854 193488 474938
rect 193168 474618 193210 474854
rect 193446 474618 193488 474854
rect 193168 474586 193488 474618
rect 223888 475174 224208 475206
rect 223888 474938 223930 475174
rect 224166 474938 224208 475174
rect 223888 474854 224208 474938
rect 223888 474618 223930 474854
rect 224166 474618 224208 474854
rect 223888 474586 224208 474618
rect 254608 475174 254928 475206
rect 254608 474938 254650 475174
rect 254886 474938 254928 475174
rect 254608 474854 254928 474938
rect 254608 474618 254650 474854
rect 254886 474618 254928 474854
rect 254608 474586 254928 474618
rect 285328 475174 285648 475206
rect 285328 474938 285370 475174
rect 285606 474938 285648 475174
rect 285328 474854 285648 474938
rect 285328 474618 285370 474854
rect 285606 474618 285648 474854
rect 285328 474586 285648 474618
rect 316048 475174 316368 475206
rect 316048 474938 316090 475174
rect 316326 474938 316368 475174
rect 316048 474854 316368 474938
rect 316048 474618 316090 474854
rect 316326 474618 316368 474854
rect 316048 474586 316368 474618
rect 346768 475174 347088 475206
rect 346768 474938 346810 475174
rect 347046 474938 347088 475174
rect 346768 474854 347088 474938
rect 346768 474618 346810 474854
rect 347046 474618 347088 474854
rect 346768 474586 347088 474618
rect 54928 471454 55248 471486
rect 54928 471218 54970 471454
rect 55206 471218 55248 471454
rect 54928 471134 55248 471218
rect 54928 470898 54970 471134
rect 55206 470898 55248 471134
rect 54928 470866 55248 470898
rect 85648 471454 85968 471486
rect 85648 471218 85690 471454
rect 85926 471218 85968 471454
rect 85648 471134 85968 471218
rect 85648 470898 85690 471134
rect 85926 470898 85968 471134
rect 85648 470866 85968 470898
rect 116368 471454 116688 471486
rect 116368 471218 116410 471454
rect 116646 471218 116688 471454
rect 116368 471134 116688 471218
rect 116368 470898 116410 471134
rect 116646 470898 116688 471134
rect 116368 470866 116688 470898
rect 147088 471454 147408 471486
rect 147088 471218 147130 471454
rect 147366 471218 147408 471454
rect 147088 471134 147408 471218
rect 147088 470898 147130 471134
rect 147366 470898 147408 471134
rect 147088 470866 147408 470898
rect 177808 471454 178128 471486
rect 177808 471218 177850 471454
rect 178086 471218 178128 471454
rect 177808 471134 178128 471218
rect 177808 470898 177850 471134
rect 178086 470898 178128 471134
rect 177808 470866 178128 470898
rect 208528 471454 208848 471486
rect 208528 471218 208570 471454
rect 208806 471218 208848 471454
rect 208528 471134 208848 471218
rect 208528 470898 208570 471134
rect 208806 470898 208848 471134
rect 208528 470866 208848 470898
rect 239248 471454 239568 471486
rect 239248 471218 239290 471454
rect 239526 471218 239568 471454
rect 239248 471134 239568 471218
rect 239248 470898 239290 471134
rect 239526 470898 239568 471134
rect 239248 470866 239568 470898
rect 269968 471454 270288 471486
rect 269968 471218 270010 471454
rect 270246 471218 270288 471454
rect 269968 471134 270288 471218
rect 269968 470898 270010 471134
rect 270246 470898 270288 471134
rect 269968 470866 270288 470898
rect 300688 471454 301008 471486
rect 300688 471218 300730 471454
rect 300966 471218 301008 471454
rect 300688 471134 301008 471218
rect 300688 470898 300730 471134
rect 300966 470898 301008 471134
rect 300688 470866 301008 470898
rect 331408 471454 331728 471486
rect 331408 471218 331450 471454
rect 331686 471218 331728 471454
rect 331408 471134 331728 471218
rect 331408 470898 331450 471134
rect 331686 470898 331728 471134
rect 331408 470866 331728 470898
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 27834 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 28454 461494
rect 27834 461174 28454 461258
rect 27834 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 28454 461174
rect 24208 435454 24528 435486
rect 24208 435218 24250 435454
rect 24486 435218 24528 435454
rect 24208 435134 24528 435218
rect 24208 434898 24250 435134
rect 24486 434898 24528 435134
rect 24208 434866 24528 434898
rect 20394 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 21014 418054
rect 20394 417734 21014 417818
rect 20394 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 21014 417734
rect 20394 382054 21014 417498
rect 27834 425494 28454 460938
rect 39568 439174 39888 439206
rect 39568 438938 39610 439174
rect 39846 438938 39888 439174
rect 39568 438854 39888 438938
rect 39568 438618 39610 438854
rect 39846 438618 39888 438854
rect 39568 438586 39888 438618
rect 70288 439174 70608 439206
rect 70288 438938 70330 439174
rect 70566 438938 70608 439174
rect 70288 438854 70608 438938
rect 70288 438618 70330 438854
rect 70566 438618 70608 438854
rect 70288 438586 70608 438618
rect 101008 439174 101328 439206
rect 101008 438938 101050 439174
rect 101286 438938 101328 439174
rect 101008 438854 101328 438938
rect 101008 438618 101050 438854
rect 101286 438618 101328 438854
rect 101008 438586 101328 438618
rect 131728 439174 132048 439206
rect 131728 438938 131770 439174
rect 132006 438938 132048 439174
rect 131728 438854 132048 438938
rect 131728 438618 131770 438854
rect 132006 438618 132048 438854
rect 131728 438586 132048 438618
rect 162448 439174 162768 439206
rect 162448 438938 162490 439174
rect 162726 438938 162768 439174
rect 162448 438854 162768 438938
rect 162448 438618 162490 438854
rect 162726 438618 162768 438854
rect 162448 438586 162768 438618
rect 193168 439174 193488 439206
rect 193168 438938 193210 439174
rect 193446 438938 193488 439174
rect 193168 438854 193488 438938
rect 193168 438618 193210 438854
rect 193446 438618 193488 438854
rect 193168 438586 193488 438618
rect 223888 439174 224208 439206
rect 223888 438938 223930 439174
rect 224166 438938 224208 439174
rect 223888 438854 224208 438938
rect 223888 438618 223930 438854
rect 224166 438618 224208 438854
rect 223888 438586 224208 438618
rect 254608 439174 254928 439206
rect 254608 438938 254650 439174
rect 254886 438938 254928 439174
rect 254608 438854 254928 438938
rect 254608 438618 254650 438854
rect 254886 438618 254928 438854
rect 254608 438586 254928 438618
rect 285328 439174 285648 439206
rect 285328 438938 285370 439174
rect 285606 438938 285648 439174
rect 285328 438854 285648 438938
rect 285328 438618 285370 438854
rect 285606 438618 285648 438854
rect 285328 438586 285648 438618
rect 316048 439174 316368 439206
rect 316048 438938 316090 439174
rect 316326 438938 316368 439174
rect 316048 438854 316368 438938
rect 316048 438618 316090 438854
rect 316326 438618 316368 438854
rect 316048 438586 316368 438618
rect 346768 439174 347088 439206
rect 346768 438938 346810 439174
rect 347046 438938 347088 439174
rect 346768 438854 347088 438938
rect 346768 438618 346810 438854
rect 347046 438618 347088 438854
rect 346768 438586 347088 438618
rect 54928 435454 55248 435486
rect 54928 435218 54970 435454
rect 55206 435218 55248 435454
rect 54928 435134 55248 435218
rect 54928 434898 54970 435134
rect 55206 434898 55248 435134
rect 54928 434866 55248 434898
rect 85648 435454 85968 435486
rect 85648 435218 85690 435454
rect 85926 435218 85968 435454
rect 85648 435134 85968 435218
rect 85648 434898 85690 435134
rect 85926 434898 85968 435134
rect 85648 434866 85968 434898
rect 116368 435454 116688 435486
rect 116368 435218 116410 435454
rect 116646 435218 116688 435454
rect 116368 435134 116688 435218
rect 116368 434898 116410 435134
rect 116646 434898 116688 435134
rect 116368 434866 116688 434898
rect 147088 435454 147408 435486
rect 147088 435218 147130 435454
rect 147366 435218 147408 435454
rect 147088 435134 147408 435218
rect 147088 434898 147130 435134
rect 147366 434898 147408 435134
rect 147088 434866 147408 434898
rect 177808 435454 178128 435486
rect 177808 435218 177850 435454
rect 178086 435218 178128 435454
rect 177808 435134 178128 435218
rect 177808 434898 177850 435134
rect 178086 434898 178128 435134
rect 177808 434866 178128 434898
rect 208528 435454 208848 435486
rect 208528 435218 208570 435454
rect 208806 435218 208848 435454
rect 208528 435134 208848 435218
rect 208528 434898 208570 435134
rect 208806 434898 208848 435134
rect 208528 434866 208848 434898
rect 239248 435454 239568 435486
rect 239248 435218 239290 435454
rect 239526 435218 239568 435454
rect 239248 435134 239568 435218
rect 239248 434898 239290 435134
rect 239526 434898 239568 435134
rect 239248 434866 239568 434898
rect 269968 435454 270288 435486
rect 269968 435218 270010 435454
rect 270246 435218 270288 435454
rect 269968 435134 270288 435218
rect 269968 434898 270010 435134
rect 270246 434898 270288 435134
rect 269968 434866 270288 434898
rect 300688 435454 301008 435486
rect 300688 435218 300730 435454
rect 300966 435218 301008 435454
rect 300688 435134 301008 435218
rect 300688 434898 300730 435134
rect 300966 434898 301008 435134
rect 300688 434866 301008 434898
rect 331408 435454 331728 435486
rect 331408 435218 331450 435454
rect 331686 435218 331728 435454
rect 331408 435134 331728 435218
rect 331408 434898 331450 435134
rect 331686 434898 331728 435134
rect 331408 434866 331728 434898
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 27834 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 28454 425494
rect 27834 425174 28454 425258
rect 27834 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 28454 425174
rect 24208 399454 24528 399486
rect 24208 399218 24250 399454
rect 24486 399218 24528 399454
rect 24208 399134 24528 399218
rect 24208 398898 24250 399134
rect 24486 398898 24528 399134
rect 24208 398866 24528 398898
rect 20394 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 21014 382054
rect 20394 381734 21014 381818
rect 20394 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 21014 381734
rect 20394 346054 21014 381498
rect 27834 389494 28454 424938
rect 39568 403174 39888 403206
rect 39568 402938 39610 403174
rect 39846 402938 39888 403174
rect 39568 402854 39888 402938
rect 39568 402618 39610 402854
rect 39846 402618 39888 402854
rect 39568 402586 39888 402618
rect 70288 403174 70608 403206
rect 70288 402938 70330 403174
rect 70566 402938 70608 403174
rect 70288 402854 70608 402938
rect 70288 402618 70330 402854
rect 70566 402618 70608 402854
rect 70288 402586 70608 402618
rect 101008 403174 101328 403206
rect 101008 402938 101050 403174
rect 101286 402938 101328 403174
rect 101008 402854 101328 402938
rect 101008 402618 101050 402854
rect 101286 402618 101328 402854
rect 101008 402586 101328 402618
rect 131728 403174 132048 403206
rect 131728 402938 131770 403174
rect 132006 402938 132048 403174
rect 131728 402854 132048 402938
rect 131728 402618 131770 402854
rect 132006 402618 132048 402854
rect 131728 402586 132048 402618
rect 162448 403174 162768 403206
rect 162448 402938 162490 403174
rect 162726 402938 162768 403174
rect 162448 402854 162768 402938
rect 162448 402618 162490 402854
rect 162726 402618 162768 402854
rect 162448 402586 162768 402618
rect 193168 403174 193488 403206
rect 193168 402938 193210 403174
rect 193446 402938 193488 403174
rect 193168 402854 193488 402938
rect 193168 402618 193210 402854
rect 193446 402618 193488 402854
rect 193168 402586 193488 402618
rect 223888 403174 224208 403206
rect 223888 402938 223930 403174
rect 224166 402938 224208 403174
rect 223888 402854 224208 402938
rect 223888 402618 223930 402854
rect 224166 402618 224208 402854
rect 223888 402586 224208 402618
rect 254608 403174 254928 403206
rect 254608 402938 254650 403174
rect 254886 402938 254928 403174
rect 254608 402854 254928 402938
rect 254608 402618 254650 402854
rect 254886 402618 254928 402854
rect 254608 402586 254928 402618
rect 285328 403174 285648 403206
rect 285328 402938 285370 403174
rect 285606 402938 285648 403174
rect 285328 402854 285648 402938
rect 285328 402618 285370 402854
rect 285606 402618 285648 402854
rect 285328 402586 285648 402618
rect 316048 403174 316368 403206
rect 316048 402938 316090 403174
rect 316326 402938 316368 403174
rect 316048 402854 316368 402938
rect 316048 402618 316090 402854
rect 316326 402618 316368 402854
rect 316048 402586 316368 402618
rect 346768 403174 347088 403206
rect 346768 402938 346810 403174
rect 347046 402938 347088 403174
rect 346768 402854 347088 402938
rect 346768 402618 346810 402854
rect 347046 402618 347088 402854
rect 346768 402586 347088 402618
rect 54928 399454 55248 399486
rect 54928 399218 54970 399454
rect 55206 399218 55248 399454
rect 54928 399134 55248 399218
rect 54928 398898 54970 399134
rect 55206 398898 55248 399134
rect 54928 398866 55248 398898
rect 85648 399454 85968 399486
rect 85648 399218 85690 399454
rect 85926 399218 85968 399454
rect 85648 399134 85968 399218
rect 85648 398898 85690 399134
rect 85926 398898 85968 399134
rect 85648 398866 85968 398898
rect 116368 399454 116688 399486
rect 116368 399218 116410 399454
rect 116646 399218 116688 399454
rect 116368 399134 116688 399218
rect 116368 398898 116410 399134
rect 116646 398898 116688 399134
rect 116368 398866 116688 398898
rect 147088 399454 147408 399486
rect 147088 399218 147130 399454
rect 147366 399218 147408 399454
rect 147088 399134 147408 399218
rect 147088 398898 147130 399134
rect 147366 398898 147408 399134
rect 147088 398866 147408 398898
rect 177808 399454 178128 399486
rect 177808 399218 177850 399454
rect 178086 399218 178128 399454
rect 177808 399134 178128 399218
rect 177808 398898 177850 399134
rect 178086 398898 178128 399134
rect 177808 398866 178128 398898
rect 208528 399454 208848 399486
rect 208528 399218 208570 399454
rect 208806 399218 208848 399454
rect 208528 399134 208848 399218
rect 208528 398898 208570 399134
rect 208806 398898 208848 399134
rect 208528 398866 208848 398898
rect 239248 399454 239568 399486
rect 239248 399218 239290 399454
rect 239526 399218 239568 399454
rect 239248 399134 239568 399218
rect 239248 398898 239290 399134
rect 239526 398898 239568 399134
rect 239248 398866 239568 398898
rect 269968 399454 270288 399486
rect 269968 399218 270010 399454
rect 270246 399218 270288 399454
rect 269968 399134 270288 399218
rect 269968 398898 270010 399134
rect 270246 398898 270288 399134
rect 269968 398866 270288 398898
rect 300688 399454 301008 399486
rect 300688 399218 300730 399454
rect 300966 399218 301008 399454
rect 300688 399134 301008 399218
rect 300688 398898 300730 399134
rect 300966 398898 301008 399134
rect 300688 398866 301008 398898
rect 331408 399454 331728 399486
rect 331408 399218 331450 399454
rect 331686 399218 331728 399454
rect 331408 399134 331728 399218
rect 331408 398898 331450 399134
rect 331686 398898 331728 399134
rect 331408 398866 331728 398898
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 27834 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 28454 389494
rect 27834 389174 28454 389258
rect 27834 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 28454 389174
rect 24208 363454 24528 363486
rect 24208 363218 24250 363454
rect 24486 363218 24528 363454
rect 24208 363134 24528 363218
rect 24208 362898 24250 363134
rect 24486 362898 24528 363134
rect 24208 362866 24528 362898
rect 20394 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 21014 346054
rect 20394 345734 21014 345818
rect 20394 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 21014 345734
rect 20394 310054 21014 345498
rect 27834 353494 28454 388938
rect 39568 367174 39888 367206
rect 39568 366938 39610 367174
rect 39846 366938 39888 367174
rect 39568 366854 39888 366938
rect 39568 366618 39610 366854
rect 39846 366618 39888 366854
rect 39568 366586 39888 366618
rect 70288 367174 70608 367206
rect 70288 366938 70330 367174
rect 70566 366938 70608 367174
rect 70288 366854 70608 366938
rect 70288 366618 70330 366854
rect 70566 366618 70608 366854
rect 70288 366586 70608 366618
rect 101008 367174 101328 367206
rect 101008 366938 101050 367174
rect 101286 366938 101328 367174
rect 101008 366854 101328 366938
rect 101008 366618 101050 366854
rect 101286 366618 101328 366854
rect 101008 366586 101328 366618
rect 131728 367174 132048 367206
rect 131728 366938 131770 367174
rect 132006 366938 132048 367174
rect 131728 366854 132048 366938
rect 131728 366618 131770 366854
rect 132006 366618 132048 366854
rect 131728 366586 132048 366618
rect 162448 367174 162768 367206
rect 162448 366938 162490 367174
rect 162726 366938 162768 367174
rect 162448 366854 162768 366938
rect 162448 366618 162490 366854
rect 162726 366618 162768 366854
rect 162448 366586 162768 366618
rect 193168 367174 193488 367206
rect 193168 366938 193210 367174
rect 193446 366938 193488 367174
rect 193168 366854 193488 366938
rect 193168 366618 193210 366854
rect 193446 366618 193488 366854
rect 193168 366586 193488 366618
rect 223888 367174 224208 367206
rect 223888 366938 223930 367174
rect 224166 366938 224208 367174
rect 223888 366854 224208 366938
rect 223888 366618 223930 366854
rect 224166 366618 224208 366854
rect 223888 366586 224208 366618
rect 254608 367174 254928 367206
rect 254608 366938 254650 367174
rect 254886 366938 254928 367174
rect 254608 366854 254928 366938
rect 254608 366618 254650 366854
rect 254886 366618 254928 366854
rect 254608 366586 254928 366618
rect 285328 367174 285648 367206
rect 285328 366938 285370 367174
rect 285606 366938 285648 367174
rect 285328 366854 285648 366938
rect 285328 366618 285370 366854
rect 285606 366618 285648 366854
rect 285328 366586 285648 366618
rect 316048 367174 316368 367206
rect 316048 366938 316090 367174
rect 316326 366938 316368 367174
rect 316048 366854 316368 366938
rect 316048 366618 316090 366854
rect 316326 366618 316368 366854
rect 316048 366586 316368 366618
rect 346768 367174 347088 367206
rect 346768 366938 346810 367174
rect 347046 366938 347088 367174
rect 346768 366854 347088 366938
rect 346768 366618 346810 366854
rect 347046 366618 347088 366854
rect 346768 366586 347088 366618
rect 54928 363454 55248 363486
rect 54928 363218 54970 363454
rect 55206 363218 55248 363454
rect 54928 363134 55248 363218
rect 54928 362898 54970 363134
rect 55206 362898 55248 363134
rect 54928 362866 55248 362898
rect 85648 363454 85968 363486
rect 85648 363218 85690 363454
rect 85926 363218 85968 363454
rect 85648 363134 85968 363218
rect 85648 362898 85690 363134
rect 85926 362898 85968 363134
rect 85648 362866 85968 362898
rect 116368 363454 116688 363486
rect 116368 363218 116410 363454
rect 116646 363218 116688 363454
rect 116368 363134 116688 363218
rect 116368 362898 116410 363134
rect 116646 362898 116688 363134
rect 116368 362866 116688 362898
rect 147088 363454 147408 363486
rect 147088 363218 147130 363454
rect 147366 363218 147408 363454
rect 147088 363134 147408 363218
rect 147088 362898 147130 363134
rect 147366 362898 147408 363134
rect 147088 362866 147408 362898
rect 177808 363454 178128 363486
rect 177808 363218 177850 363454
rect 178086 363218 178128 363454
rect 177808 363134 178128 363218
rect 177808 362898 177850 363134
rect 178086 362898 178128 363134
rect 177808 362866 178128 362898
rect 208528 363454 208848 363486
rect 208528 363218 208570 363454
rect 208806 363218 208848 363454
rect 208528 363134 208848 363218
rect 208528 362898 208570 363134
rect 208806 362898 208848 363134
rect 208528 362866 208848 362898
rect 239248 363454 239568 363486
rect 239248 363218 239290 363454
rect 239526 363218 239568 363454
rect 239248 363134 239568 363218
rect 239248 362898 239290 363134
rect 239526 362898 239568 363134
rect 239248 362866 239568 362898
rect 269968 363454 270288 363486
rect 269968 363218 270010 363454
rect 270246 363218 270288 363454
rect 269968 363134 270288 363218
rect 269968 362898 270010 363134
rect 270246 362898 270288 363134
rect 269968 362866 270288 362898
rect 300688 363454 301008 363486
rect 300688 363218 300730 363454
rect 300966 363218 301008 363454
rect 300688 363134 301008 363218
rect 300688 362898 300730 363134
rect 300966 362898 301008 363134
rect 300688 362866 301008 362898
rect 331408 363454 331728 363486
rect 331408 363218 331450 363454
rect 331686 363218 331728 363454
rect 331408 363134 331728 363218
rect 331408 362898 331450 363134
rect 331686 362898 331728 363134
rect 331408 362866 331728 362898
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 27834 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 28454 353494
rect 27834 353174 28454 353258
rect 27834 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 28454 353174
rect 24208 327454 24528 327486
rect 24208 327218 24250 327454
rect 24486 327218 24528 327454
rect 24208 327134 24528 327218
rect 24208 326898 24250 327134
rect 24486 326898 24528 327134
rect 24208 326866 24528 326898
rect 20394 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 21014 310054
rect 20394 309734 21014 309818
rect 20394 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 21014 309734
rect 20394 274054 21014 309498
rect 27834 317494 28454 352938
rect 39568 331174 39888 331206
rect 39568 330938 39610 331174
rect 39846 330938 39888 331174
rect 39568 330854 39888 330938
rect 39568 330618 39610 330854
rect 39846 330618 39888 330854
rect 39568 330586 39888 330618
rect 70288 331174 70608 331206
rect 70288 330938 70330 331174
rect 70566 330938 70608 331174
rect 70288 330854 70608 330938
rect 70288 330618 70330 330854
rect 70566 330618 70608 330854
rect 70288 330586 70608 330618
rect 101008 331174 101328 331206
rect 101008 330938 101050 331174
rect 101286 330938 101328 331174
rect 101008 330854 101328 330938
rect 101008 330618 101050 330854
rect 101286 330618 101328 330854
rect 101008 330586 101328 330618
rect 131728 331174 132048 331206
rect 131728 330938 131770 331174
rect 132006 330938 132048 331174
rect 131728 330854 132048 330938
rect 131728 330618 131770 330854
rect 132006 330618 132048 330854
rect 131728 330586 132048 330618
rect 162448 331174 162768 331206
rect 162448 330938 162490 331174
rect 162726 330938 162768 331174
rect 162448 330854 162768 330938
rect 162448 330618 162490 330854
rect 162726 330618 162768 330854
rect 162448 330586 162768 330618
rect 193168 331174 193488 331206
rect 193168 330938 193210 331174
rect 193446 330938 193488 331174
rect 193168 330854 193488 330938
rect 193168 330618 193210 330854
rect 193446 330618 193488 330854
rect 193168 330586 193488 330618
rect 223888 331174 224208 331206
rect 223888 330938 223930 331174
rect 224166 330938 224208 331174
rect 223888 330854 224208 330938
rect 223888 330618 223930 330854
rect 224166 330618 224208 330854
rect 223888 330586 224208 330618
rect 254608 331174 254928 331206
rect 254608 330938 254650 331174
rect 254886 330938 254928 331174
rect 254608 330854 254928 330938
rect 254608 330618 254650 330854
rect 254886 330618 254928 330854
rect 254608 330586 254928 330618
rect 285328 331174 285648 331206
rect 285328 330938 285370 331174
rect 285606 330938 285648 331174
rect 285328 330854 285648 330938
rect 285328 330618 285370 330854
rect 285606 330618 285648 330854
rect 285328 330586 285648 330618
rect 316048 331174 316368 331206
rect 316048 330938 316090 331174
rect 316326 330938 316368 331174
rect 316048 330854 316368 330938
rect 316048 330618 316090 330854
rect 316326 330618 316368 330854
rect 316048 330586 316368 330618
rect 346768 331174 347088 331206
rect 346768 330938 346810 331174
rect 347046 330938 347088 331174
rect 346768 330854 347088 330938
rect 346768 330618 346810 330854
rect 347046 330618 347088 330854
rect 346768 330586 347088 330618
rect 54928 327454 55248 327486
rect 54928 327218 54970 327454
rect 55206 327218 55248 327454
rect 54928 327134 55248 327218
rect 54928 326898 54970 327134
rect 55206 326898 55248 327134
rect 54928 326866 55248 326898
rect 85648 327454 85968 327486
rect 85648 327218 85690 327454
rect 85926 327218 85968 327454
rect 85648 327134 85968 327218
rect 85648 326898 85690 327134
rect 85926 326898 85968 327134
rect 85648 326866 85968 326898
rect 116368 327454 116688 327486
rect 116368 327218 116410 327454
rect 116646 327218 116688 327454
rect 116368 327134 116688 327218
rect 116368 326898 116410 327134
rect 116646 326898 116688 327134
rect 116368 326866 116688 326898
rect 147088 327454 147408 327486
rect 147088 327218 147130 327454
rect 147366 327218 147408 327454
rect 147088 327134 147408 327218
rect 147088 326898 147130 327134
rect 147366 326898 147408 327134
rect 147088 326866 147408 326898
rect 177808 327454 178128 327486
rect 177808 327218 177850 327454
rect 178086 327218 178128 327454
rect 177808 327134 178128 327218
rect 177808 326898 177850 327134
rect 178086 326898 178128 327134
rect 177808 326866 178128 326898
rect 208528 327454 208848 327486
rect 208528 327218 208570 327454
rect 208806 327218 208848 327454
rect 208528 327134 208848 327218
rect 208528 326898 208570 327134
rect 208806 326898 208848 327134
rect 208528 326866 208848 326898
rect 239248 327454 239568 327486
rect 239248 327218 239290 327454
rect 239526 327218 239568 327454
rect 239248 327134 239568 327218
rect 239248 326898 239290 327134
rect 239526 326898 239568 327134
rect 239248 326866 239568 326898
rect 269968 327454 270288 327486
rect 269968 327218 270010 327454
rect 270246 327218 270288 327454
rect 269968 327134 270288 327218
rect 269968 326898 270010 327134
rect 270246 326898 270288 327134
rect 269968 326866 270288 326898
rect 300688 327454 301008 327486
rect 300688 327218 300730 327454
rect 300966 327218 301008 327454
rect 300688 327134 301008 327218
rect 300688 326898 300730 327134
rect 300966 326898 301008 327134
rect 300688 326866 301008 326898
rect 331408 327454 331728 327486
rect 331408 327218 331450 327454
rect 331686 327218 331728 327454
rect 331408 327134 331728 327218
rect 331408 326898 331450 327134
rect 331686 326898 331728 327134
rect 331408 326866 331728 326898
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 27834 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 28454 317494
rect 27834 317174 28454 317258
rect 27834 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 28454 317174
rect 24208 291454 24528 291486
rect 24208 291218 24250 291454
rect 24486 291218 24528 291454
rect 24208 291134 24528 291218
rect 24208 290898 24250 291134
rect 24486 290898 24528 291134
rect 24208 290866 24528 290898
rect 20394 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 21014 274054
rect 20394 273734 21014 273818
rect 20394 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 21014 273734
rect 20394 238054 21014 273498
rect 27834 281494 28454 316938
rect 39568 295174 39888 295206
rect 39568 294938 39610 295174
rect 39846 294938 39888 295174
rect 39568 294854 39888 294938
rect 39568 294618 39610 294854
rect 39846 294618 39888 294854
rect 39568 294586 39888 294618
rect 70288 295174 70608 295206
rect 70288 294938 70330 295174
rect 70566 294938 70608 295174
rect 70288 294854 70608 294938
rect 70288 294618 70330 294854
rect 70566 294618 70608 294854
rect 70288 294586 70608 294618
rect 101008 295174 101328 295206
rect 101008 294938 101050 295174
rect 101286 294938 101328 295174
rect 101008 294854 101328 294938
rect 101008 294618 101050 294854
rect 101286 294618 101328 294854
rect 101008 294586 101328 294618
rect 131728 295174 132048 295206
rect 131728 294938 131770 295174
rect 132006 294938 132048 295174
rect 131728 294854 132048 294938
rect 131728 294618 131770 294854
rect 132006 294618 132048 294854
rect 131728 294586 132048 294618
rect 162448 295174 162768 295206
rect 162448 294938 162490 295174
rect 162726 294938 162768 295174
rect 162448 294854 162768 294938
rect 162448 294618 162490 294854
rect 162726 294618 162768 294854
rect 162448 294586 162768 294618
rect 193168 295174 193488 295206
rect 193168 294938 193210 295174
rect 193446 294938 193488 295174
rect 193168 294854 193488 294938
rect 193168 294618 193210 294854
rect 193446 294618 193488 294854
rect 193168 294586 193488 294618
rect 223888 295174 224208 295206
rect 223888 294938 223930 295174
rect 224166 294938 224208 295174
rect 223888 294854 224208 294938
rect 223888 294618 223930 294854
rect 224166 294618 224208 294854
rect 223888 294586 224208 294618
rect 254608 295174 254928 295206
rect 254608 294938 254650 295174
rect 254886 294938 254928 295174
rect 254608 294854 254928 294938
rect 254608 294618 254650 294854
rect 254886 294618 254928 294854
rect 254608 294586 254928 294618
rect 285328 295174 285648 295206
rect 285328 294938 285370 295174
rect 285606 294938 285648 295174
rect 285328 294854 285648 294938
rect 285328 294618 285370 294854
rect 285606 294618 285648 294854
rect 285328 294586 285648 294618
rect 316048 295174 316368 295206
rect 316048 294938 316090 295174
rect 316326 294938 316368 295174
rect 316048 294854 316368 294938
rect 316048 294618 316090 294854
rect 316326 294618 316368 294854
rect 316048 294586 316368 294618
rect 346768 295174 347088 295206
rect 346768 294938 346810 295174
rect 347046 294938 347088 295174
rect 346768 294854 347088 294938
rect 346768 294618 346810 294854
rect 347046 294618 347088 294854
rect 346768 294586 347088 294618
rect 54928 291454 55248 291486
rect 54928 291218 54970 291454
rect 55206 291218 55248 291454
rect 54928 291134 55248 291218
rect 54928 290898 54970 291134
rect 55206 290898 55248 291134
rect 54928 290866 55248 290898
rect 85648 291454 85968 291486
rect 85648 291218 85690 291454
rect 85926 291218 85968 291454
rect 85648 291134 85968 291218
rect 85648 290898 85690 291134
rect 85926 290898 85968 291134
rect 85648 290866 85968 290898
rect 116368 291454 116688 291486
rect 116368 291218 116410 291454
rect 116646 291218 116688 291454
rect 116368 291134 116688 291218
rect 116368 290898 116410 291134
rect 116646 290898 116688 291134
rect 116368 290866 116688 290898
rect 147088 291454 147408 291486
rect 147088 291218 147130 291454
rect 147366 291218 147408 291454
rect 147088 291134 147408 291218
rect 147088 290898 147130 291134
rect 147366 290898 147408 291134
rect 147088 290866 147408 290898
rect 177808 291454 178128 291486
rect 177808 291218 177850 291454
rect 178086 291218 178128 291454
rect 177808 291134 178128 291218
rect 177808 290898 177850 291134
rect 178086 290898 178128 291134
rect 177808 290866 178128 290898
rect 208528 291454 208848 291486
rect 208528 291218 208570 291454
rect 208806 291218 208848 291454
rect 208528 291134 208848 291218
rect 208528 290898 208570 291134
rect 208806 290898 208848 291134
rect 208528 290866 208848 290898
rect 239248 291454 239568 291486
rect 239248 291218 239290 291454
rect 239526 291218 239568 291454
rect 239248 291134 239568 291218
rect 239248 290898 239290 291134
rect 239526 290898 239568 291134
rect 239248 290866 239568 290898
rect 269968 291454 270288 291486
rect 269968 291218 270010 291454
rect 270246 291218 270288 291454
rect 269968 291134 270288 291218
rect 269968 290898 270010 291134
rect 270246 290898 270288 291134
rect 269968 290866 270288 290898
rect 300688 291454 301008 291486
rect 300688 291218 300730 291454
rect 300966 291218 301008 291454
rect 300688 291134 301008 291218
rect 300688 290898 300730 291134
rect 300966 290898 301008 291134
rect 300688 290866 301008 290898
rect 331408 291454 331728 291486
rect 331408 291218 331450 291454
rect 331686 291218 331728 291454
rect 331408 291134 331728 291218
rect 331408 290898 331450 291134
rect 331686 290898 331728 291134
rect 331408 290866 331728 290898
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 27834 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 28454 281494
rect 27834 281174 28454 281258
rect 27834 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 28454 281174
rect 24208 255454 24528 255486
rect 24208 255218 24250 255454
rect 24486 255218 24528 255454
rect 24208 255134 24528 255218
rect 24208 254898 24250 255134
rect 24486 254898 24528 255134
rect 24208 254866 24528 254898
rect 20394 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 21014 238054
rect 20394 237734 21014 237818
rect 20394 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 21014 237734
rect 20394 202054 21014 237498
rect 27834 245494 28454 280938
rect 39568 259174 39888 259206
rect 39568 258938 39610 259174
rect 39846 258938 39888 259174
rect 39568 258854 39888 258938
rect 39568 258618 39610 258854
rect 39846 258618 39888 258854
rect 39568 258586 39888 258618
rect 70288 259174 70608 259206
rect 70288 258938 70330 259174
rect 70566 258938 70608 259174
rect 70288 258854 70608 258938
rect 70288 258618 70330 258854
rect 70566 258618 70608 258854
rect 70288 258586 70608 258618
rect 101008 259174 101328 259206
rect 101008 258938 101050 259174
rect 101286 258938 101328 259174
rect 101008 258854 101328 258938
rect 101008 258618 101050 258854
rect 101286 258618 101328 258854
rect 101008 258586 101328 258618
rect 131728 259174 132048 259206
rect 131728 258938 131770 259174
rect 132006 258938 132048 259174
rect 131728 258854 132048 258938
rect 131728 258618 131770 258854
rect 132006 258618 132048 258854
rect 131728 258586 132048 258618
rect 162448 259174 162768 259206
rect 162448 258938 162490 259174
rect 162726 258938 162768 259174
rect 162448 258854 162768 258938
rect 162448 258618 162490 258854
rect 162726 258618 162768 258854
rect 162448 258586 162768 258618
rect 193168 259174 193488 259206
rect 193168 258938 193210 259174
rect 193446 258938 193488 259174
rect 193168 258854 193488 258938
rect 193168 258618 193210 258854
rect 193446 258618 193488 258854
rect 193168 258586 193488 258618
rect 223888 259174 224208 259206
rect 223888 258938 223930 259174
rect 224166 258938 224208 259174
rect 223888 258854 224208 258938
rect 223888 258618 223930 258854
rect 224166 258618 224208 258854
rect 223888 258586 224208 258618
rect 254608 259174 254928 259206
rect 254608 258938 254650 259174
rect 254886 258938 254928 259174
rect 254608 258854 254928 258938
rect 254608 258618 254650 258854
rect 254886 258618 254928 258854
rect 254608 258586 254928 258618
rect 285328 259174 285648 259206
rect 285328 258938 285370 259174
rect 285606 258938 285648 259174
rect 285328 258854 285648 258938
rect 285328 258618 285370 258854
rect 285606 258618 285648 258854
rect 285328 258586 285648 258618
rect 316048 259174 316368 259206
rect 316048 258938 316090 259174
rect 316326 258938 316368 259174
rect 316048 258854 316368 258938
rect 316048 258618 316090 258854
rect 316326 258618 316368 258854
rect 316048 258586 316368 258618
rect 346768 259174 347088 259206
rect 346768 258938 346810 259174
rect 347046 258938 347088 259174
rect 346768 258854 347088 258938
rect 346768 258618 346810 258854
rect 347046 258618 347088 258854
rect 346768 258586 347088 258618
rect 54928 255454 55248 255486
rect 54928 255218 54970 255454
rect 55206 255218 55248 255454
rect 54928 255134 55248 255218
rect 54928 254898 54970 255134
rect 55206 254898 55248 255134
rect 54928 254866 55248 254898
rect 85648 255454 85968 255486
rect 85648 255218 85690 255454
rect 85926 255218 85968 255454
rect 85648 255134 85968 255218
rect 85648 254898 85690 255134
rect 85926 254898 85968 255134
rect 85648 254866 85968 254898
rect 116368 255454 116688 255486
rect 116368 255218 116410 255454
rect 116646 255218 116688 255454
rect 116368 255134 116688 255218
rect 116368 254898 116410 255134
rect 116646 254898 116688 255134
rect 116368 254866 116688 254898
rect 147088 255454 147408 255486
rect 147088 255218 147130 255454
rect 147366 255218 147408 255454
rect 147088 255134 147408 255218
rect 147088 254898 147130 255134
rect 147366 254898 147408 255134
rect 147088 254866 147408 254898
rect 177808 255454 178128 255486
rect 177808 255218 177850 255454
rect 178086 255218 178128 255454
rect 177808 255134 178128 255218
rect 177808 254898 177850 255134
rect 178086 254898 178128 255134
rect 177808 254866 178128 254898
rect 208528 255454 208848 255486
rect 208528 255218 208570 255454
rect 208806 255218 208848 255454
rect 208528 255134 208848 255218
rect 208528 254898 208570 255134
rect 208806 254898 208848 255134
rect 208528 254866 208848 254898
rect 239248 255454 239568 255486
rect 239248 255218 239290 255454
rect 239526 255218 239568 255454
rect 239248 255134 239568 255218
rect 239248 254898 239290 255134
rect 239526 254898 239568 255134
rect 239248 254866 239568 254898
rect 269968 255454 270288 255486
rect 269968 255218 270010 255454
rect 270246 255218 270288 255454
rect 269968 255134 270288 255218
rect 269968 254898 270010 255134
rect 270246 254898 270288 255134
rect 269968 254866 270288 254898
rect 300688 255454 301008 255486
rect 300688 255218 300730 255454
rect 300966 255218 301008 255454
rect 300688 255134 301008 255218
rect 300688 254898 300730 255134
rect 300966 254898 301008 255134
rect 300688 254866 301008 254898
rect 331408 255454 331728 255486
rect 331408 255218 331450 255454
rect 331686 255218 331728 255454
rect 331408 255134 331728 255218
rect 331408 254898 331450 255134
rect 331686 254898 331728 255134
rect 331408 254866 331728 254898
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 27834 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 28454 245494
rect 27834 245174 28454 245258
rect 27834 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 28454 245174
rect 24208 219454 24528 219486
rect 24208 219218 24250 219454
rect 24486 219218 24528 219454
rect 24208 219134 24528 219218
rect 24208 218898 24250 219134
rect 24486 218898 24528 219134
rect 24208 218866 24528 218898
rect 20394 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 21014 202054
rect 20394 201734 21014 201818
rect 20394 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 21014 201734
rect 20394 166054 21014 201498
rect 27834 209494 28454 244938
rect 39568 223174 39888 223206
rect 39568 222938 39610 223174
rect 39846 222938 39888 223174
rect 39568 222854 39888 222938
rect 39568 222618 39610 222854
rect 39846 222618 39888 222854
rect 39568 222586 39888 222618
rect 70288 223174 70608 223206
rect 70288 222938 70330 223174
rect 70566 222938 70608 223174
rect 70288 222854 70608 222938
rect 70288 222618 70330 222854
rect 70566 222618 70608 222854
rect 70288 222586 70608 222618
rect 101008 223174 101328 223206
rect 101008 222938 101050 223174
rect 101286 222938 101328 223174
rect 101008 222854 101328 222938
rect 101008 222618 101050 222854
rect 101286 222618 101328 222854
rect 101008 222586 101328 222618
rect 131728 223174 132048 223206
rect 131728 222938 131770 223174
rect 132006 222938 132048 223174
rect 131728 222854 132048 222938
rect 131728 222618 131770 222854
rect 132006 222618 132048 222854
rect 131728 222586 132048 222618
rect 162448 223174 162768 223206
rect 162448 222938 162490 223174
rect 162726 222938 162768 223174
rect 162448 222854 162768 222938
rect 162448 222618 162490 222854
rect 162726 222618 162768 222854
rect 162448 222586 162768 222618
rect 193168 223174 193488 223206
rect 193168 222938 193210 223174
rect 193446 222938 193488 223174
rect 193168 222854 193488 222938
rect 193168 222618 193210 222854
rect 193446 222618 193488 222854
rect 193168 222586 193488 222618
rect 223888 223174 224208 223206
rect 223888 222938 223930 223174
rect 224166 222938 224208 223174
rect 223888 222854 224208 222938
rect 223888 222618 223930 222854
rect 224166 222618 224208 222854
rect 223888 222586 224208 222618
rect 254608 223174 254928 223206
rect 254608 222938 254650 223174
rect 254886 222938 254928 223174
rect 254608 222854 254928 222938
rect 254608 222618 254650 222854
rect 254886 222618 254928 222854
rect 254608 222586 254928 222618
rect 285328 223174 285648 223206
rect 285328 222938 285370 223174
rect 285606 222938 285648 223174
rect 285328 222854 285648 222938
rect 285328 222618 285370 222854
rect 285606 222618 285648 222854
rect 285328 222586 285648 222618
rect 316048 223174 316368 223206
rect 316048 222938 316090 223174
rect 316326 222938 316368 223174
rect 316048 222854 316368 222938
rect 316048 222618 316090 222854
rect 316326 222618 316368 222854
rect 316048 222586 316368 222618
rect 346768 223174 347088 223206
rect 346768 222938 346810 223174
rect 347046 222938 347088 223174
rect 346768 222854 347088 222938
rect 346768 222618 346810 222854
rect 347046 222618 347088 222854
rect 346768 222586 347088 222618
rect 54928 219454 55248 219486
rect 54928 219218 54970 219454
rect 55206 219218 55248 219454
rect 54928 219134 55248 219218
rect 54928 218898 54970 219134
rect 55206 218898 55248 219134
rect 54928 218866 55248 218898
rect 85648 219454 85968 219486
rect 85648 219218 85690 219454
rect 85926 219218 85968 219454
rect 85648 219134 85968 219218
rect 85648 218898 85690 219134
rect 85926 218898 85968 219134
rect 85648 218866 85968 218898
rect 116368 219454 116688 219486
rect 116368 219218 116410 219454
rect 116646 219218 116688 219454
rect 116368 219134 116688 219218
rect 116368 218898 116410 219134
rect 116646 218898 116688 219134
rect 116368 218866 116688 218898
rect 147088 219454 147408 219486
rect 147088 219218 147130 219454
rect 147366 219218 147408 219454
rect 147088 219134 147408 219218
rect 147088 218898 147130 219134
rect 147366 218898 147408 219134
rect 147088 218866 147408 218898
rect 177808 219454 178128 219486
rect 177808 219218 177850 219454
rect 178086 219218 178128 219454
rect 177808 219134 178128 219218
rect 177808 218898 177850 219134
rect 178086 218898 178128 219134
rect 177808 218866 178128 218898
rect 208528 219454 208848 219486
rect 208528 219218 208570 219454
rect 208806 219218 208848 219454
rect 208528 219134 208848 219218
rect 208528 218898 208570 219134
rect 208806 218898 208848 219134
rect 208528 218866 208848 218898
rect 239248 219454 239568 219486
rect 239248 219218 239290 219454
rect 239526 219218 239568 219454
rect 239248 219134 239568 219218
rect 239248 218898 239290 219134
rect 239526 218898 239568 219134
rect 239248 218866 239568 218898
rect 269968 219454 270288 219486
rect 269968 219218 270010 219454
rect 270246 219218 270288 219454
rect 269968 219134 270288 219218
rect 269968 218898 270010 219134
rect 270246 218898 270288 219134
rect 269968 218866 270288 218898
rect 300688 219454 301008 219486
rect 300688 219218 300730 219454
rect 300966 219218 301008 219454
rect 300688 219134 301008 219218
rect 300688 218898 300730 219134
rect 300966 218898 301008 219134
rect 300688 218866 301008 218898
rect 331408 219454 331728 219486
rect 331408 219218 331450 219454
rect 331686 219218 331728 219454
rect 331408 219134 331728 219218
rect 331408 218898 331450 219134
rect 331686 218898 331728 219134
rect 331408 218866 331728 218898
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 27834 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 28454 209494
rect 27834 209174 28454 209258
rect 27834 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 28454 209174
rect 24208 183454 24528 183486
rect 24208 183218 24250 183454
rect 24486 183218 24528 183454
rect 24208 183134 24528 183218
rect 24208 182898 24250 183134
rect 24486 182898 24528 183134
rect 24208 182866 24528 182898
rect 20394 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 21014 166054
rect 20394 165734 21014 165818
rect 20394 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 21014 165734
rect 20394 130054 21014 165498
rect 27834 173494 28454 208938
rect 39568 187174 39888 187206
rect 39568 186938 39610 187174
rect 39846 186938 39888 187174
rect 39568 186854 39888 186938
rect 39568 186618 39610 186854
rect 39846 186618 39888 186854
rect 39568 186586 39888 186618
rect 70288 187174 70608 187206
rect 70288 186938 70330 187174
rect 70566 186938 70608 187174
rect 70288 186854 70608 186938
rect 70288 186618 70330 186854
rect 70566 186618 70608 186854
rect 70288 186586 70608 186618
rect 101008 187174 101328 187206
rect 101008 186938 101050 187174
rect 101286 186938 101328 187174
rect 101008 186854 101328 186938
rect 101008 186618 101050 186854
rect 101286 186618 101328 186854
rect 101008 186586 101328 186618
rect 131728 187174 132048 187206
rect 131728 186938 131770 187174
rect 132006 186938 132048 187174
rect 131728 186854 132048 186938
rect 131728 186618 131770 186854
rect 132006 186618 132048 186854
rect 131728 186586 132048 186618
rect 162448 187174 162768 187206
rect 162448 186938 162490 187174
rect 162726 186938 162768 187174
rect 162448 186854 162768 186938
rect 162448 186618 162490 186854
rect 162726 186618 162768 186854
rect 162448 186586 162768 186618
rect 193168 187174 193488 187206
rect 193168 186938 193210 187174
rect 193446 186938 193488 187174
rect 193168 186854 193488 186938
rect 193168 186618 193210 186854
rect 193446 186618 193488 186854
rect 193168 186586 193488 186618
rect 223888 187174 224208 187206
rect 223888 186938 223930 187174
rect 224166 186938 224208 187174
rect 223888 186854 224208 186938
rect 223888 186618 223930 186854
rect 224166 186618 224208 186854
rect 223888 186586 224208 186618
rect 254608 187174 254928 187206
rect 254608 186938 254650 187174
rect 254886 186938 254928 187174
rect 254608 186854 254928 186938
rect 254608 186618 254650 186854
rect 254886 186618 254928 186854
rect 254608 186586 254928 186618
rect 285328 187174 285648 187206
rect 285328 186938 285370 187174
rect 285606 186938 285648 187174
rect 285328 186854 285648 186938
rect 285328 186618 285370 186854
rect 285606 186618 285648 186854
rect 285328 186586 285648 186618
rect 316048 187174 316368 187206
rect 316048 186938 316090 187174
rect 316326 186938 316368 187174
rect 316048 186854 316368 186938
rect 316048 186618 316090 186854
rect 316326 186618 316368 186854
rect 316048 186586 316368 186618
rect 346768 187174 347088 187206
rect 346768 186938 346810 187174
rect 347046 186938 347088 187174
rect 346768 186854 347088 186938
rect 346768 186618 346810 186854
rect 347046 186618 347088 186854
rect 346768 186586 347088 186618
rect 54928 183454 55248 183486
rect 54928 183218 54970 183454
rect 55206 183218 55248 183454
rect 54928 183134 55248 183218
rect 54928 182898 54970 183134
rect 55206 182898 55248 183134
rect 54928 182866 55248 182898
rect 85648 183454 85968 183486
rect 85648 183218 85690 183454
rect 85926 183218 85968 183454
rect 85648 183134 85968 183218
rect 85648 182898 85690 183134
rect 85926 182898 85968 183134
rect 85648 182866 85968 182898
rect 116368 183454 116688 183486
rect 116368 183218 116410 183454
rect 116646 183218 116688 183454
rect 116368 183134 116688 183218
rect 116368 182898 116410 183134
rect 116646 182898 116688 183134
rect 116368 182866 116688 182898
rect 147088 183454 147408 183486
rect 147088 183218 147130 183454
rect 147366 183218 147408 183454
rect 147088 183134 147408 183218
rect 147088 182898 147130 183134
rect 147366 182898 147408 183134
rect 147088 182866 147408 182898
rect 177808 183454 178128 183486
rect 177808 183218 177850 183454
rect 178086 183218 178128 183454
rect 177808 183134 178128 183218
rect 177808 182898 177850 183134
rect 178086 182898 178128 183134
rect 177808 182866 178128 182898
rect 208528 183454 208848 183486
rect 208528 183218 208570 183454
rect 208806 183218 208848 183454
rect 208528 183134 208848 183218
rect 208528 182898 208570 183134
rect 208806 182898 208848 183134
rect 208528 182866 208848 182898
rect 239248 183454 239568 183486
rect 239248 183218 239290 183454
rect 239526 183218 239568 183454
rect 239248 183134 239568 183218
rect 239248 182898 239290 183134
rect 239526 182898 239568 183134
rect 239248 182866 239568 182898
rect 269968 183454 270288 183486
rect 269968 183218 270010 183454
rect 270246 183218 270288 183454
rect 269968 183134 270288 183218
rect 269968 182898 270010 183134
rect 270246 182898 270288 183134
rect 269968 182866 270288 182898
rect 300688 183454 301008 183486
rect 300688 183218 300730 183454
rect 300966 183218 301008 183454
rect 300688 183134 301008 183218
rect 300688 182898 300730 183134
rect 300966 182898 301008 183134
rect 300688 182866 301008 182898
rect 331408 183454 331728 183486
rect 331408 183218 331450 183454
rect 331686 183218 331728 183454
rect 331408 183134 331728 183218
rect 331408 182898 331450 183134
rect 331686 182898 331728 183134
rect 331408 182866 331728 182898
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 27834 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 28454 173494
rect 27834 173174 28454 173258
rect 27834 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 28454 173174
rect 24208 147454 24528 147486
rect 24208 147218 24250 147454
rect 24486 147218 24528 147454
rect 24208 147134 24528 147218
rect 24208 146898 24250 147134
rect 24486 146898 24528 147134
rect 24208 146866 24528 146898
rect 20394 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 21014 130054
rect 20394 129734 21014 129818
rect 20394 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 21014 129734
rect 20394 94054 21014 129498
rect 27834 137494 28454 172938
rect 39568 151174 39888 151206
rect 39568 150938 39610 151174
rect 39846 150938 39888 151174
rect 39568 150854 39888 150938
rect 39568 150618 39610 150854
rect 39846 150618 39888 150854
rect 39568 150586 39888 150618
rect 70288 151174 70608 151206
rect 70288 150938 70330 151174
rect 70566 150938 70608 151174
rect 70288 150854 70608 150938
rect 70288 150618 70330 150854
rect 70566 150618 70608 150854
rect 70288 150586 70608 150618
rect 101008 151174 101328 151206
rect 101008 150938 101050 151174
rect 101286 150938 101328 151174
rect 101008 150854 101328 150938
rect 101008 150618 101050 150854
rect 101286 150618 101328 150854
rect 101008 150586 101328 150618
rect 131728 151174 132048 151206
rect 131728 150938 131770 151174
rect 132006 150938 132048 151174
rect 131728 150854 132048 150938
rect 131728 150618 131770 150854
rect 132006 150618 132048 150854
rect 131728 150586 132048 150618
rect 162448 151174 162768 151206
rect 162448 150938 162490 151174
rect 162726 150938 162768 151174
rect 162448 150854 162768 150938
rect 162448 150618 162490 150854
rect 162726 150618 162768 150854
rect 162448 150586 162768 150618
rect 193168 151174 193488 151206
rect 193168 150938 193210 151174
rect 193446 150938 193488 151174
rect 193168 150854 193488 150938
rect 193168 150618 193210 150854
rect 193446 150618 193488 150854
rect 193168 150586 193488 150618
rect 223888 151174 224208 151206
rect 223888 150938 223930 151174
rect 224166 150938 224208 151174
rect 223888 150854 224208 150938
rect 223888 150618 223930 150854
rect 224166 150618 224208 150854
rect 223888 150586 224208 150618
rect 254608 151174 254928 151206
rect 254608 150938 254650 151174
rect 254886 150938 254928 151174
rect 254608 150854 254928 150938
rect 254608 150618 254650 150854
rect 254886 150618 254928 150854
rect 254608 150586 254928 150618
rect 285328 151174 285648 151206
rect 285328 150938 285370 151174
rect 285606 150938 285648 151174
rect 285328 150854 285648 150938
rect 285328 150618 285370 150854
rect 285606 150618 285648 150854
rect 285328 150586 285648 150618
rect 316048 151174 316368 151206
rect 316048 150938 316090 151174
rect 316326 150938 316368 151174
rect 316048 150854 316368 150938
rect 316048 150618 316090 150854
rect 316326 150618 316368 150854
rect 316048 150586 316368 150618
rect 346768 151174 347088 151206
rect 346768 150938 346810 151174
rect 347046 150938 347088 151174
rect 346768 150854 347088 150938
rect 346768 150618 346810 150854
rect 347046 150618 347088 150854
rect 346768 150586 347088 150618
rect 54928 147454 55248 147486
rect 54928 147218 54970 147454
rect 55206 147218 55248 147454
rect 54928 147134 55248 147218
rect 54928 146898 54970 147134
rect 55206 146898 55248 147134
rect 54928 146866 55248 146898
rect 85648 147454 85968 147486
rect 85648 147218 85690 147454
rect 85926 147218 85968 147454
rect 85648 147134 85968 147218
rect 85648 146898 85690 147134
rect 85926 146898 85968 147134
rect 85648 146866 85968 146898
rect 116368 147454 116688 147486
rect 116368 147218 116410 147454
rect 116646 147218 116688 147454
rect 116368 147134 116688 147218
rect 116368 146898 116410 147134
rect 116646 146898 116688 147134
rect 116368 146866 116688 146898
rect 147088 147454 147408 147486
rect 147088 147218 147130 147454
rect 147366 147218 147408 147454
rect 147088 147134 147408 147218
rect 147088 146898 147130 147134
rect 147366 146898 147408 147134
rect 147088 146866 147408 146898
rect 177808 147454 178128 147486
rect 177808 147218 177850 147454
rect 178086 147218 178128 147454
rect 177808 147134 178128 147218
rect 177808 146898 177850 147134
rect 178086 146898 178128 147134
rect 177808 146866 178128 146898
rect 208528 147454 208848 147486
rect 208528 147218 208570 147454
rect 208806 147218 208848 147454
rect 208528 147134 208848 147218
rect 208528 146898 208570 147134
rect 208806 146898 208848 147134
rect 208528 146866 208848 146898
rect 239248 147454 239568 147486
rect 239248 147218 239290 147454
rect 239526 147218 239568 147454
rect 239248 147134 239568 147218
rect 239248 146898 239290 147134
rect 239526 146898 239568 147134
rect 239248 146866 239568 146898
rect 269968 147454 270288 147486
rect 269968 147218 270010 147454
rect 270246 147218 270288 147454
rect 269968 147134 270288 147218
rect 269968 146898 270010 147134
rect 270246 146898 270288 147134
rect 269968 146866 270288 146898
rect 300688 147454 301008 147486
rect 300688 147218 300730 147454
rect 300966 147218 301008 147454
rect 300688 147134 301008 147218
rect 300688 146898 300730 147134
rect 300966 146898 301008 147134
rect 300688 146866 301008 146898
rect 331408 147454 331728 147486
rect 331408 147218 331450 147454
rect 331686 147218 331728 147454
rect 331408 147134 331728 147218
rect 331408 146898 331450 147134
rect 331686 146898 331728 147134
rect 331408 146866 331728 146898
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 27834 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 28454 137494
rect 27834 137174 28454 137258
rect 27834 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 28454 137174
rect 24208 111454 24528 111486
rect 24208 111218 24250 111454
rect 24486 111218 24528 111454
rect 24208 111134 24528 111218
rect 24208 110898 24250 111134
rect 24486 110898 24528 111134
rect 24208 110866 24528 110898
rect 20394 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 21014 94054
rect 20394 93734 21014 93818
rect 20394 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 21014 93734
rect 20394 58054 21014 93498
rect 27834 101494 28454 136938
rect 39568 115174 39888 115206
rect 39568 114938 39610 115174
rect 39846 114938 39888 115174
rect 39568 114854 39888 114938
rect 39568 114618 39610 114854
rect 39846 114618 39888 114854
rect 39568 114586 39888 114618
rect 70288 115174 70608 115206
rect 70288 114938 70330 115174
rect 70566 114938 70608 115174
rect 70288 114854 70608 114938
rect 70288 114618 70330 114854
rect 70566 114618 70608 114854
rect 70288 114586 70608 114618
rect 101008 115174 101328 115206
rect 101008 114938 101050 115174
rect 101286 114938 101328 115174
rect 101008 114854 101328 114938
rect 101008 114618 101050 114854
rect 101286 114618 101328 114854
rect 101008 114586 101328 114618
rect 131728 115174 132048 115206
rect 131728 114938 131770 115174
rect 132006 114938 132048 115174
rect 131728 114854 132048 114938
rect 131728 114618 131770 114854
rect 132006 114618 132048 114854
rect 131728 114586 132048 114618
rect 162448 115174 162768 115206
rect 162448 114938 162490 115174
rect 162726 114938 162768 115174
rect 162448 114854 162768 114938
rect 162448 114618 162490 114854
rect 162726 114618 162768 114854
rect 162448 114586 162768 114618
rect 193168 115174 193488 115206
rect 193168 114938 193210 115174
rect 193446 114938 193488 115174
rect 193168 114854 193488 114938
rect 193168 114618 193210 114854
rect 193446 114618 193488 114854
rect 193168 114586 193488 114618
rect 223888 115174 224208 115206
rect 223888 114938 223930 115174
rect 224166 114938 224208 115174
rect 223888 114854 224208 114938
rect 223888 114618 223930 114854
rect 224166 114618 224208 114854
rect 223888 114586 224208 114618
rect 254608 115174 254928 115206
rect 254608 114938 254650 115174
rect 254886 114938 254928 115174
rect 254608 114854 254928 114938
rect 254608 114618 254650 114854
rect 254886 114618 254928 114854
rect 254608 114586 254928 114618
rect 285328 115174 285648 115206
rect 285328 114938 285370 115174
rect 285606 114938 285648 115174
rect 285328 114854 285648 114938
rect 285328 114618 285370 114854
rect 285606 114618 285648 114854
rect 285328 114586 285648 114618
rect 316048 115174 316368 115206
rect 316048 114938 316090 115174
rect 316326 114938 316368 115174
rect 316048 114854 316368 114938
rect 316048 114618 316090 114854
rect 316326 114618 316368 114854
rect 316048 114586 316368 114618
rect 346768 115174 347088 115206
rect 346768 114938 346810 115174
rect 347046 114938 347088 115174
rect 346768 114854 347088 114938
rect 346768 114618 346810 114854
rect 347046 114618 347088 114854
rect 346768 114586 347088 114618
rect 54928 111454 55248 111486
rect 54928 111218 54970 111454
rect 55206 111218 55248 111454
rect 54928 111134 55248 111218
rect 54928 110898 54970 111134
rect 55206 110898 55248 111134
rect 54928 110866 55248 110898
rect 85648 111454 85968 111486
rect 85648 111218 85690 111454
rect 85926 111218 85968 111454
rect 85648 111134 85968 111218
rect 85648 110898 85690 111134
rect 85926 110898 85968 111134
rect 85648 110866 85968 110898
rect 116368 111454 116688 111486
rect 116368 111218 116410 111454
rect 116646 111218 116688 111454
rect 116368 111134 116688 111218
rect 116368 110898 116410 111134
rect 116646 110898 116688 111134
rect 116368 110866 116688 110898
rect 147088 111454 147408 111486
rect 147088 111218 147130 111454
rect 147366 111218 147408 111454
rect 147088 111134 147408 111218
rect 147088 110898 147130 111134
rect 147366 110898 147408 111134
rect 147088 110866 147408 110898
rect 177808 111454 178128 111486
rect 177808 111218 177850 111454
rect 178086 111218 178128 111454
rect 177808 111134 178128 111218
rect 177808 110898 177850 111134
rect 178086 110898 178128 111134
rect 177808 110866 178128 110898
rect 208528 111454 208848 111486
rect 208528 111218 208570 111454
rect 208806 111218 208848 111454
rect 208528 111134 208848 111218
rect 208528 110898 208570 111134
rect 208806 110898 208848 111134
rect 208528 110866 208848 110898
rect 239248 111454 239568 111486
rect 239248 111218 239290 111454
rect 239526 111218 239568 111454
rect 239248 111134 239568 111218
rect 239248 110898 239290 111134
rect 239526 110898 239568 111134
rect 239248 110866 239568 110898
rect 269968 111454 270288 111486
rect 269968 111218 270010 111454
rect 270246 111218 270288 111454
rect 269968 111134 270288 111218
rect 269968 110898 270010 111134
rect 270246 110898 270288 111134
rect 269968 110866 270288 110898
rect 300688 111454 301008 111486
rect 300688 111218 300730 111454
rect 300966 111218 301008 111454
rect 300688 111134 301008 111218
rect 300688 110898 300730 111134
rect 300966 110898 301008 111134
rect 300688 110866 301008 110898
rect 331408 111454 331728 111486
rect 331408 111218 331450 111454
rect 331686 111218 331728 111454
rect 331408 111134 331728 111218
rect 331408 110898 331450 111134
rect 331686 110898 331728 111134
rect 331408 110866 331728 110898
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 27834 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 28454 101494
rect 27834 101174 28454 101258
rect 27834 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 28454 101174
rect 24208 75454 24528 75486
rect 24208 75218 24250 75454
rect 24486 75218 24528 75454
rect 24208 75134 24528 75218
rect 24208 74898 24250 75134
rect 24486 74898 24528 75134
rect 24208 74866 24528 74898
rect 20394 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 21014 58054
rect 20394 57734 21014 57818
rect 20394 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 21014 57734
rect 20394 22054 21014 57498
rect 27834 65494 28454 100938
rect 39568 79174 39888 79206
rect 39568 78938 39610 79174
rect 39846 78938 39888 79174
rect 39568 78854 39888 78938
rect 39568 78618 39610 78854
rect 39846 78618 39888 78854
rect 39568 78586 39888 78618
rect 70288 79174 70608 79206
rect 70288 78938 70330 79174
rect 70566 78938 70608 79174
rect 70288 78854 70608 78938
rect 70288 78618 70330 78854
rect 70566 78618 70608 78854
rect 70288 78586 70608 78618
rect 101008 79174 101328 79206
rect 101008 78938 101050 79174
rect 101286 78938 101328 79174
rect 101008 78854 101328 78938
rect 101008 78618 101050 78854
rect 101286 78618 101328 78854
rect 101008 78586 101328 78618
rect 131728 79174 132048 79206
rect 131728 78938 131770 79174
rect 132006 78938 132048 79174
rect 131728 78854 132048 78938
rect 131728 78618 131770 78854
rect 132006 78618 132048 78854
rect 131728 78586 132048 78618
rect 162448 79174 162768 79206
rect 162448 78938 162490 79174
rect 162726 78938 162768 79174
rect 162448 78854 162768 78938
rect 162448 78618 162490 78854
rect 162726 78618 162768 78854
rect 162448 78586 162768 78618
rect 193168 79174 193488 79206
rect 193168 78938 193210 79174
rect 193446 78938 193488 79174
rect 193168 78854 193488 78938
rect 193168 78618 193210 78854
rect 193446 78618 193488 78854
rect 193168 78586 193488 78618
rect 223888 79174 224208 79206
rect 223888 78938 223930 79174
rect 224166 78938 224208 79174
rect 223888 78854 224208 78938
rect 223888 78618 223930 78854
rect 224166 78618 224208 78854
rect 223888 78586 224208 78618
rect 254608 79174 254928 79206
rect 254608 78938 254650 79174
rect 254886 78938 254928 79174
rect 254608 78854 254928 78938
rect 254608 78618 254650 78854
rect 254886 78618 254928 78854
rect 254608 78586 254928 78618
rect 285328 79174 285648 79206
rect 285328 78938 285370 79174
rect 285606 78938 285648 79174
rect 285328 78854 285648 78938
rect 285328 78618 285370 78854
rect 285606 78618 285648 78854
rect 285328 78586 285648 78618
rect 316048 79174 316368 79206
rect 316048 78938 316090 79174
rect 316326 78938 316368 79174
rect 316048 78854 316368 78938
rect 316048 78618 316090 78854
rect 316326 78618 316368 78854
rect 316048 78586 316368 78618
rect 346768 79174 347088 79206
rect 346768 78938 346810 79174
rect 347046 78938 347088 79174
rect 346768 78854 347088 78938
rect 346768 78618 346810 78854
rect 347046 78618 347088 78854
rect 346768 78586 347088 78618
rect 54928 75454 55248 75486
rect 54928 75218 54970 75454
rect 55206 75218 55248 75454
rect 54928 75134 55248 75218
rect 54928 74898 54970 75134
rect 55206 74898 55248 75134
rect 54928 74866 55248 74898
rect 85648 75454 85968 75486
rect 85648 75218 85690 75454
rect 85926 75218 85968 75454
rect 85648 75134 85968 75218
rect 85648 74898 85690 75134
rect 85926 74898 85968 75134
rect 85648 74866 85968 74898
rect 116368 75454 116688 75486
rect 116368 75218 116410 75454
rect 116646 75218 116688 75454
rect 116368 75134 116688 75218
rect 116368 74898 116410 75134
rect 116646 74898 116688 75134
rect 116368 74866 116688 74898
rect 147088 75454 147408 75486
rect 147088 75218 147130 75454
rect 147366 75218 147408 75454
rect 147088 75134 147408 75218
rect 147088 74898 147130 75134
rect 147366 74898 147408 75134
rect 147088 74866 147408 74898
rect 177808 75454 178128 75486
rect 177808 75218 177850 75454
rect 178086 75218 178128 75454
rect 177808 75134 178128 75218
rect 177808 74898 177850 75134
rect 178086 74898 178128 75134
rect 177808 74866 178128 74898
rect 208528 75454 208848 75486
rect 208528 75218 208570 75454
rect 208806 75218 208848 75454
rect 208528 75134 208848 75218
rect 208528 74898 208570 75134
rect 208806 74898 208848 75134
rect 208528 74866 208848 74898
rect 239248 75454 239568 75486
rect 239248 75218 239290 75454
rect 239526 75218 239568 75454
rect 239248 75134 239568 75218
rect 239248 74898 239290 75134
rect 239526 74898 239568 75134
rect 239248 74866 239568 74898
rect 269968 75454 270288 75486
rect 269968 75218 270010 75454
rect 270246 75218 270288 75454
rect 269968 75134 270288 75218
rect 269968 74898 270010 75134
rect 270246 74898 270288 75134
rect 269968 74866 270288 74898
rect 300688 75454 301008 75486
rect 300688 75218 300730 75454
rect 300966 75218 301008 75454
rect 300688 75134 301008 75218
rect 300688 74898 300730 75134
rect 300966 74898 301008 75134
rect 300688 74866 301008 74898
rect 331408 75454 331728 75486
rect 331408 75218 331450 75454
rect 331686 75218 331728 75454
rect 331408 75134 331728 75218
rect 331408 74898 331450 75134
rect 331686 74898 331728 75134
rect 331408 74866 331728 74898
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 27834 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 28454 65494
rect 27834 65174 28454 65258
rect 27834 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 28454 65174
rect 22139 49604 22205 49605
rect 22139 49540 22140 49604
rect 22204 49540 22205 49604
rect 22139 49539 22205 49540
rect 22142 46613 22202 49539
rect 22139 46612 22205 46613
rect 22139 46548 22140 46612
rect 22204 46548 22205 46612
rect 22139 46547 22205 46548
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20394 -5146 21014 21498
rect 20394 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 21014 -5146
rect 20394 -5466 21014 -5382
rect 20394 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 21014 -5466
rect 20394 -7654 21014 -5702
rect 24114 25774 24734 45068
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 24114 -6106 24734 25218
rect 24114 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 24734 -6106
rect 24114 -6426 24734 -6342
rect 24114 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 24734 -6426
rect 24114 -7654 24734 -6662
rect 27834 29494 28454 64938
rect 27834 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 28454 29494
rect 27834 29174 28454 29258
rect 27834 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 28454 29174
rect 27834 -7066 28454 28938
rect 27834 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 28454 -7066
rect 27834 -7386 28454 -7302
rect 27834 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 28454 -7386
rect 27834 -7654 28454 -7622
rect 37794 39454 38414 49367
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 43174 42134 49367
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 46894 45854 49367
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 48954 14614 49574 49367
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 48954 -3226 49574 14058
rect 48954 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 49574 -3226
rect 48954 -3546 49574 -3462
rect 48954 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 49574 -3546
rect 48954 -7654 49574 -3782
rect 52674 18334 53294 49367
rect 52674 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 53294 18334
rect 52674 18014 53294 18098
rect 52674 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 53294 18014
rect 52674 -4186 53294 17778
rect 52674 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 53294 -4186
rect 52674 -4506 53294 -4422
rect 52674 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 53294 -4506
rect 52674 -7654 53294 -4742
rect 56394 22054 57014 49367
rect 56394 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 57014 22054
rect 56394 21734 57014 21818
rect 56394 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 57014 21734
rect 56394 -5146 57014 21498
rect 56394 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 57014 -5146
rect 56394 -5466 57014 -5382
rect 56394 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 57014 -5466
rect 56394 -7654 57014 -5702
rect 60114 25774 60734 49367
rect 60114 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 60734 25774
rect 60114 25454 60734 25538
rect 60114 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 60734 25454
rect 60114 -6106 60734 25218
rect 60114 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 60734 -6106
rect 60114 -6426 60734 -6342
rect 60114 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 60734 -6426
rect 60114 -7654 60734 -6662
rect 63834 29494 64454 49367
rect 63834 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 64454 29494
rect 63834 29174 64454 29258
rect 63834 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 64454 29174
rect 63834 -7066 64454 28938
rect 63834 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 64454 -7066
rect 63834 -7386 64454 -7302
rect 63834 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 64454 -7386
rect 63834 -7654 64454 -7622
rect 73794 39454 74414 49367
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 43174 78134 49367
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 46894 81854 49367
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 84954 14614 85574 49367
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 84954 -3226 85574 14058
rect 84954 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 85574 -3226
rect 84954 -3546 85574 -3462
rect 84954 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 85574 -3546
rect 84954 -7654 85574 -3782
rect 88674 18334 89294 49367
rect 88674 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 89294 18334
rect 88674 18014 89294 18098
rect 88674 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 89294 18014
rect 88674 -4186 89294 17778
rect 88674 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 89294 -4186
rect 88674 -4506 89294 -4422
rect 88674 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 89294 -4506
rect 88674 -7654 89294 -4742
rect 92394 22054 93014 49367
rect 92394 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 93014 22054
rect 92394 21734 93014 21818
rect 92394 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 93014 21734
rect 92394 -5146 93014 21498
rect 92394 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 93014 -5146
rect 92394 -5466 93014 -5382
rect 92394 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 93014 -5466
rect 92394 -7654 93014 -5702
rect 96114 25774 96734 49367
rect 96114 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 96734 25774
rect 96114 25454 96734 25538
rect 96114 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 96734 25454
rect 96114 -6106 96734 25218
rect 96114 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 96734 -6106
rect 96114 -6426 96734 -6342
rect 96114 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 96734 -6426
rect 96114 -7654 96734 -6662
rect 99834 29494 100454 49367
rect 99834 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 100454 29494
rect 99834 29174 100454 29258
rect 99834 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 100454 29174
rect 99834 -7066 100454 28938
rect 99834 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 100454 -7066
rect 99834 -7386 100454 -7302
rect 99834 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 100454 -7386
rect 99834 -7654 100454 -7622
rect 109794 39454 110414 49367
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 43174 114134 49367
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 46894 117854 49367
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 120954 14614 121574 49367
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 120954 -3226 121574 14058
rect 120954 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 121574 -3226
rect 120954 -3546 121574 -3462
rect 120954 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 121574 -3546
rect 120954 -7654 121574 -3782
rect 124674 18334 125294 49367
rect 124674 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 125294 18334
rect 124674 18014 125294 18098
rect 124674 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 125294 18014
rect 124674 -4186 125294 17778
rect 124674 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 125294 -4186
rect 124674 -4506 125294 -4422
rect 124674 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 125294 -4506
rect 124674 -7654 125294 -4742
rect 128394 22054 129014 49367
rect 128394 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 129014 22054
rect 128394 21734 129014 21818
rect 128394 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 129014 21734
rect 128394 -5146 129014 21498
rect 128394 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 129014 -5146
rect 128394 -5466 129014 -5382
rect 128394 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 129014 -5466
rect 128394 -7654 129014 -5702
rect 132114 25774 132734 49367
rect 132114 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 132734 25774
rect 132114 25454 132734 25538
rect 132114 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 132734 25454
rect 132114 -6106 132734 25218
rect 132114 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 132734 -6106
rect 132114 -6426 132734 -6342
rect 132114 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 132734 -6426
rect 132114 -7654 132734 -6662
rect 135834 29494 136454 49367
rect 135834 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 136454 29494
rect 135834 29174 136454 29258
rect 135834 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 136454 29174
rect 135834 -7066 136454 28938
rect 135834 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 136454 -7066
rect 135834 -7386 136454 -7302
rect 135834 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 136454 -7386
rect 135834 -7654 136454 -7622
rect 145794 39454 146414 49367
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 43174 150134 49367
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 46894 153854 49367
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 156954 14614 157574 49367
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 156954 -3226 157574 14058
rect 156954 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 157574 -3226
rect 156954 -3546 157574 -3462
rect 156954 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 157574 -3546
rect 156954 -7654 157574 -3782
rect 160674 18334 161294 49367
rect 160674 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 161294 18334
rect 160674 18014 161294 18098
rect 160674 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 161294 18014
rect 160674 -4186 161294 17778
rect 160674 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 161294 -4186
rect 160674 -4506 161294 -4422
rect 160674 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 161294 -4506
rect 160674 -7654 161294 -4742
rect 164394 22054 165014 49367
rect 164394 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 165014 22054
rect 164394 21734 165014 21818
rect 164394 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 165014 21734
rect 164394 -5146 165014 21498
rect 164394 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 165014 -5146
rect 164394 -5466 165014 -5382
rect 164394 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 165014 -5466
rect 164394 -7654 165014 -5702
rect 168114 25774 168734 49367
rect 168114 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 168734 25774
rect 168114 25454 168734 25538
rect 168114 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 168734 25454
rect 168114 -6106 168734 25218
rect 168114 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 168734 -6106
rect 168114 -6426 168734 -6342
rect 168114 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 168734 -6426
rect 168114 -7654 168734 -6662
rect 171834 29494 172454 49367
rect 171834 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 172454 29494
rect 171834 29174 172454 29258
rect 171834 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 172454 29174
rect 171834 -7066 172454 28938
rect 171834 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 172454 -7066
rect 171834 -7386 172454 -7302
rect 171834 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 172454 -7386
rect 171834 -7654 172454 -7622
rect 181794 39454 182414 49367
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 43174 186134 49367
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 46894 189854 49367
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 192954 14614 193574 45068
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 192954 -3226 193574 14058
rect 192954 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 193574 -3226
rect 192954 -3546 193574 -3462
rect 192954 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 193574 -3546
rect 192954 -7654 193574 -3782
rect 196674 18334 197294 49367
rect 196674 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 197294 18334
rect 196674 18014 197294 18098
rect 196674 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 197294 18014
rect 196674 -4186 197294 17778
rect 196674 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 197294 -4186
rect 196674 -4506 197294 -4422
rect 196674 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 197294 -4506
rect 196674 -7654 197294 -4742
rect 200394 22054 201014 49367
rect 200394 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 201014 22054
rect 200394 21734 201014 21818
rect 200394 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 201014 21734
rect 200394 -5146 201014 21498
rect 200394 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 201014 -5146
rect 200394 -5466 201014 -5382
rect 200394 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 201014 -5466
rect 200394 -7654 201014 -5702
rect 204114 25774 204734 49367
rect 204114 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 204734 25774
rect 204114 25454 204734 25538
rect 204114 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 204734 25454
rect 204114 -6106 204734 25218
rect 204114 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 204734 -6106
rect 204114 -6426 204734 -6342
rect 204114 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 204734 -6426
rect 204114 -7654 204734 -6662
rect 207834 29494 208454 49367
rect 207834 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 208454 29494
rect 207834 29174 208454 29258
rect 207834 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 208454 29174
rect 207834 -7066 208454 28938
rect 207834 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 208454 -7066
rect 207834 -7386 208454 -7302
rect 207834 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 208454 -7386
rect 207834 -7654 208454 -7622
rect 217794 39454 218414 49367
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 43174 222134 49367
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 46894 225854 49367
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 228954 14614 229574 49367
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228954 -3226 229574 14058
rect 228954 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 229574 -3226
rect 228954 -3546 229574 -3462
rect 228954 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 229574 -3546
rect 228954 -7654 229574 -3782
rect 232674 18334 233294 49367
rect 232674 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 233294 18334
rect 232674 18014 233294 18098
rect 232674 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 233294 18014
rect 232674 -4186 233294 17778
rect 232674 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 233294 -4186
rect 232674 -4506 233294 -4422
rect 232674 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 233294 -4506
rect 232674 -7654 233294 -4742
rect 236394 22054 237014 49367
rect 236394 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 237014 22054
rect 236394 21734 237014 21818
rect 236394 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 237014 21734
rect 236394 -5146 237014 21498
rect 236394 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 237014 -5146
rect 236394 -5466 237014 -5382
rect 236394 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 237014 -5466
rect 236394 -7654 237014 -5702
rect 240114 25774 240734 49367
rect 240114 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 240734 25774
rect 240114 25454 240734 25538
rect 240114 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 240734 25454
rect 240114 -6106 240734 25218
rect 240114 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 240734 -6106
rect 240114 -6426 240734 -6342
rect 240114 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 240734 -6426
rect 240114 -7654 240734 -6662
rect 243834 29494 244454 49367
rect 243834 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 244454 29494
rect 243834 29174 244454 29258
rect 243834 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 244454 29174
rect 243834 -7066 244454 28938
rect 243834 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 244454 -7066
rect 243834 -7386 244454 -7302
rect 243834 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 244454 -7386
rect 243834 -7654 244454 -7622
rect 253794 39454 254414 49367
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 43174 258134 49367
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 46894 261854 49367
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -2266 261854 10338
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 264954 14614 265574 49367
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 264954 -3226 265574 14058
rect 264954 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 265574 -3226
rect 264954 -3546 265574 -3462
rect 264954 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 265574 -3546
rect 264954 -7654 265574 -3782
rect 268674 18334 269294 49367
rect 268674 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 269294 18334
rect 268674 18014 269294 18098
rect 268674 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 269294 18014
rect 268674 -4186 269294 17778
rect 268674 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 269294 -4186
rect 268674 -4506 269294 -4422
rect 268674 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 269294 -4506
rect 268674 -7654 269294 -4742
rect 272394 22054 273014 49367
rect 272394 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 273014 22054
rect 272394 21734 273014 21818
rect 272394 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 273014 21734
rect 272394 -5146 273014 21498
rect 272394 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 273014 -5146
rect 272394 -5466 273014 -5382
rect 272394 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 273014 -5466
rect 272394 -7654 273014 -5702
rect 276114 25774 276734 49367
rect 276114 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 276734 25774
rect 276114 25454 276734 25538
rect 276114 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 276734 25454
rect 276114 -6106 276734 25218
rect 276114 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 276734 -6106
rect 276114 -6426 276734 -6342
rect 276114 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 276734 -6426
rect 276114 -7654 276734 -6662
rect 279834 29494 280454 49367
rect 279834 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 280454 29494
rect 279834 29174 280454 29258
rect 279834 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 280454 29174
rect 279834 -7066 280454 28938
rect 279834 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 280454 -7066
rect 279834 -7386 280454 -7302
rect 279834 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 280454 -7386
rect 279834 -7654 280454 -7622
rect 289794 39454 290414 49367
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 43174 294134 49367
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 46894 297854 49367
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 300954 14614 301574 45068
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 300954 -3226 301574 14058
rect 300954 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 301574 -3226
rect 300954 -3546 301574 -3462
rect 300954 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 301574 -3546
rect 300954 -7654 301574 -3782
rect 304674 18334 305294 49367
rect 304674 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 305294 18334
rect 304674 18014 305294 18098
rect 304674 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 305294 18014
rect 304674 -4186 305294 17778
rect 304674 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 305294 -4186
rect 304674 -4506 305294 -4422
rect 304674 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 305294 -4506
rect 304674 -7654 305294 -4742
rect 308394 22054 309014 49367
rect 308394 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 309014 22054
rect 308394 21734 309014 21818
rect 308394 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 309014 21734
rect 308394 -5146 309014 21498
rect 308394 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 309014 -5146
rect 308394 -5466 309014 -5382
rect 308394 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 309014 -5466
rect 308394 -7654 309014 -5702
rect 312114 25774 312734 49367
rect 312114 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 312734 25774
rect 312114 25454 312734 25538
rect 312114 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 312734 25454
rect 312114 -6106 312734 25218
rect 312114 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 312734 -6106
rect 312114 -6426 312734 -6342
rect 312114 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 312734 -6426
rect 312114 -7654 312734 -6662
rect 315834 29494 316454 45068
rect 315834 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 316454 29494
rect 315834 29174 316454 29258
rect 315834 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 316454 29174
rect 315834 -7066 316454 28938
rect 315834 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 316454 -7066
rect 315834 -7386 316454 -7302
rect 315834 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 316454 -7386
rect 315834 -7654 316454 -7622
rect 325794 39454 326414 49367
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 43174 330134 49367
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 46894 333854 49367
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 336954 14614 337574 49367
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 336954 -3226 337574 14058
rect 336954 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 337574 -3226
rect 336954 -3546 337574 -3462
rect 336954 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 337574 -3546
rect 336954 -7654 337574 -3782
rect 340674 18334 341294 49367
rect 340674 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 341294 18334
rect 340674 18014 341294 18098
rect 340674 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 341294 18014
rect 340674 -4186 341294 17778
rect 340674 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 341294 -4186
rect 340674 -4506 341294 -4422
rect 340674 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 341294 -4506
rect 340674 -7654 341294 -4742
rect 344394 22054 345014 49367
rect 344394 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 345014 22054
rect 344394 21734 345014 21818
rect 344394 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 345014 21734
rect 344394 -5146 345014 21498
rect 344394 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 345014 -5146
rect 344394 -5466 345014 -5382
rect 344394 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 345014 -5466
rect 344394 -7654 345014 -5702
rect 348114 25774 348734 49367
rect 348114 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 348734 25774
rect 348114 25454 348734 25538
rect 348114 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 348734 25454
rect 348114 -6106 348734 25218
rect 348114 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 348734 -6106
rect 348114 -6426 348734 -6342
rect 348114 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 348734 -6426
rect 348114 -7654 348734 -6662
rect 351834 29494 352454 49367
rect 351834 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 352454 29494
rect 351834 29174 352454 29258
rect 351834 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 352454 29174
rect 351834 -7066 352454 28938
rect 351834 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 352454 -7066
rect 351834 -7386 352454 -7302
rect 351834 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 352454 -7386
rect 351834 -7654 352454 -7622
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 372954 -3226 373574 14058
rect 372954 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 373574 -3226
rect 372954 -3546 373574 -3462
rect 372954 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 373574 -3546
rect 372954 -7654 373574 -3782
rect 376674 708678 377294 711590
rect 376674 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 377294 708678
rect 376674 708358 377294 708442
rect 376674 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 377294 708358
rect 376674 666334 377294 708122
rect 376674 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 377294 666334
rect 376674 666014 377294 666098
rect 376674 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 377294 666014
rect 376674 630334 377294 665778
rect 376674 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 377294 630334
rect 376674 630014 377294 630098
rect 376674 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 377294 630014
rect 376674 594334 377294 629778
rect 376674 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 377294 594334
rect 376674 594014 377294 594098
rect 376674 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 377294 594014
rect 376674 558334 377294 593778
rect 376674 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 377294 558334
rect 376674 558014 377294 558098
rect 376674 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 377294 558014
rect 376674 522334 377294 557778
rect 376674 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 377294 522334
rect 376674 522014 377294 522098
rect 376674 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 377294 522014
rect 376674 486334 377294 521778
rect 376674 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 377294 486334
rect 376674 486014 377294 486098
rect 376674 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 377294 486014
rect 376674 450334 377294 485778
rect 376674 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 377294 450334
rect 376674 450014 377294 450098
rect 376674 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 377294 450014
rect 376674 414334 377294 449778
rect 376674 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 377294 414334
rect 376674 414014 377294 414098
rect 376674 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 377294 414014
rect 376674 378334 377294 413778
rect 376674 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 377294 378334
rect 376674 378014 377294 378098
rect 376674 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 377294 378014
rect 376674 342334 377294 377778
rect 376674 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 377294 342334
rect 376674 342014 377294 342098
rect 376674 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 377294 342014
rect 376674 306334 377294 341778
rect 376674 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 377294 306334
rect 376674 306014 377294 306098
rect 376674 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 377294 306014
rect 376674 270334 377294 305778
rect 376674 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 377294 270334
rect 376674 270014 377294 270098
rect 376674 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 377294 270014
rect 376674 234334 377294 269778
rect 376674 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 377294 234334
rect 376674 234014 377294 234098
rect 376674 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 377294 234014
rect 376674 198334 377294 233778
rect 376674 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 377294 198334
rect 376674 198014 377294 198098
rect 376674 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 377294 198014
rect 376674 162334 377294 197778
rect 376674 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 377294 162334
rect 376674 162014 377294 162098
rect 376674 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 377294 162014
rect 376674 126334 377294 161778
rect 376674 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 377294 126334
rect 376674 126014 377294 126098
rect 376674 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 377294 126014
rect 376674 90334 377294 125778
rect 376674 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 377294 90334
rect 376674 90014 377294 90098
rect 376674 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 377294 90014
rect 376674 54334 377294 89778
rect 376674 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 377294 54334
rect 376674 54014 377294 54098
rect 376674 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 377294 54014
rect 376674 18334 377294 53778
rect 376674 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 377294 18334
rect 376674 18014 377294 18098
rect 376674 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 377294 18014
rect 376674 -4186 377294 17778
rect 376674 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 377294 -4186
rect 376674 -4506 377294 -4422
rect 376674 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 377294 -4506
rect 376674 -7654 377294 -4742
rect 380394 709638 381014 711590
rect 380394 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 381014 709638
rect 380394 709318 381014 709402
rect 380394 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 381014 709318
rect 380394 670054 381014 709082
rect 380394 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 381014 670054
rect 380394 669734 381014 669818
rect 380394 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 381014 669734
rect 380394 634054 381014 669498
rect 380394 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 381014 634054
rect 380394 633734 381014 633818
rect 380394 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 381014 633734
rect 380394 598054 381014 633498
rect 380394 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 381014 598054
rect 380394 597734 381014 597818
rect 380394 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 381014 597734
rect 380394 562054 381014 597498
rect 380394 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 381014 562054
rect 380394 561734 381014 561818
rect 380394 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 381014 561734
rect 380394 526054 381014 561498
rect 380394 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 381014 526054
rect 380394 525734 381014 525818
rect 380394 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 381014 525734
rect 380394 490054 381014 525498
rect 380394 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 381014 490054
rect 380394 489734 381014 489818
rect 380394 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 381014 489734
rect 380394 454054 381014 489498
rect 380394 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 381014 454054
rect 380394 453734 381014 453818
rect 380394 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 381014 453734
rect 380394 418054 381014 453498
rect 380394 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 381014 418054
rect 380394 417734 381014 417818
rect 380394 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 381014 417734
rect 380394 382054 381014 417498
rect 380394 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 381014 382054
rect 380394 381734 381014 381818
rect 380394 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 381014 381734
rect 380394 346054 381014 381498
rect 380394 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 381014 346054
rect 380394 345734 381014 345818
rect 380394 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 381014 345734
rect 380394 310054 381014 345498
rect 380394 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 381014 310054
rect 380394 309734 381014 309818
rect 380394 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 381014 309734
rect 380394 274054 381014 309498
rect 380394 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 381014 274054
rect 380394 273734 381014 273818
rect 380394 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 381014 273734
rect 380394 238054 381014 273498
rect 380394 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 381014 238054
rect 380394 237734 381014 237818
rect 380394 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 381014 237734
rect 380394 202054 381014 237498
rect 380394 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 381014 202054
rect 380394 201734 381014 201818
rect 380394 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 381014 201734
rect 380394 166054 381014 201498
rect 380394 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 381014 166054
rect 380394 165734 381014 165818
rect 380394 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 381014 165734
rect 380394 130054 381014 165498
rect 380394 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 381014 130054
rect 380394 129734 381014 129818
rect 380394 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 381014 129734
rect 380394 94054 381014 129498
rect 380394 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 381014 94054
rect 380394 93734 381014 93818
rect 380394 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 381014 93734
rect 380394 58054 381014 93498
rect 380394 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 381014 58054
rect 380394 57734 381014 57818
rect 380394 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 381014 57734
rect 380394 22054 381014 57498
rect 380394 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 381014 22054
rect 380394 21734 381014 21818
rect 380394 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 381014 21734
rect 380394 -5146 381014 21498
rect 380394 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 381014 -5146
rect 380394 -5466 381014 -5382
rect 380394 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 381014 -5466
rect 380394 -7654 381014 -5702
rect 384114 710598 384734 711590
rect 384114 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 384734 710598
rect 384114 710278 384734 710362
rect 384114 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 384734 710278
rect 384114 673774 384734 710042
rect 384114 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 384734 673774
rect 384114 673454 384734 673538
rect 384114 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 384734 673454
rect 384114 637774 384734 673218
rect 384114 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 384734 637774
rect 384114 637454 384734 637538
rect 384114 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 384734 637454
rect 384114 601774 384734 637218
rect 384114 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 384734 601774
rect 384114 601454 384734 601538
rect 384114 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 384734 601454
rect 384114 565774 384734 601218
rect 384114 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 384734 565774
rect 384114 565454 384734 565538
rect 384114 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 384734 565454
rect 384114 529774 384734 565218
rect 384114 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 384734 529774
rect 384114 529454 384734 529538
rect 384114 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 384734 529454
rect 384114 493774 384734 529218
rect 384114 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 384734 493774
rect 384114 493454 384734 493538
rect 384114 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 384734 493454
rect 384114 457774 384734 493218
rect 384114 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 384734 457774
rect 384114 457454 384734 457538
rect 384114 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 384734 457454
rect 384114 421774 384734 457218
rect 384114 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 384734 421774
rect 384114 421454 384734 421538
rect 384114 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 384734 421454
rect 384114 385774 384734 421218
rect 384114 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 384734 385774
rect 384114 385454 384734 385538
rect 384114 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 384734 385454
rect 384114 349774 384734 385218
rect 384114 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 384734 349774
rect 384114 349454 384734 349538
rect 384114 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 384734 349454
rect 384114 313774 384734 349218
rect 384114 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 384734 313774
rect 384114 313454 384734 313538
rect 384114 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 384734 313454
rect 384114 277774 384734 313218
rect 384114 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 384734 277774
rect 384114 277454 384734 277538
rect 384114 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 384734 277454
rect 384114 241774 384734 277218
rect 384114 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 384734 241774
rect 384114 241454 384734 241538
rect 384114 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 384734 241454
rect 384114 205774 384734 241218
rect 384114 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 384734 205774
rect 384114 205454 384734 205538
rect 384114 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 384734 205454
rect 384114 169774 384734 205218
rect 384114 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 384734 169774
rect 384114 169454 384734 169538
rect 384114 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 384734 169454
rect 384114 133774 384734 169218
rect 384114 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 384734 133774
rect 384114 133454 384734 133538
rect 384114 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 384734 133454
rect 384114 97774 384734 133218
rect 384114 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 384734 97774
rect 384114 97454 384734 97538
rect 384114 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 384734 97454
rect 384114 61774 384734 97218
rect 387834 711558 388454 711590
rect 387834 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 388454 711558
rect 387834 711238 388454 711322
rect 387834 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 388454 711238
rect 387834 677494 388454 711002
rect 387834 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 388454 677494
rect 387834 677174 388454 677258
rect 387834 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 388454 677174
rect 387834 641494 388454 676938
rect 387834 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 388454 641494
rect 387834 641174 388454 641258
rect 387834 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 388454 641174
rect 387834 605494 388454 640938
rect 387834 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 388454 605494
rect 387834 605174 388454 605258
rect 387834 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 388454 605174
rect 387834 569494 388454 604938
rect 387834 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 388454 569494
rect 387834 569174 388454 569258
rect 387834 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 388454 569174
rect 387834 533494 388454 568938
rect 387834 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 388454 533494
rect 387834 533174 388454 533258
rect 387834 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 388454 533174
rect 387834 497494 388454 532938
rect 387834 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 388454 497494
rect 387834 497174 388454 497258
rect 387834 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 388454 497174
rect 387834 461494 388454 496938
rect 387834 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 388454 461494
rect 387834 461174 388454 461258
rect 387834 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 388454 461174
rect 387834 425494 388454 460938
rect 387834 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 388454 425494
rect 387834 425174 388454 425258
rect 387834 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 388454 425174
rect 387834 389494 388454 424938
rect 387834 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 388454 389494
rect 387834 389174 388454 389258
rect 387834 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 388454 389174
rect 387834 353494 388454 388938
rect 387834 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 388454 353494
rect 387834 353174 388454 353258
rect 387834 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 388454 353174
rect 387834 317494 388454 352938
rect 387834 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 388454 317494
rect 387834 317174 388454 317258
rect 387834 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 388454 317174
rect 387834 281494 388454 316938
rect 387834 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 388454 281494
rect 387834 281174 388454 281258
rect 387834 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 388454 281174
rect 387834 245494 388454 280938
rect 387834 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 388454 245494
rect 387834 245174 388454 245258
rect 387834 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 388454 245174
rect 387834 209494 388454 244938
rect 387834 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 388454 209494
rect 387834 209174 388454 209258
rect 387834 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 388454 209174
rect 387834 173494 388454 208938
rect 387834 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 388454 173494
rect 387834 173174 388454 173258
rect 387834 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 388454 173174
rect 387834 137494 388454 172938
rect 387834 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 388454 137494
rect 387834 137174 388454 137258
rect 387834 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 388454 137174
rect 387834 101494 388454 136938
rect 387834 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 388454 101494
rect 387834 101174 388454 101258
rect 387834 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 388454 101174
rect 387834 92137 388454 100938
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 92137 398414 110898
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 404417 327454 404737 327486
rect 404417 327218 404459 327454
rect 404695 327218 404737 327454
rect 404417 327134 404737 327218
rect 404417 326898 404459 327134
rect 404695 326898 404737 327134
rect 404417 326866 404737 326898
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 92137 402134 114618
rect 405234 298894 405854 334338
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 407890 331174 408210 331206
rect 407890 330938 407932 331174
rect 408168 330938 408210 331174
rect 407890 330854 408210 330938
rect 407890 330618 407932 330854
rect 408168 330618 408210 330854
rect 407890 330586 408210 330618
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 104460 405854 118338
rect 408954 302614 409574 338058
rect 412674 708678 413294 711590
rect 412674 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 413294 708678
rect 412674 708358 413294 708442
rect 412674 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 413294 708358
rect 412674 666334 413294 708122
rect 412674 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 413294 666334
rect 412674 666014 413294 666098
rect 412674 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 413294 666014
rect 412674 630334 413294 665778
rect 412674 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 413294 630334
rect 412674 630014 413294 630098
rect 412674 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 413294 630014
rect 412674 594334 413294 629778
rect 412674 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 413294 594334
rect 412674 594014 413294 594098
rect 412674 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 413294 594014
rect 412674 558334 413294 593778
rect 412674 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 413294 558334
rect 412674 558014 413294 558098
rect 412674 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 413294 558014
rect 412674 522334 413294 557778
rect 412674 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 413294 522334
rect 412674 522014 413294 522098
rect 412674 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 413294 522014
rect 412674 486334 413294 521778
rect 412674 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 413294 486334
rect 412674 486014 413294 486098
rect 412674 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 413294 486014
rect 412674 450334 413294 485778
rect 412674 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 413294 450334
rect 412674 450014 413294 450098
rect 412674 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 413294 450014
rect 412674 414334 413294 449778
rect 412674 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 413294 414334
rect 412674 414014 413294 414098
rect 412674 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 413294 414014
rect 412674 378334 413294 413778
rect 412674 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 413294 378334
rect 412674 378014 413294 378098
rect 412674 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 413294 378014
rect 412674 342334 413294 377778
rect 412674 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 413294 342334
rect 412674 342014 413294 342098
rect 412674 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 413294 342014
rect 411363 327454 411683 327486
rect 411363 327218 411405 327454
rect 411641 327218 411683 327454
rect 411363 327134 411683 327218
rect 411363 326898 411405 327134
rect 411641 326898 411683 327134
rect 411363 326866 411683 326898
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 92137 409574 122058
rect 412674 306334 413294 341778
rect 416394 709638 417014 711590
rect 416394 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 417014 709638
rect 416394 709318 417014 709402
rect 416394 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 417014 709318
rect 416394 670054 417014 709082
rect 416394 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 417014 670054
rect 416394 669734 417014 669818
rect 416394 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 417014 669734
rect 416394 634054 417014 669498
rect 416394 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 417014 634054
rect 416394 633734 417014 633818
rect 416394 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 417014 633734
rect 416394 598054 417014 633498
rect 416394 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 417014 598054
rect 416394 597734 417014 597818
rect 416394 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 417014 597734
rect 416394 562054 417014 597498
rect 416394 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 417014 562054
rect 416394 561734 417014 561818
rect 416394 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 417014 561734
rect 416394 526054 417014 561498
rect 416394 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 417014 526054
rect 416394 525734 417014 525818
rect 416394 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 417014 525734
rect 416394 490054 417014 525498
rect 416394 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 417014 490054
rect 416394 489734 417014 489818
rect 416394 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 417014 489734
rect 416394 454054 417014 489498
rect 416394 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 417014 454054
rect 416394 453734 417014 453818
rect 416394 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 417014 453734
rect 416394 418054 417014 453498
rect 416394 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 417014 418054
rect 416394 417734 417014 417818
rect 416394 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 417014 417734
rect 416394 382054 417014 417498
rect 416394 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 417014 382054
rect 416394 381734 417014 381818
rect 416394 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 417014 381734
rect 416394 346054 417014 381498
rect 416394 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 417014 346054
rect 416394 345734 417014 345818
rect 416394 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 417014 345734
rect 414836 331174 415156 331206
rect 414836 330938 414878 331174
rect 415114 330938 415156 331174
rect 414836 330854 415156 330938
rect 414836 330618 414878 330854
rect 415114 330618 415156 330854
rect 414836 330586 415156 330618
rect 412674 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 413294 306334
rect 412674 306014 413294 306098
rect 412674 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 413294 306014
rect 412674 270334 413294 305778
rect 412674 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 413294 270334
rect 412674 270014 413294 270098
rect 412674 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 413294 270014
rect 412674 234334 413294 269778
rect 412674 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 413294 234334
rect 412674 234014 413294 234098
rect 412674 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 413294 234014
rect 412674 198334 413294 233778
rect 412674 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 413294 198334
rect 412674 198014 413294 198098
rect 412674 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 413294 198014
rect 412674 162334 413294 197778
rect 412674 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 413294 162334
rect 412674 162014 413294 162098
rect 412674 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 413294 162014
rect 412674 126334 413294 161778
rect 416394 310054 417014 345498
rect 420114 710598 420734 711590
rect 420114 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 420734 710598
rect 420114 710278 420734 710362
rect 420114 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 420734 710278
rect 420114 673774 420734 710042
rect 420114 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 420734 673774
rect 420114 673454 420734 673538
rect 420114 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 420734 673454
rect 420114 637774 420734 673218
rect 420114 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 420734 637774
rect 420114 637454 420734 637538
rect 420114 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 420734 637454
rect 420114 601774 420734 637218
rect 420114 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 420734 601774
rect 420114 601454 420734 601538
rect 420114 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 420734 601454
rect 420114 565774 420734 601218
rect 420114 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 420734 565774
rect 420114 565454 420734 565538
rect 420114 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 420734 565454
rect 420114 529774 420734 565218
rect 420114 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 420734 529774
rect 420114 529454 420734 529538
rect 420114 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 420734 529454
rect 420114 493774 420734 529218
rect 420114 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 420734 493774
rect 420114 493454 420734 493538
rect 420114 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 420734 493454
rect 420114 457774 420734 493218
rect 420114 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 420734 457774
rect 420114 457454 420734 457538
rect 420114 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 420734 457454
rect 420114 421774 420734 457218
rect 423834 711558 424454 711590
rect 423834 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 424454 711558
rect 423834 711238 424454 711322
rect 423834 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 424454 711238
rect 423834 677494 424454 711002
rect 423834 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 424454 677494
rect 423834 677174 424454 677258
rect 423834 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 424454 677174
rect 423834 641494 424454 676938
rect 423834 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 424454 641494
rect 423834 641174 424454 641258
rect 423834 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 424454 641174
rect 423834 605494 424454 640938
rect 423834 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 424454 605494
rect 423834 605174 424454 605258
rect 423834 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 424454 605174
rect 423834 569494 424454 604938
rect 423834 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 424454 569494
rect 423834 569174 424454 569258
rect 423834 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 424454 569174
rect 423834 533494 424454 568938
rect 423834 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 424454 533494
rect 423834 533174 424454 533258
rect 423834 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 424454 533174
rect 423834 497494 424454 532938
rect 423834 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 424454 497494
rect 423834 497174 424454 497258
rect 423834 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 424454 497174
rect 423834 461494 424454 496938
rect 423834 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 424454 461494
rect 423834 461174 424454 461258
rect 423834 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 424454 461174
rect 423834 444412 424454 460938
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 442833 434414 470898
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 444412 438134 474618
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444235 700364 444301 700365
rect 444235 700300 444236 700364
rect 444300 700300 444301 700364
rect 444235 700299 444301 700300
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442833 441854 478338
rect 426624 439174 426944 439206
rect 426624 438938 426666 439174
rect 426902 438938 426944 439174
rect 426624 438854 426944 438938
rect 426624 438618 426666 438854
rect 426902 438618 426944 438854
rect 426624 438586 426944 438618
rect 432305 439174 432625 439206
rect 432305 438938 432347 439174
rect 432583 438938 432625 439174
rect 432305 438854 432625 438938
rect 432305 438618 432347 438854
rect 432583 438618 432625 438854
rect 432305 438586 432625 438618
rect 437986 439174 438306 439206
rect 437986 438938 438028 439174
rect 438264 438938 438306 439174
rect 437986 438854 438306 438938
rect 437986 438618 438028 438854
rect 438264 438618 438306 438854
rect 437986 438586 438306 438618
rect 443667 439174 443987 439206
rect 443667 438938 443709 439174
rect 443945 438938 443987 439174
rect 443667 438854 443987 438938
rect 443667 438618 443709 438854
rect 443945 438618 443987 438854
rect 443667 438586 443987 438618
rect 423784 435454 424104 435486
rect 423784 435218 423826 435454
rect 424062 435218 424104 435454
rect 423784 435134 424104 435218
rect 423784 434898 423826 435134
rect 424062 434898 424104 435134
rect 423784 434866 424104 434898
rect 429465 435454 429785 435486
rect 429465 435218 429507 435454
rect 429743 435218 429785 435454
rect 429465 435134 429785 435218
rect 429465 434898 429507 435134
rect 429743 434898 429785 435134
rect 429465 434866 429785 434898
rect 435146 435454 435466 435486
rect 435146 435218 435188 435454
rect 435424 435218 435466 435454
rect 435146 435134 435466 435218
rect 435146 434898 435188 435134
rect 435424 434898 435466 435134
rect 435146 434866 435466 434898
rect 440827 435454 441147 435486
rect 440827 435218 440869 435454
rect 441105 435218 441147 435454
rect 440827 435134 441147 435218
rect 440827 434898 440869 435134
rect 441105 434898 441147 435134
rect 440827 434866 441147 434898
rect 420114 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 420734 421774
rect 420114 421454 420734 421538
rect 420114 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 420734 421454
rect 420114 385774 420734 421218
rect 420114 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 420734 385774
rect 420114 385454 420734 385538
rect 420114 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 420734 385454
rect 420114 349774 420734 385218
rect 420114 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 420734 349774
rect 420114 349454 420734 349538
rect 420114 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 420734 349454
rect 418309 327454 418629 327486
rect 418309 327218 418351 327454
rect 418587 327218 418629 327454
rect 418309 327134 418629 327218
rect 418309 326898 418351 327134
rect 418587 326898 418629 327134
rect 418309 326866 418629 326898
rect 416394 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 417014 310054
rect 416394 309734 417014 309818
rect 416394 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 417014 309734
rect 416394 274054 417014 309498
rect 416394 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 417014 274054
rect 416394 273734 417014 273818
rect 416394 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 417014 273734
rect 416394 238054 417014 273498
rect 416394 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 417014 238054
rect 416394 237734 417014 237818
rect 416394 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 417014 237734
rect 416394 202054 417014 237498
rect 416394 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 417014 202054
rect 416394 201734 417014 201818
rect 416394 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 417014 201734
rect 416394 166054 417014 201498
rect 416394 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 417014 166054
rect 416394 165734 417014 165818
rect 416394 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 417014 165734
rect 416394 157249 417014 165498
rect 420114 313774 420734 349218
rect 423834 389494 424454 420068
rect 423834 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 424454 389494
rect 423834 389174 424454 389258
rect 423834 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 424454 389174
rect 423834 353494 424454 388938
rect 423834 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 424454 353494
rect 423834 353174 424454 353258
rect 423834 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 424454 353174
rect 421419 334116 421485 334117
rect 421419 334052 421420 334116
rect 421484 334052 421485 334116
rect 421419 334051 421485 334052
rect 420114 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 420734 313774
rect 420114 313454 420734 313538
rect 420114 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 420734 313454
rect 420114 277774 420734 313218
rect 420114 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 420734 277774
rect 420114 277454 420734 277538
rect 420114 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 420734 277454
rect 420114 241774 420734 277218
rect 420114 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 420734 241774
rect 420114 241454 420734 241538
rect 420114 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 420734 241454
rect 420114 205774 420734 241218
rect 420114 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 420734 205774
rect 420114 205454 420734 205538
rect 420114 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 420734 205454
rect 420114 169774 420734 205218
rect 420114 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 420734 169774
rect 420114 169454 420734 169538
rect 420114 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 420734 169454
rect 420114 157249 420734 169218
rect 421422 162757 421482 334051
rect 421782 331174 422102 331206
rect 421782 330938 421824 331174
rect 422060 330938 422102 331174
rect 421782 330854 422102 330938
rect 421782 330618 421824 330854
rect 422060 330618 422102 330854
rect 421782 330586 422102 330618
rect 423834 317494 424454 352938
rect 433794 399454 434414 422599
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 428411 336836 428477 336837
rect 428411 336772 428412 336836
rect 428476 336772 428477 336836
rect 428411 336771 428477 336772
rect 425835 334388 425901 334389
rect 425835 334324 425836 334388
rect 425900 334324 425901 334388
rect 425835 334323 425901 334324
rect 425255 327454 425575 327486
rect 425255 327218 425297 327454
rect 425533 327218 425575 327454
rect 425255 327134 425575 327218
rect 425255 326898 425297 327134
rect 425533 326898 425575 327134
rect 425255 326866 425575 326898
rect 423834 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 424454 317494
rect 423834 317174 424454 317258
rect 423834 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 424454 317174
rect 423834 281494 424454 316938
rect 423834 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 424454 281494
rect 423834 281174 424454 281258
rect 423834 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 424454 281174
rect 423834 245494 424454 280938
rect 423834 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 424454 245494
rect 423834 245174 424454 245258
rect 423834 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 424454 245174
rect 423834 209494 424454 244938
rect 423834 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 424454 209494
rect 423834 209174 424454 209258
rect 423834 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 424454 209174
rect 423834 173494 424454 208938
rect 423834 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 424454 173494
rect 423834 173174 424454 173258
rect 423834 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 424454 173174
rect 421419 162756 421485 162757
rect 421419 162692 421420 162756
rect 421484 162692 421485 162756
rect 421419 162691 421485 162692
rect 423834 157249 424454 172938
rect 425838 162757 425898 334323
rect 428414 162757 428474 336771
rect 428728 331174 429048 331206
rect 428728 330938 428770 331174
rect 429006 330938 429048 331174
rect 428728 330854 429048 330938
rect 428728 330618 428770 330854
rect 429006 330618 429048 330854
rect 428728 330586 429048 330618
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 425835 162756 425901 162757
rect 425835 162692 425836 162756
rect 425900 162692 425901 162756
rect 425835 162691 425901 162692
rect 428411 162756 428477 162757
rect 428411 162692 428412 162756
rect 428476 162692 428477 162756
rect 428411 162691 428477 162692
rect 433794 157249 434414 182898
rect 437514 403174 438134 420068
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 157249 438134 186618
rect 441234 406894 441854 422599
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 444238 321061 444298 700299
rect 444954 698614 445574 707162
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 448674 708678 449294 711590
rect 448674 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 449294 708678
rect 448674 708358 449294 708442
rect 448674 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 449294 708358
rect 447731 692068 447797 692069
rect 447731 692004 447732 692068
rect 447796 692004 447797 692068
rect 447731 692003 447797 692004
rect 446259 689348 446325 689349
rect 446259 689284 446260 689348
rect 446324 689284 446325 689348
rect 446259 689283 446325 689284
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444235 321060 444301 321061
rect 444235 320996 444236 321060
rect 444300 320996 444301 321060
rect 444235 320995 444301 320996
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 157249 441854 190338
rect 444954 302614 445574 338058
rect 446262 319973 446322 689283
rect 446259 319972 446325 319973
rect 446259 319908 446260 319972
rect 446324 319908 446325 319972
rect 446259 319907 446325 319908
rect 447734 319701 447794 692003
rect 447915 684316 447981 684317
rect 447915 684252 447916 684316
rect 447980 684252 447981 684316
rect 447915 684251 447981 684252
rect 447918 321333 447978 684251
rect 448674 666334 449294 708122
rect 452394 709638 453014 711590
rect 452394 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 453014 709638
rect 452394 709318 453014 709402
rect 452394 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 453014 709318
rect 449571 700500 449637 700501
rect 449571 700436 449572 700500
rect 449636 700436 449637 700500
rect 449571 700435 449637 700436
rect 448674 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 449294 666334
rect 448674 666014 449294 666098
rect 448674 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 449294 666014
rect 448674 630334 449294 665778
rect 448674 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 449294 630334
rect 448674 630014 449294 630098
rect 448674 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 449294 630014
rect 448674 594334 449294 629778
rect 448674 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 449294 594334
rect 448674 594014 449294 594098
rect 448674 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 449294 594014
rect 448674 558334 449294 593778
rect 448674 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 449294 558334
rect 448674 558014 449294 558098
rect 448674 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 449294 558014
rect 448674 522334 449294 557778
rect 448674 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 449294 522334
rect 448674 522014 449294 522098
rect 448674 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 449294 522014
rect 448674 486334 449294 521778
rect 448674 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 449294 486334
rect 448674 486014 449294 486098
rect 448674 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 449294 486014
rect 448674 450334 449294 485778
rect 448674 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 449294 450334
rect 448674 450014 449294 450098
rect 448674 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 449294 450014
rect 448674 414334 449294 449778
rect 448674 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 449294 414334
rect 448674 414014 449294 414098
rect 448674 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 449294 414014
rect 448283 395316 448349 395317
rect 448283 395252 448284 395316
rect 448348 395252 448349 395316
rect 448283 395251 448349 395252
rect 448286 346221 448346 395251
rect 448674 378334 449294 413778
rect 448674 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 449294 378334
rect 448674 378014 449294 378098
rect 448674 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 449294 378014
rect 448283 346220 448349 346221
rect 448283 346156 448284 346220
rect 448348 346156 448349 346220
rect 448283 346155 448349 346156
rect 448674 342334 449294 377778
rect 448674 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 449294 342334
rect 448674 342014 449294 342098
rect 448674 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 449294 342014
rect 447915 321332 447981 321333
rect 447915 321268 447916 321332
rect 447980 321268 447981 321332
rect 447915 321267 447981 321268
rect 447731 319700 447797 319701
rect 447731 319636 447732 319700
rect 447796 319636 447797 319700
rect 447731 319635 447797 319636
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 159644 445574 194058
rect 448674 306334 449294 341778
rect 449574 321197 449634 700435
rect 452394 670054 453014 709082
rect 452394 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 453014 670054
rect 452394 669734 453014 669818
rect 452394 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 453014 669734
rect 452394 634054 453014 669498
rect 452394 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 453014 634054
rect 452394 633734 453014 633818
rect 452394 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 453014 633734
rect 452394 598054 453014 633498
rect 452394 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 453014 598054
rect 452394 597734 453014 597818
rect 452394 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 453014 597734
rect 452394 562054 453014 597498
rect 452394 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 453014 562054
rect 452394 561734 453014 561818
rect 452394 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 453014 561734
rect 452394 526054 453014 561498
rect 452394 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 453014 526054
rect 452394 525734 453014 525818
rect 452394 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 453014 525734
rect 452394 517884 453014 525498
rect 456114 710598 456734 711590
rect 456114 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 456734 710598
rect 456114 710278 456734 710362
rect 456114 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 456734 710278
rect 456114 673774 456734 710042
rect 456114 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 456734 673774
rect 456114 673454 456734 673538
rect 456114 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 456734 673454
rect 456114 637774 456734 673218
rect 459834 711558 460454 711590
rect 459834 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 460454 711558
rect 459834 711238 460454 711322
rect 459834 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 460454 711238
rect 459834 677494 460454 711002
rect 459834 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 460454 677494
rect 459834 677174 460454 677258
rect 459834 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 460454 677174
rect 459834 669073 460454 676938
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 669073 470414 686898
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 669073 474134 690618
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 669073 477854 694338
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 669073 481574 698058
rect 488394 709638 489014 711590
rect 488394 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 489014 709638
rect 488394 709318 489014 709402
rect 488394 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 489014 709318
rect 488394 670054 489014 709082
rect 488394 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 489014 670054
rect 488394 669734 489014 669818
rect 488394 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 489014 669734
rect 488394 669073 489014 669498
rect 492114 710598 492734 711590
rect 492114 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 492734 710598
rect 492114 710278 492734 710362
rect 492114 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 492734 710278
rect 492114 673774 492734 710042
rect 492114 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 492734 673774
rect 492114 673454 492734 673538
rect 492114 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 492734 673454
rect 492114 669073 492734 673218
rect 495834 711558 496454 711590
rect 495834 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 496454 711558
rect 495834 711238 496454 711322
rect 495834 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 496454 711238
rect 495834 677494 496454 711002
rect 495834 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 496454 677494
rect 495834 677174 496454 677258
rect 495834 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 496454 677174
rect 495834 669073 496454 676938
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 669073 506414 686898
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 669073 510134 690618
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 669073 513854 694338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 669073 517574 698058
rect 520674 708678 521294 711590
rect 520674 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 521294 708678
rect 520674 708358 521294 708442
rect 520674 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 521294 708358
rect 520674 666334 521294 708122
rect 520674 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 521294 666334
rect 520674 666014 521294 666098
rect 520674 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 521294 666014
rect 458035 665276 458101 665277
rect 458035 665212 458036 665276
rect 458100 665212 458101 665276
rect 458035 665211 458101 665212
rect 456114 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 456734 637774
rect 456114 637454 456734 637538
rect 456114 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 456734 637454
rect 456114 601774 456734 637218
rect 456114 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 456734 601774
rect 456114 601454 456734 601538
rect 456114 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 456734 601454
rect 456114 565774 456734 601218
rect 456114 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 456734 565774
rect 456114 565454 456734 565538
rect 456114 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 456734 565454
rect 456114 529774 456734 565218
rect 456114 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 456734 529774
rect 456114 529454 456734 529538
rect 456114 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 456734 529454
rect 456114 517884 456734 529218
rect 458038 517581 458098 665211
rect 459139 655756 459205 655757
rect 459139 655692 459140 655756
rect 459204 655692 459205 655756
rect 459139 655691 459205 655692
rect 458955 647732 459021 647733
rect 458955 647668 458956 647732
rect 459020 647668 459021 647732
rect 458955 647667 459021 647668
rect 458035 517580 458101 517581
rect 458035 517516 458036 517580
rect 458100 517516 458101 517580
rect 458035 517515 458101 517516
rect 451043 516764 451109 516765
rect 451043 516700 451044 516764
rect 451108 516700 451109 516764
rect 451043 516699 451109 516700
rect 450491 514384 450557 514385
rect 450491 514320 450492 514384
rect 450556 514320 450557 514384
rect 450491 514319 450557 514320
rect 450494 328677 450554 514319
rect 451046 335370 451106 516699
rect 453382 511174 453702 511206
rect 453382 510938 453424 511174
rect 453660 510938 453702 511174
rect 453382 510854 453702 510938
rect 453382 510618 453424 510854
rect 453660 510618 453702 510854
rect 453382 510586 453702 510618
rect 455820 511174 456140 511206
rect 455820 510938 455862 511174
rect 456098 510938 456140 511174
rect 455820 510854 456140 510938
rect 455820 510618 455862 510854
rect 456098 510618 456140 510854
rect 455820 510586 456140 510618
rect 458258 511174 458578 511206
rect 458258 510938 458300 511174
rect 458536 510938 458578 511174
rect 458258 510854 458578 510938
rect 458258 510618 458300 510854
rect 458536 510618 458578 510854
rect 458258 510586 458578 510618
rect 452163 507454 452483 507486
rect 452163 507218 452205 507454
rect 452441 507218 452483 507454
rect 452163 507134 452483 507218
rect 452163 506898 452205 507134
rect 452441 506898 452483 507134
rect 452163 506866 452483 506898
rect 454601 507454 454921 507486
rect 454601 507218 454643 507454
rect 454879 507218 454921 507454
rect 454601 507134 454921 507218
rect 454601 506898 454643 507134
rect 454879 506898 454921 507134
rect 454601 506866 454921 506898
rect 457039 507454 457359 507486
rect 457039 507218 457081 507454
rect 457317 507218 457359 507454
rect 457039 507134 457359 507218
rect 457039 506898 457081 507134
rect 457317 506898 457359 507134
rect 457039 506866 457359 506898
rect 450678 335310 451106 335370
rect 452394 490054 453014 500068
rect 452394 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 453014 490054
rect 452394 489734 453014 489818
rect 452394 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 453014 489734
rect 452394 454054 453014 489498
rect 452394 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 453014 454054
rect 452394 453734 453014 453818
rect 452394 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 453014 453734
rect 452394 418054 453014 453498
rect 452394 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 453014 418054
rect 452394 417734 453014 417818
rect 452394 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 453014 417734
rect 452394 382054 453014 417498
rect 452394 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 453014 382054
rect 452394 381734 453014 381818
rect 452394 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 453014 381734
rect 452394 346054 453014 381498
rect 456114 493774 456734 500068
rect 456114 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 456734 493774
rect 456114 493454 456734 493538
rect 456114 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 456734 493454
rect 456114 457774 456734 493218
rect 456114 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 456734 457774
rect 456114 457454 456734 457538
rect 456114 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 456734 457454
rect 456114 421774 456734 457218
rect 458958 428501 459018 647667
rect 459142 598229 459202 655691
rect 479568 655174 479888 655206
rect 479568 654938 479610 655174
rect 479846 654938 479888 655174
rect 479568 654854 479888 654938
rect 479568 654618 479610 654854
rect 479846 654618 479888 654854
rect 479568 654586 479888 654618
rect 510288 655174 510608 655206
rect 510288 654938 510330 655174
rect 510566 654938 510608 655174
rect 510288 654854 510608 654938
rect 510288 654618 510330 654854
rect 510566 654618 510608 654854
rect 510288 654586 510608 654618
rect 464208 651454 464528 651486
rect 464208 651218 464250 651454
rect 464486 651218 464528 651454
rect 464208 651134 464528 651218
rect 464208 650898 464250 651134
rect 464486 650898 464528 651134
rect 464208 650866 464528 650898
rect 494928 651454 495248 651486
rect 494928 651218 494970 651454
rect 495206 651218 495248 651454
rect 494928 651134 495248 651218
rect 494928 650898 494970 651134
rect 495206 650898 495248 651134
rect 494928 650866 495248 650898
rect 520674 630334 521294 665778
rect 520674 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 521294 630334
rect 520674 630014 521294 630098
rect 520674 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 521294 630014
rect 479568 619174 479888 619206
rect 479568 618938 479610 619174
rect 479846 618938 479888 619174
rect 479568 618854 479888 618938
rect 479568 618618 479610 618854
rect 479846 618618 479888 618854
rect 479568 618586 479888 618618
rect 510288 619174 510608 619206
rect 510288 618938 510330 619174
rect 510566 618938 510608 619174
rect 510288 618854 510608 618938
rect 510288 618618 510330 618854
rect 510566 618618 510608 618854
rect 510288 618586 510608 618618
rect 464208 615454 464528 615486
rect 464208 615218 464250 615454
rect 464486 615218 464528 615454
rect 464208 615134 464528 615218
rect 464208 614898 464250 615134
rect 464486 614898 464528 615134
rect 464208 614866 464528 614898
rect 494928 615454 495248 615486
rect 494928 615218 494970 615454
rect 495206 615218 495248 615454
rect 494928 615134 495248 615218
rect 494928 614898 494970 615134
rect 495206 614898 495248 615134
rect 494928 614866 495248 614898
rect 459139 598228 459205 598229
rect 459139 598164 459140 598228
rect 459204 598164 459205 598228
rect 459139 598163 459205 598164
rect 459834 569494 460454 601103
rect 459834 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 460454 569494
rect 459834 569174 460454 569258
rect 459834 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 460454 569174
rect 459834 533494 460454 568938
rect 459834 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 460454 533494
rect 459834 533174 460454 533258
rect 459834 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 460454 533174
rect 459834 517884 460454 532938
rect 469794 579454 470414 601103
rect 472019 599588 472085 599589
rect 472019 599524 472020 599588
rect 472084 599524 472085 599588
rect 472019 599523 472085 599524
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 460696 511174 461016 511206
rect 460696 510938 460738 511174
rect 460974 510938 461016 511174
rect 460696 510854 461016 510938
rect 460696 510618 460738 510854
rect 460974 510618 461016 510854
rect 460696 510586 461016 510618
rect 459477 507454 459797 507486
rect 459477 507218 459519 507454
rect 459755 507218 459797 507454
rect 459477 507134 459797 507218
rect 459477 506898 459519 507134
rect 459755 506898 459797 507134
rect 459477 506866 459797 506898
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 459834 497494 460454 500068
rect 459834 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 460454 497494
rect 459834 497174 460454 497258
rect 459834 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 460454 497174
rect 459834 461494 460454 496938
rect 459834 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 460454 461494
rect 459834 461174 460454 461258
rect 459834 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 460454 461174
rect 458955 428500 459021 428501
rect 458955 428436 458956 428500
rect 459020 428436 459021 428500
rect 458955 428435 459021 428436
rect 456114 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 456734 421774
rect 456114 421454 456734 421538
rect 456114 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 456734 421454
rect 456114 385774 456734 421218
rect 456114 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 456734 385774
rect 456114 385454 456734 385538
rect 456114 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 456734 385454
rect 454208 363454 454528 363486
rect 454208 363218 454250 363454
rect 454486 363218 454528 363454
rect 454208 363134 454528 363218
rect 454208 362898 454250 363134
rect 454486 362898 454528 363134
rect 454208 362866 454528 362898
rect 452394 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 453014 346054
rect 452394 345734 453014 345818
rect 452394 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 453014 345734
rect 450678 329221 450738 335310
rect 450675 329220 450741 329221
rect 450675 329156 450676 329220
rect 450740 329156 450741 329220
rect 450675 329155 450741 329156
rect 450491 328676 450557 328677
rect 450491 328612 450492 328676
rect 450556 328612 450557 328676
rect 450491 328611 450557 328612
rect 449571 321196 449637 321197
rect 449571 321132 449572 321196
rect 449636 321132 449637 321196
rect 449571 321131 449637 321132
rect 448674 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 449294 306334
rect 448674 306014 449294 306098
rect 448674 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 449294 306014
rect 448674 270334 449294 305778
rect 448674 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 449294 270334
rect 448674 270014 449294 270098
rect 448674 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 449294 270014
rect 448674 234334 449294 269778
rect 448674 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 449294 234334
rect 448674 234014 449294 234098
rect 448674 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 449294 234014
rect 448674 198334 449294 233778
rect 448674 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 449294 198334
rect 448674 198014 449294 198098
rect 448674 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 449294 198014
rect 448674 162334 449294 197778
rect 448674 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 449294 162334
rect 448674 162014 449294 162098
rect 448674 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 449294 162014
rect 429568 151174 429888 151206
rect 429568 150938 429610 151174
rect 429846 150938 429888 151174
rect 429568 150854 429888 150938
rect 429568 150618 429610 150854
rect 429846 150618 429888 150854
rect 429568 150586 429888 150618
rect 414208 147454 414528 147486
rect 414208 147218 414250 147454
rect 414486 147218 414528 147454
rect 414208 147134 414528 147218
rect 414208 146898 414250 147134
rect 414486 146898 414528 147134
rect 414208 146866 414528 146898
rect 444928 147454 445248 147486
rect 444928 147218 444970 147454
rect 445206 147218 445248 147454
rect 444928 147134 445248 147218
rect 444928 146898 444970 147134
rect 445206 146898 445248 147134
rect 444928 146866 445248 146898
rect 412674 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 413294 126334
rect 412674 126014 413294 126098
rect 412674 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 413294 126014
rect 412674 92137 413294 125778
rect 416394 94054 417014 127767
rect 416394 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 417014 94054
rect 416394 93734 417014 93818
rect 416394 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 417014 93734
rect 416394 92137 417014 93498
rect 420114 97774 420734 127767
rect 420114 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 420734 97774
rect 420114 97454 420734 97538
rect 420114 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 420734 97454
rect 420114 92137 420734 97218
rect 423834 101494 424454 127767
rect 423834 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 424454 101494
rect 423834 101174 424454 101258
rect 423834 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 424454 101174
rect 423834 92137 424454 100938
rect 448674 126334 449294 161778
rect 448674 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 449294 126334
rect 448674 126014 449294 126098
rect 448674 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 449294 126014
rect 448674 92137 449294 125778
rect 452394 310054 453014 345498
rect 456114 349774 456734 385218
rect 456114 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 456734 349774
rect 456114 349454 456734 349538
rect 456114 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 456734 349454
rect 454208 327454 454528 327486
rect 454208 327218 454250 327454
rect 454486 327218 454528 327454
rect 454208 327134 454528 327218
rect 454208 326898 454250 327134
rect 454486 326898 454528 327134
rect 454208 326866 454528 326898
rect 452394 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 453014 310054
rect 452394 309734 453014 309818
rect 452394 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 453014 309734
rect 452394 274054 453014 309498
rect 452394 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 453014 274054
rect 452394 273734 453014 273818
rect 452394 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 453014 273734
rect 452394 238054 453014 273498
rect 452394 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 453014 238054
rect 452394 237734 453014 237818
rect 452394 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 453014 237734
rect 452394 202054 453014 237498
rect 452394 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 453014 202054
rect 452394 201734 453014 201818
rect 452394 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 453014 201734
rect 452394 166054 453014 201498
rect 452394 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 453014 166054
rect 452394 165734 453014 165818
rect 452394 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 453014 165734
rect 452394 130054 453014 165498
rect 452394 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 453014 130054
rect 452394 129734 453014 129818
rect 452394 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 453014 129734
rect 452394 94054 453014 129498
rect 452394 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 453014 94054
rect 452394 93734 453014 93818
rect 452394 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 453014 93734
rect 452394 92137 453014 93498
rect 456114 313774 456734 349218
rect 456114 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 456734 313774
rect 456114 313454 456734 313538
rect 456114 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 456734 313454
rect 456114 277774 456734 313218
rect 456114 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 456734 277774
rect 456114 277454 456734 277538
rect 456114 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 456734 277454
rect 456114 241774 456734 277218
rect 456114 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 456734 241774
rect 456114 241454 456734 241538
rect 456114 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 456734 241454
rect 456114 205774 456734 241218
rect 456114 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 456734 205774
rect 456114 205454 456734 205538
rect 456114 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 456734 205454
rect 456114 169774 456734 205218
rect 456114 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 456734 169774
rect 456114 169454 456734 169538
rect 456114 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 456734 169454
rect 456114 133774 456734 169218
rect 456114 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 456734 133774
rect 456114 133454 456734 133538
rect 456114 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 456734 133454
rect 456114 97774 456734 133218
rect 456114 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 456734 97774
rect 456114 97454 456734 97538
rect 456114 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 456734 97454
rect 456114 92137 456734 97218
rect 459834 425494 460454 460938
rect 459834 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 460454 425494
rect 459834 425174 460454 425258
rect 459834 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 460454 425174
rect 459834 389494 460454 424938
rect 459834 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 460454 389494
rect 459834 389174 460454 389258
rect 459834 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 460454 389174
rect 459834 353494 460454 388938
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 385580 470414 398898
rect 472022 388925 472082 599523
rect 472203 589932 472269 589933
rect 472203 589868 472204 589932
rect 472268 589868 472269 589932
rect 472203 589867 472269 589868
rect 472206 389061 472266 589867
rect 473514 583174 474134 601103
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 477234 586894 477854 601103
rect 478827 598228 478893 598229
rect 478827 598164 478828 598228
rect 478892 598164 478893 598228
rect 478827 598163 478893 598164
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 474411 518124 474477 518125
rect 474411 518060 474412 518124
rect 474476 518060 474477 518124
rect 474411 518059 474477 518060
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 453692 474134 474618
rect 473416 435454 473736 435486
rect 473416 435218 473458 435454
rect 473694 435218 473736 435454
rect 473416 435134 473736 435218
rect 473416 434898 473458 435134
rect 473694 434898 473736 435134
rect 473416 434866 473736 434898
rect 474414 389061 474474 518059
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 475888 439174 476208 439206
rect 475888 438938 475930 439174
rect 476166 438938 476208 439174
rect 475888 438854 476208 438938
rect 475888 438618 475930 438854
rect 476166 438618 476208 438854
rect 475888 438586 476208 438618
rect 477234 406894 477854 442338
rect 478361 435454 478681 435486
rect 478361 435218 478403 435454
rect 478639 435218 478681 435454
rect 478361 435134 478681 435218
rect 478361 434898 478403 435134
rect 478639 434898 478681 435134
rect 478361 434866 478681 434898
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 472203 389060 472269 389061
rect 472203 388996 472204 389060
rect 472268 388996 472269 389060
rect 472203 388995 472269 388996
rect 474411 389060 474477 389061
rect 474411 388996 474412 389060
rect 474476 388996 474477 389060
rect 474411 388995 474477 388996
rect 472019 388924 472085 388925
rect 472019 388860 472020 388924
rect 472084 388860 472085 388924
rect 472019 388859 472085 388860
rect 477234 385225 477854 406338
rect 478830 389061 478890 598163
rect 480954 590614 481574 601103
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 484674 594334 485294 601103
rect 484674 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 485294 594334
rect 484674 594014 485294 594098
rect 484674 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 485294 594014
rect 484674 558334 485294 593778
rect 484674 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 485294 558334
rect 484674 558014 485294 558098
rect 484674 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 485294 558014
rect 484674 522334 485294 557778
rect 484674 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 485294 522334
rect 484674 522014 485294 522098
rect 484674 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 485294 522014
rect 484674 517884 485294 521778
rect 488394 598054 489014 601103
rect 488394 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 489014 598054
rect 488394 597734 489014 597818
rect 488394 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 489014 597734
rect 488394 562054 489014 597498
rect 488394 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 489014 562054
rect 488394 561734 489014 561818
rect 488394 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 489014 561734
rect 488394 526054 489014 561498
rect 488394 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 489014 526054
rect 488394 525734 489014 525818
rect 488394 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 489014 525734
rect 488394 517884 489014 525498
rect 492114 565774 492734 601103
rect 492114 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 492734 565774
rect 492114 565454 492734 565538
rect 492114 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 492734 565454
rect 492114 529774 492734 565218
rect 492114 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 492734 529774
rect 492114 529454 492734 529538
rect 492114 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 492734 529454
rect 482691 517580 482757 517581
rect 482691 517516 482692 517580
rect 482756 517516 482757 517580
rect 482691 517515 482757 517516
rect 482163 507454 482483 507486
rect 482163 507218 482205 507454
rect 482441 507218 482483 507454
rect 482163 507134 482483 507218
rect 482163 506898 482205 507134
rect 482441 506898 482483 507134
rect 482163 506866 482483 506898
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 453692 481574 482058
rect 482694 462909 482754 517515
rect 483382 511174 483702 511206
rect 483382 510938 483424 511174
rect 483660 510938 483702 511174
rect 483382 510854 483702 510938
rect 483382 510618 483424 510854
rect 483660 510618 483702 510854
rect 483382 510586 483702 510618
rect 485820 511174 486140 511206
rect 485820 510938 485862 511174
rect 486098 510938 486140 511174
rect 485820 510854 486140 510938
rect 485820 510618 485862 510854
rect 486098 510618 486140 510854
rect 485820 510586 486140 510618
rect 488258 511174 488578 511206
rect 488258 510938 488300 511174
rect 488536 510938 488578 511174
rect 488258 510854 488578 510938
rect 488258 510618 488300 510854
rect 488536 510618 488578 510854
rect 488258 510586 488578 510618
rect 490696 511174 491016 511206
rect 490696 510938 490738 511174
rect 490974 510938 491016 511174
rect 490696 510854 491016 510938
rect 490696 510618 490738 510854
rect 490974 510618 491016 510854
rect 490696 510586 491016 510618
rect 484601 507454 484921 507486
rect 484601 507218 484643 507454
rect 484879 507218 484921 507454
rect 484601 507134 484921 507218
rect 484601 506898 484643 507134
rect 484879 506898 484921 507134
rect 484601 506866 484921 506898
rect 487039 507454 487359 507486
rect 487039 507218 487081 507454
rect 487317 507218 487359 507454
rect 487039 507134 487359 507218
rect 487039 506898 487081 507134
rect 487317 506898 487359 507134
rect 487039 506866 487359 506898
rect 489477 507454 489797 507486
rect 489477 507218 489519 507454
rect 489755 507218 489797 507454
rect 489477 507134 489797 507218
rect 489477 506898 489519 507134
rect 489755 506898 489797 507134
rect 489477 506866 489797 506898
rect 484674 486334 485294 500068
rect 484674 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 485294 486334
rect 484674 486014 485294 486098
rect 484674 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 485294 486014
rect 482691 462908 482757 462909
rect 482691 462844 482692 462908
rect 482756 462844 482757 462908
rect 482691 462843 482757 462844
rect 484674 450334 485294 485778
rect 488394 490054 489014 500068
rect 489315 496908 489381 496909
rect 489315 496844 489316 496908
rect 489380 496844 489381 496908
rect 489315 496843 489381 496844
rect 488394 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 489014 490054
rect 488394 489734 489014 489818
rect 488394 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 489014 489734
rect 488394 454007 489014 489498
rect 488394 453771 488426 454007
rect 488662 453771 488746 454007
rect 488982 453771 489014 454007
rect 488394 453692 489014 453771
rect 484674 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 485294 450334
rect 484674 450014 485294 450098
rect 484674 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 485294 450014
rect 480833 439174 481153 439206
rect 480833 438938 480875 439174
rect 481111 438938 481153 439174
rect 480833 438854 481153 438938
rect 480833 438618 480875 438854
rect 481111 438618 481153 438854
rect 480833 438586 481153 438618
rect 483306 435454 483626 435486
rect 483306 435218 483348 435454
rect 483584 435218 483626 435454
rect 483306 435134 483626 435218
rect 483306 434898 483348 435134
rect 483584 434898 483626 435134
rect 483306 434866 483626 434898
rect 484674 414334 485294 449778
rect 485778 439174 486098 439206
rect 485778 438938 485820 439174
rect 486056 438938 486098 439174
rect 485778 438854 486098 438938
rect 485778 438618 485820 438854
rect 486056 438618 486098 438854
rect 485778 438586 486098 438618
rect 488251 435454 488571 435486
rect 488251 435218 488293 435454
rect 488529 435218 488571 435454
rect 488251 435134 488571 435218
rect 488251 434898 488293 435134
rect 488529 434898 488571 435134
rect 488251 434866 488571 434898
rect 484674 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 485294 414334
rect 484674 414014 485294 414098
rect 484674 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 485294 414014
rect 478827 389060 478893 389061
rect 478827 388996 478828 389060
rect 478892 388996 478893 389060
rect 478827 388995 478893 388996
rect 484674 385580 485294 413778
rect 489318 387021 489378 496843
rect 492114 493774 492734 529218
rect 492114 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 492734 493774
rect 492114 493454 492734 493538
rect 492114 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 492734 493454
rect 492114 457774 492734 493218
rect 492114 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 492734 457774
rect 492114 457454 492734 457538
rect 492114 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 492734 457454
rect 490723 439174 491043 439206
rect 490723 438938 490765 439174
rect 491001 438938 491043 439174
rect 490723 438854 491043 438938
rect 490723 438618 490765 438854
rect 491001 438618 491043 438854
rect 490723 438586 491043 438618
rect 492114 421774 492734 457218
rect 492114 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 492734 421774
rect 492114 421454 492734 421538
rect 492114 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 492734 421454
rect 489315 387020 489381 387021
rect 489315 386956 489316 387020
rect 489380 386956 489381 387020
rect 489315 386955 489381 386956
rect 492114 385225 492734 421218
rect 495834 569494 496454 601103
rect 495834 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 496454 569494
rect 495834 569174 496454 569258
rect 495834 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 496454 569174
rect 495834 533494 496454 568938
rect 495834 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 496454 533494
rect 495834 533174 496454 533258
rect 495834 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 496454 533174
rect 495834 497494 496454 532938
rect 495834 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 496454 497494
rect 495834 497174 496454 497258
rect 495834 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 496454 497174
rect 495834 461494 496454 496938
rect 495834 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 496454 461494
rect 495834 461174 496454 461258
rect 495834 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 496454 461174
rect 495834 425494 496454 460938
rect 495834 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 496454 425494
rect 495834 425174 496454 425258
rect 495834 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 496454 425174
rect 495834 389494 496454 424938
rect 495834 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 496454 389494
rect 495834 389174 496454 389258
rect 495834 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 496454 389174
rect 469568 367174 469888 367206
rect 469568 366938 469610 367174
rect 469846 366938 469888 367174
rect 469568 366854 469888 366938
rect 469568 366618 469610 366854
rect 469846 366618 469888 366854
rect 469568 366586 469888 366618
rect 484928 363454 485248 363486
rect 484928 363218 484970 363454
rect 485206 363218 485248 363454
rect 484928 363134 485248 363218
rect 484928 362898 484970 363134
rect 485206 362898 485248 363134
rect 484928 362866 485248 362898
rect 459834 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 460454 353494
rect 459834 353174 460454 353258
rect 459834 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 460454 353174
rect 459834 317494 460454 352938
rect 495834 353494 496454 388938
rect 505794 579454 506414 601103
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 500288 367174 500608 367206
rect 500288 366938 500330 367174
rect 500566 366938 500608 367174
rect 500288 366854 500608 366938
rect 500288 366618 500330 366854
rect 500566 366618 500608 366854
rect 500288 366586 500608 366618
rect 495834 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 496454 353494
rect 495834 353174 496454 353258
rect 495834 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 496454 353174
rect 469568 331174 469888 331206
rect 469568 330938 469610 331174
rect 469846 330938 469888 331174
rect 469568 330854 469888 330938
rect 469568 330618 469610 330854
rect 469846 330618 469888 330854
rect 469568 330586 469888 330618
rect 484928 327454 485248 327486
rect 484928 327218 484970 327454
rect 485206 327218 485248 327454
rect 484928 327134 485248 327218
rect 484928 326898 484970 327134
rect 485206 326898 485248 327134
rect 484928 326866 485248 326898
rect 459834 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 460454 317494
rect 459834 317174 460454 317258
rect 459834 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 460454 317174
rect 459834 281494 460454 316938
rect 459834 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 460454 281494
rect 459834 281174 460454 281258
rect 459834 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 460454 281174
rect 459834 245494 460454 280938
rect 477234 298894 477854 322287
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 259417 477854 262338
rect 480954 302614 481574 322287
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 259417 481574 266058
rect 484674 306334 485294 322068
rect 484674 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 485294 306334
rect 484674 306014 485294 306098
rect 484674 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 485294 306014
rect 484674 270334 485294 305778
rect 484674 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 485294 270334
rect 484674 270014 485294 270098
rect 484674 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 485294 270014
rect 484674 259417 485294 269778
rect 488394 310054 489014 322287
rect 488394 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 489014 310054
rect 488394 309734 489014 309818
rect 488394 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 489014 309734
rect 488394 274054 489014 309498
rect 488394 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 489014 274054
rect 488394 273734 489014 273818
rect 488394 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 489014 273734
rect 488394 259417 489014 273498
rect 492114 313774 492734 322287
rect 492114 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 492734 313774
rect 492114 313454 492734 313538
rect 492114 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 492734 313454
rect 492114 277774 492734 313218
rect 492114 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 492734 277774
rect 492114 277454 492734 277538
rect 492114 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 492734 277454
rect 492114 259417 492734 277218
rect 495834 317494 496454 352938
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 500288 331174 500608 331206
rect 500288 330938 500330 331174
rect 500566 330938 500608 331174
rect 500288 330854 500608 330938
rect 500288 330618 500330 330854
rect 500566 330618 500608 330854
rect 500288 330586 500608 330618
rect 495834 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 496454 317494
rect 495834 317174 496454 317258
rect 495834 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 496454 317174
rect 495834 281494 496454 316938
rect 495834 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 496454 281494
rect 495834 281174 496454 281258
rect 495834 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 496454 281174
rect 495834 259417 496454 280938
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 509514 583174 510134 601103
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 513234 586894 513854 601103
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 510659 333028 510725 333029
rect 510659 332964 510660 333028
rect 510724 332964 510725 333028
rect 510659 332963 510725 332964
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509187 322692 509253 322693
rect 509187 322628 509188 322692
rect 509252 322628 509253 322692
rect 509187 322627 509253 322628
rect 509190 321570 509250 322627
rect 509190 321510 509434 321570
rect 509374 318810 509434 321510
rect 509006 318750 509434 318810
rect 509006 306237 509066 318750
rect 509003 306236 509069 306237
rect 509003 306172 509004 306236
rect 509068 306172 509069 306236
rect 509003 306171 509069 306172
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 259417 506414 290898
rect 509514 295174 510134 330618
rect 510291 326500 510357 326501
rect 510291 326436 510292 326500
rect 510356 326436 510357 326500
rect 510291 326435 510357 326436
rect 510294 322693 510354 326435
rect 510291 322692 510357 322693
rect 510291 322628 510292 322692
rect 510356 322628 510357 322692
rect 510291 322627 510357 322628
rect 510662 297669 510722 332963
rect 510843 325956 510909 325957
rect 510843 325892 510844 325956
rect 510908 325892 510909 325956
rect 510843 325891 510909 325892
rect 510846 322285 510906 325891
rect 511211 324324 511277 324325
rect 511211 324260 511212 324324
rect 511276 324260 511277 324324
rect 511211 324259 511277 324260
rect 511027 323780 511093 323781
rect 511027 323716 511028 323780
rect 511092 323716 511093 323780
rect 511027 323715 511093 323716
rect 510843 322284 510909 322285
rect 510843 322220 510844 322284
rect 510908 322220 510909 322284
rect 510843 322219 510909 322220
rect 511030 322010 511090 323715
rect 510846 321950 511090 322010
rect 510846 305965 510906 321950
rect 511214 321570 511274 324259
rect 511030 321510 511274 321570
rect 510843 305964 510909 305965
rect 510843 305900 510844 305964
rect 510908 305900 510909 305964
rect 510843 305899 510909 305900
rect 511030 305829 511090 321510
rect 511027 305828 511093 305829
rect 511027 305764 511028 305828
rect 511092 305764 511093 305828
rect 511027 305763 511093 305764
rect 513234 298894 513854 334338
rect 516954 590614 517574 601103
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 515075 330308 515141 330309
rect 515075 330244 515076 330308
rect 515140 330244 515141 330308
rect 515075 330243 515141 330244
rect 514891 329764 514957 329765
rect 514891 329700 514892 329764
rect 514956 329700 514957 329764
rect 514891 329699 514957 329700
rect 514155 328676 514221 328677
rect 514155 328612 514156 328676
rect 514220 328612 514221 328676
rect 514155 328611 514221 328612
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 510659 297668 510725 297669
rect 510659 297604 510660 297668
rect 510724 297604 510725 297668
rect 510659 297603 510725 297604
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259417 510134 294618
rect 513234 262894 513854 298338
rect 514158 294541 514218 328611
rect 514894 297533 514954 329699
rect 514891 297532 514957 297533
rect 514891 297468 514892 297532
rect 514956 297468 514957 297532
rect 514891 297467 514957 297468
rect 514155 294540 514221 294541
rect 514155 294476 514156 294540
rect 514220 294476 514221 294540
rect 514155 294475 514221 294476
rect 515078 291821 515138 330243
rect 516954 302614 517574 338058
rect 520674 594334 521294 629778
rect 520674 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 521294 594334
rect 520674 594014 521294 594098
rect 520674 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 521294 594014
rect 520674 558334 521294 593778
rect 520674 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 521294 558334
rect 520674 558014 521294 558098
rect 520674 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 521294 558014
rect 520674 522334 521294 557778
rect 520674 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 521294 522334
rect 520674 522014 521294 522098
rect 520674 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 521294 522014
rect 520674 486334 521294 521778
rect 520674 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 521294 486334
rect 520674 486014 521294 486098
rect 520674 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 521294 486014
rect 520674 450334 521294 485778
rect 520674 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 521294 450334
rect 520674 450014 521294 450098
rect 520674 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 521294 450014
rect 520674 414334 521294 449778
rect 520674 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 521294 414334
rect 520674 414014 521294 414098
rect 520674 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 521294 414014
rect 520674 378334 521294 413778
rect 520674 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 521294 378334
rect 520674 378014 521294 378098
rect 520674 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 521294 378014
rect 520674 342334 521294 377778
rect 520674 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 521294 342334
rect 520674 342014 521294 342098
rect 520674 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 521294 342014
rect 518019 332484 518085 332485
rect 518019 332420 518020 332484
rect 518084 332420 518085 332484
rect 518019 332419 518085 332420
rect 517835 324868 517901 324869
rect 517835 324804 517836 324868
rect 517900 324804 517901 324868
rect 517835 324803 517901 324804
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 515075 291820 515141 291821
rect 515075 291756 515076 291820
rect 515140 291756 515141 291820
rect 515075 291755 515141 291756
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 259417 513854 262338
rect 516954 266614 517574 302058
rect 517838 297397 517898 324803
rect 518022 306917 518082 332419
rect 518019 306916 518085 306917
rect 518019 306852 518020 306916
rect 518084 306852 518085 306916
rect 518019 306851 518085 306852
rect 520674 306334 521294 341778
rect 520674 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 521294 306334
rect 520674 306014 521294 306098
rect 520674 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 521294 306014
rect 517835 297396 517901 297397
rect 517835 297332 517836 297396
rect 517900 297332 517901 297396
rect 517835 297331 517901 297332
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 259417 517574 266058
rect 520674 270334 521294 305778
rect 520674 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 521294 270334
rect 520674 270014 521294 270098
rect 520674 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 521294 270014
rect 520674 259417 521294 269778
rect 524394 709638 525014 711590
rect 524394 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 525014 709638
rect 524394 709318 525014 709402
rect 524394 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 525014 709318
rect 524394 670054 525014 709082
rect 528114 710598 528734 711590
rect 528114 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 528734 710598
rect 528114 710278 528734 710362
rect 528114 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 528734 710278
rect 526299 699820 526365 699821
rect 526299 699756 526300 699820
rect 526364 699756 526365 699820
rect 526299 699755 526365 699756
rect 524394 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 525014 670054
rect 524394 669734 525014 669818
rect 524394 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 525014 669734
rect 524394 634054 525014 669498
rect 525648 651454 525968 651486
rect 525648 651218 525690 651454
rect 525926 651218 525968 651454
rect 525648 651134 525968 651218
rect 525648 650898 525690 651134
rect 525926 650898 525968 651134
rect 525648 650866 525968 650898
rect 524394 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 525014 634054
rect 524394 633734 525014 633818
rect 524394 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 525014 633734
rect 524394 598054 525014 633498
rect 525648 615454 525968 615486
rect 525648 615218 525690 615454
rect 525926 615218 525968 615454
rect 525648 615134 525968 615218
rect 525648 614898 525690 615134
rect 525926 614898 525968 615134
rect 525648 614866 525968 614898
rect 524394 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 525014 598054
rect 524394 597734 525014 597818
rect 524394 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 525014 597734
rect 524394 562054 525014 597498
rect 524394 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 525014 562054
rect 524394 561734 525014 561818
rect 524394 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 525014 561734
rect 524394 526054 525014 561498
rect 524394 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 525014 526054
rect 524394 525734 525014 525818
rect 524394 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 525014 525734
rect 524394 490054 525014 525498
rect 524394 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 525014 490054
rect 524394 489734 525014 489818
rect 524394 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 525014 489734
rect 524394 454054 525014 489498
rect 524394 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 525014 454054
rect 524394 453734 525014 453818
rect 524394 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 525014 453734
rect 524394 418054 525014 453498
rect 525164 435454 525484 435486
rect 525164 435218 525206 435454
rect 525442 435218 525484 435454
rect 525164 435134 525484 435218
rect 525164 434898 525206 435134
rect 525442 434898 525484 435134
rect 525164 434866 525484 434898
rect 524394 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 525014 418054
rect 524394 417734 525014 417818
rect 524394 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 525014 417734
rect 524394 382054 525014 417498
rect 524394 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 525014 382054
rect 524394 381734 525014 381818
rect 524394 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 525014 381734
rect 524394 346054 525014 381498
rect 524394 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 525014 346054
rect 524394 345734 525014 345818
rect 524394 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 525014 345734
rect 524394 310054 525014 345498
rect 526302 322829 526362 699755
rect 528114 673774 528734 710042
rect 531834 711558 532454 711590
rect 531834 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 532454 711558
rect 531834 711238 532454 711322
rect 531834 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 532454 711238
rect 530531 700364 530597 700365
rect 530531 700300 530532 700364
rect 530596 700300 530597 700364
rect 530531 700299 530597 700300
rect 528114 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 528734 673774
rect 528114 673454 528734 673538
rect 528114 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 528734 673454
rect 528114 637774 528734 673218
rect 528114 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 528734 637774
rect 528114 637454 528734 637538
rect 528114 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 528734 637454
rect 528114 601774 528734 637218
rect 528114 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 528734 601774
rect 528114 601454 528734 601538
rect 528114 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 528734 601454
rect 528114 565774 528734 601218
rect 528114 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 528734 565774
rect 528114 565454 528734 565538
rect 528114 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 528734 565454
rect 528114 529774 528734 565218
rect 528114 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 528734 529774
rect 528114 529454 528734 529538
rect 528114 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 528734 529454
rect 528114 493774 528734 529218
rect 528114 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 528734 493774
rect 528114 493454 528734 493538
rect 528114 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 528734 493454
rect 528114 457774 528734 493218
rect 528114 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 528734 457774
rect 528114 457454 528734 457538
rect 528114 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 528734 457454
rect 528114 421774 528734 457218
rect 529384 439174 529704 439206
rect 529384 438938 529426 439174
rect 529662 438938 529704 439174
rect 529384 438854 529704 438938
rect 529384 438618 529426 438854
rect 529662 438618 529704 438854
rect 529384 438586 529704 438618
rect 528114 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 528734 421774
rect 528114 421454 528734 421538
rect 528114 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 528734 421454
rect 528114 385774 528734 421218
rect 528114 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 528734 385774
rect 528114 385454 528734 385538
rect 528114 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 528734 385454
rect 528114 349774 528734 385218
rect 528114 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 528734 349774
rect 528114 349454 528734 349538
rect 528114 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 528734 349454
rect 526299 322828 526365 322829
rect 526299 322764 526300 322828
rect 526364 322764 526365 322828
rect 526299 322763 526365 322764
rect 524394 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 525014 310054
rect 524394 309734 525014 309818
rect 524394 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 525014 309734
rect 524394 274054 525014 309498
rect 524394 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 525014 274054
rect 524394 273734 525014 273818
rect 524394 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 525014 273734
rect 524394 259417 525014 273498
rect 528114 313774 528734 349218
rect 530534 321333 530594 700299
rect 531834 677494 532454 711002
rect 531834 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 532454 677494
rect 531834 677174 532454 677258
rect 531834 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 532454 677174
rect 531834 641494 532454 676938
rect 531834 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 532454 641494
rect 531834 641174 532454 641258
rect 531834 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 532454 641174
rect 531834 605494 532454 640938
rect 531834 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 532454 605494
rect 531834 605174 532454 605258
rect 531834 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 532454 605174
rect 531834 569494 532454 604938
rect 531834 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 532454 569494
rect 531834 569174 532454 569258
rect 531834 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 532454 569174
rect 531834 533494 532454 568938
rect 531834 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 532454 533494
rect 531834 533174 532454 533258
rect 531834 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 532454 533174
rect 531834 497494 532454 532938
rect 531834 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 532454 497494
rect 531834 497174 532454 497258
rect 531834 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 532454 497174
rect 531834 461494 532454 496938
rect 531834 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 532454 461494
rect 531834 461174 532454 461258
rect 531834 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 532454 461174
rect 531834 425494 532454 460938
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 460836 542414 470898
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 537825 439174 538145 439206
rect 537825 438938 537867 439174
rect 538103 438938 538145 439174
rect 537825 438854 538145 438938
rect 537825 438618 537867 438854
rect 538103 438618 538145 438854
rect 537825 438586 538145 438618
rect 545514 439174 546134 474618
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 533605 435454 533925 435486
rect 533605 435218 533647 435454
rect 533883 435218 533925 435454
rect 533605 435134 533925 435218
rect 533605 434898 533647 435134
rect 533883 434898 533925 435134
rect 533605 434866 533925 434898
rect 542046 435454 542366 435486
rect 542046 435218 542088 435454
rect 542324 435218 542366 435454
rect 542046 435134 542366 435218
rect 542046 434898 542088 435134
rect 542324 434898 542366 435134
rect 542046 434866 542366 434898
rect 531834 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 532454 425494
rect 531834 425174 532454 425258
rect 531834 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 532454 425174
rect 531834 389494 532454 424938
rect 531834 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 532454 389494
rect 531834 389174 532454 389258
rect 531834 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 532454 389174
rect 531834 353494 532454 388938
rect 531834 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 532454 353494
rect 531834 353174 532454 353258
rect 531834 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 532454 353174
rect 530531 321332 530597 321333
rect 530531 321268 530532 321332
rect 530596 321268 530597 321332
rect 530531 321267 530597 321268
rect 528114 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 528734 313774
rect 528114 313454 528734 313538
rect 528114 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 528734 313454
rect 528114 277774 528734 313218
rect 528114 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 528734 277774
rect 528114 277454 528734 277538
rect 528114 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 528734 277454
rect 528114 259417 528734 277218
rect 531834 317494 532454 352938
rect 541794 399454 542414 425068
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 538811 319564 538877 319565
rect 538811 319500 538812 319564
rect 538876 319500 538877 319564
rect 538811 319499 538877 319500
rect 531834 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 532454 317494
rect 531834 317174 532454 317258
rect 531834 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 532454 317174
rect 531834 281494 532454 316938
rect 538259 313988 538325 313989
rect 538259 313924 538260 313988
rect 538324 313924 538325 313988
rect 538259 313923 538325 313924
rect 531834 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 532454 281494
rect 531834 281174 532454 281258
rect 531834 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 532454 281174
rect 479568 259174 479888 259206
rect 479568 258938 479610 259174
rect 479846 258938 479888 259174
rect 479568 258854 479888 258938
rect 479568 258618 479610 258854
rect 479846 258618 479888 258854
rect 479568 258586 479888 258618
rect 510288 259174 510608 259206
rect 510288 258938 510330 259174
rect 510566 258938 510608 259174
rect 510288 258854 510608 258938
rect 510288 258618 510330 258854
rect 510566 258618 510608 258854
rect 510288 258586 510608 258618
rect 464208 255454 464528 255486
rect 464208 255218 464250 255454
rect 464486 255218 464528 255454
rect 464208 255134 464528 255218
rect 464208 254898 464250 255134
rect 464486 254898 464528 255134
rect 464208 254866 464528 254898
rect 494928 255454 495248 255486
rect 494928 255218 494970 255454
rect 495206 255218 495248 255454
rect 494928 255134 495248 255218
rect 494928 254898 494970 255134
rect 495206 254898 495248 255134
rect 494928 254866 495248 254898
rect 525648 255454 525968 255486
rect 525648 255218 525690 255454
rect 525926 255218 525968 255454
rect 525648 255134 525968 255218
rect 525648 254898 525690 255134
rect 525926 254898 525968 255134
rect 525648 254866 525968 254898
rect 459834 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 460454 245494
rect 459834 245174 460454 245258
rect 459834 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 460454 245174
rect 459834 209494 460454 244938
rect 531834 245494 532454 280938
rect 531834 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 532454 245494
rect 531834 245174 532454 245258
rect 531834 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 532454 245174
rect 479568 223174 479888 223206
rect 479568 222938 479610 223174
rect 479846 222938 479888 223174
rect 479568 222854 479888 222938
rect 479568 222618 479610 222854
rect 479846 222618 479888 222854
rect 479568 222586 479888 222618
rect 510288 223174 510608 223206
rect 510288 222938 510330 223174
rect 510566 222938 510608 223174
rect 510288 222854 510608 222938
rect 510288 222618 510330 222854
rect 510566 222618 510608 222854
rect 510288 222586 510608 222618
rect 464208 219454 464528 219486
rect 464208 219218 464250 219454
rect 464486 219218 464528 219454
rect 464208 219134 464528 219218
rect 464208 218898 464250 219134
rect 464486 218898 464528 219134
rect 464208 218866 464528 218898
rect 494928 219454 495248 219486
rect 494928 219218 494970 219454
rect 495206 219218 495248 219454
rect 494928 219134 495248 219218
rect 494928 218898 494970 219134
rect 495206 218898 495248 219134
rect 494928 218866 495248 218898
rect 525648 219454 525968 219486
rect 525648 219218 525690 219454
rect 525926 219218 525968 219454
rect 525648 219134 525968 219218
rect 525648 218898 525690 219134
rect 525926 218898 525968 219134
rect 525648 218866 525968 218898
rect 459834 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 460454 209494
rect 459834 209174 460454 209258
rect 459834 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 460454 209174
rect 459834 173494 460454 208938
rect 531834 209494 532454 244938
rect 531834 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 532454 209494
rect 531834 209174 532454 209258
rect 531834 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 532454 209174
rect 459834 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 460454 173494
rect 459834 173174 460454 173258
rect 459834 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 460454 173174
rect 459834 137494 460454 172938
rect 459834 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 460454 137494
rect 459834 137174 460454 137258
rect 459834 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 460454 137174
rect 459834 101494 460454 136938
rect 459834 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 460454 101494
rect 459834 101174 460454 101258
rect 459834 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 460454 101174
rect 405568 79174 405888 79206
rect 405568 78938 405610 79174
rect 405846 78938 405888 79174
rect 405568 78854 405888 78938
rect 405568 78618 405610 78854
rect 405846 78618 405888 78854
rect 405568 78586 405888 78618
rect 436288 79174 436608 79206
rect 436288 78938 436330 79174
rect 436566 78938 436608 79174
rect 436288 78854 436608 78938
rect 436288 78618 436330 78854
rect 436566 78618 436608 78854
rect 436288 78586 436608 78618
rect 390208 75454 390528 75486
rect 390208 75218 390250 75454
rect 390486 75218 390528 75454
rect 390208 75134 390528 75218
rect 390208 74898 390250 75134
rect 390486 74898 390528 75134
rect 390208 74866 390528 74898
rect 420928 75454 421248 75486
rect 420928 75218 420970 75454
rect 421206 75218 421248 75454
rect 420928 75134 421248 75218
rect 420928 74898 420970 75134
rect 421206 74898 421248 75134
rect 420928 74866 421248 74898
rect 451648 75454 451968 75486
rect 451648 75218 451690 75454
rect 451926 75218 451968 75454
rect 451648 75134 451968 75218
rect 451648 74898 451690 75134
rect 451926 74898 451968 75134
rect 451648 74866 451968 74898
rect 384114 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 384734 61774
rect 384114 61454 384734 61538
rect 384114 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 384734 61454
rect 384114 25774 384734 61218
rect 459834 65494 460454 100938
rect 459834 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 460454 65494
rect 459834 65174 460454 65258
rect 459834 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 460454 65174
rect 405568 43174 405888 43206
rect 405568 42938 405610 43174
rect 405846 42938 405888 43174
rect 405568 42854 405888 42938
rect 405568 42618 405610 42854
rect 405846 42618 405888 42854
rect 405568 42586 405888 42618
rect 436288 43174 436608 43206
rect 436288 42938 436330 43174
rect 436566 42938 436608 43174
rect 436288 42854 436608 42938
rect 436288 42618 436330 42854
rect 436566 42618 436608 42854
rect 436288 42586 436608 42618
rect 390208 39454 390528 39486
rect 390208 39218 390250 39454
rect 390486 39218 390528 39454
rect 390208 39134 390528 39218
rect 390208 38898 390250 39134
rect 390486 38898 390528 39134
rect 390208 38866 390528 38898
rect 420928 39454 421248 39486
rect 420928 39218 420970 39454
rect 421206 39218 421248 39454
rect 420928 39134 421248 39218
rect 420928 38898 420970 39134
rect 421206 38898 421248 39134
rect 420928 38866 421248 38898
rect 451648 39454 451968 39486
rect 451648 39218 451690 39454
rect 451926 39218 451968 39454
rect 451648 39134 451968 39218
rect 451648 38898 451690 39134
rect 451926 38898 451968 39134
rect 451648 38866 451968 38898
rect 384114 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 384734 25774
rect 384114 25454 384734 25538
rect 384114 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 384734 25454
rect 384114 -6106 384734 25218
rect 384114 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 384734 -6106
rect 384114 -6426 384734 -6342
rect 384114 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 384734 -6426
rect 384114 -7654 384734 -6662
rect 387834 29494 388454 31919
rect 387834 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 388454 29494
rect 387834 29174 388454 29258
rect 387834 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 388454 29174
rect 387834 -7066 388454 28938
rect 387834 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 388454 -7066
rect 387834 -7386 388454 -7302
rect 387834 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 388454 -7386
rect 387834 -7654 388454 -7622
rect 397794 3454 398414 31919
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 7174 402134 31919
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 10894 405854 30068
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 408954 14614 409574 31919
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 408954 -3226 409574 14058
rect 408954 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 409574 -3226
rect 408954 -3546 409574 -3462
rect 408954 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 409574 -3546
rect 408954 -7654 409574 -3782
rect 412674 18334 413294 31919
rect 412674 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 413294 18334
rect 412674 18014 413294 18098
rect 412674 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 413294 18014
rect 412674 -4186 413294 17778
rect 412674 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 413294 -4186
rect 412674 -4506 413294 -4422
rect 412674 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 413294 -4506
rect 412674 -7654 413294 -4742
rect 416394 22054 417014 31919
rect 416394 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 417014 22054
rect 416394 21734 417014 21818
rect 416394 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 417014 21734
rect 416394 -5146 417014 21498
rect 416394 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 417014 -5146
rect 416394 -5466 417014 -5382
rect 416394 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 417014 -5466
rect 416394 -7654 417014 -5702
rect 420114 25774 420734 31919
rect 420114 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 420734 25774
rect 420114 25454 420734 25538
rect 420114 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 420734 25454
rect 420114 -6106 420734 25218
rect 420114 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 420734 -6106
rect 420114 -6426 420734 -6342
rect 420114 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 420734 -6426
rect 420114 -7654 420734 -6662
rect 423834 29494 424454 31919
rect 423834 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 424454 29494
rect 423834 29174 424454 29258
rect 423834 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 424454 29174
rect 423834 -7066 424454 28938
rect 423834 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 424454 -7066
rect 423834 -7386 424454 -7302
rect 423834 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 424454 -7386
rect 423834 -7654 424454 -7622
rect 433794 3454 434414 31919
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 7174 438134 31919
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 10894 441854 31919
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 444954 14614 445574 31919
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 444954 -3226 445574 14058
rect 444954 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 445574 -3226
rect 444954 -3546 445574 -3462
rect 444954 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 445574 -3546
rect 444954 -7654 445574 -3782
rect 448674 18334 449294 31919
rect 448674 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 449294 18334
rect 448674 18014 449294 18098
rect 448674 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 449294 18014
rect 448674 -4186 449294 17778
rect 448674 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 449294 -4186
rect 448674 -4506 449294 -4422
rect 448674 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 449294 -4506
rect 448674 -7654 449294 -4742
rect 452394 22054 453014 31919
rect 452394 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 453014 22054
rect 452394 21734 453014 21818
rect 452394 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 453014 21734
rect 452394 -5146 453014 21498
rect 452394 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 453014 -5146
rect 452394 -5466 453014 -5382
rect 452394 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 453014 -5466
rect 452394 -7654 453014 -5702
rect 456114 25774 456734 31919
rect 456114 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 456734 25774
rect 456114 25454 456734 25538
rect 456114 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 456734 25454
rect 456114 -6106 456734 25218
rect 456114 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 456734 -6106
rect 456114 -6426 456734 -6342
rect 456114 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 456734 -6426
rect 456114 -7654 456734 -6662
rect 459834 29494 460454 64938
rect 459834 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 460454 29494
rect 459834 29174 460454 29258
rect 459834 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 460454 29174
rect 459834 -7066 460454 28938
rect 459834 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 460454 -7066
rect 459834 -7386 460454 -7302
rect 459834 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 460454 -7386
rect 459834 -7654 460454 -7622
rect 469794 183454 470414 201919
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 187174 474134 201919
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 190894 477854 201919
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 480954 194614 481574 201919
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 484674 198334 485294 201919
rect 484674 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 485294 198334
rect 484674 198014 485294 198098
rect 484674 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 485294 198014
rect 484674 162334 485294 197778
rect 484674 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 485294 162334
rect 484674 162014 485294 162098
rect 484674 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 485294 162014
rect 484674 126334 485294 161778
rect 488394 166054 489014 201919
rect 488394 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 489014 166054
rect 488394 165734 489014 165818
rect 488394 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 489014 165734
rect 488394 139281 489014 165498
rect 505794 183454 506414 201919
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 139281 506414 146898
rect 509514 187174 510134 201919
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 139281 510134 150618
rect 513234 190894 513854 201919
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 139281 513854 154338
rect 516954 194614 517574 201919
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 139281 517574 158058
rect 520674 198334 521294 201919
rect 520674 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 521294 198334
rect 520674 198014 521294 198098
rect 520674 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 521294 198014
rect 520674 162334 521294 197778
rect 520674 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 521294 162334
rect 520674 162014 521294 162098
rect 520674 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 521294 162014
rect 520674 139281 521294 161778
rect 524394 166054 525014 201919
rect 524394 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 525014 166054
rect 524394 165734 525014 165818
rect 524394 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 525014 165734
rect 524394 139281 525014 165498
rect 531834 173494 532454 208938
rect 531834 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 532454 173494
rect 531834 173174 532454 173258
rect 531834 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 532454 173174
rect 531834 139281 532454 172938
rect 538262 137730 538322 313923
rect 538814 137869 538874 319499
rect 541794 291454 542414 326898
rect 545514 403174 546134 438618
rect 546266 439174 546586 439206
rect 546266 438938 546308 439174
rect 546544 438938 546586 439174
rect 546266 438854 546586 438938
rect 546266 438618 546308 438854
rect 546544 438618 546586 438854
rect 546266 438586 546586 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 542675 318068 542741 318069
rect 542675 318004 542676 318068
rect 542740 318004 542741 318068
rect 542675 318003 542741 318004
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 538811 137868 538877 137869
rect 538811 137804 538812 137868
rect 538876 137804 538877 137868
rect 538811 137803 538877 137804
rect 538262 137670 539426 137730
rect 539366 133381 539426 137670
rect 539363 133380 539429 133381
rect 539363 133316 539364 133380
rect 539428 133316 539429 133380
rect 539363 133315 539429 133316
rect 484674 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 485294 126334
rect 484674 126014 485294 126098
rect 484674 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 485294 126014
rect 484208 111454 484528 111486
rect 484208 111218 484250 111454
rect 484486 111218 484528 111454
rect 484208 111134 484528 111218
rect 484208 110898 484250 111134
rect 484486 110898 484528 111134
rect 484208 110866 484528 110898
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 480954 -3226 481574 14058
rect 480954 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 481574 -3226
rect 480954 -3546 481574 -3462
rect 480954 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 481574 -3546
rect 480954 -7654 481574 -3782
rect 484674 90334 485294 125778
rect 499568 115174 499888 115206
rect 499568 114938 499610 115174
rect 499846 114938 499888 115174
rect 499568 114854 499888 114938
rect 499568 114618 499610 114854
rect 499846 114618 499888 114854
rect 499568 114586 499888 114618
rect 530288 115174 530608 115206
rect 530288 114938 530330 115174
rect 530566 114938 530608 115174
rect 530288 114854 530608 114938
rect 530288 114618 530330 114854
rect 530566 114618 530608 114854
rect 530288 114586 530608 114618
rect 514928 111454 515248 111486
rect 514928 111218 514970 111454
rect 515206 111218 515248 111454
rect 514928 111134 515248 111218
rect 514928 110898 514970 111134
rect 515206 110898 515248 111134
rect 514928 110866 515248 110898
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 484674 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 485294 90334
rect 484674 90014 485294 90098
rect 484674 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 485294 90014
rect 484674 54334 485294 89778
rect 484674 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 485294 54334
rect 484674 54014 485294 54098
rect 484674 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 485294 54014
rect 484674 18334 485294 53778
rect 484674 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 485294 18334
rect 484674 18014 485294 18098
rect 484674 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 485294 18014
rect 484674 -4186 485294 17778
rect 484674 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 485294 -4186
rect 484674 -4506 485294 -4422
rect 484674 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 485294 -4506
rect 484674 -7654 485294 -4742
rect 488394 58054 489014 82599
rect 488394 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 489014 58054
rect 488394 57734 489014 57818
rect 488394 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 489014 57734
rect 488394 22054 489014 57498
rect 488394 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 489014 22054
rect 488394 21734 489014 21818
rect 488394 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 489014 21734
rect 488394 -5146 489014 21498
rect 488394 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 489014 -5146
rect 488394 -5466 489014 -5382
rect 488394 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 489014 -5466
rect 488394 -7654 489014 -5702
rect 492114 61774 492734 82599
rect 492114 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 492734 61774
rect 492114 61454 492734 61538
rect 492114 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 492734 61454
rect 492114 25774 492734 61218
rect 492114 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 492734 25774
rect 492114 25454 492734 25538
rect 492114 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 492734 25454
rect 492114 -6106 492734 25218
rect 492114 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 492734 -6106
rect 492114 -6426 492734 -6342
rect 492114 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 492734 -6426
rect 492114 -7654 492734 -6662
rect 495834 65494 496454 82599
rect 495834 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 496454 65494
rect 495834 65174 496454 65258
rect 495834 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 496454 65174
rect 495834 29494 496454 64938
rect 495834 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 496454 29494
rect 495834 29174 496454 29258
rect 495834 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 496454 29174
rect 495834 -7066 496454 28938
rect 495834 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 496454 -7066
rect 495834 -7386 496454 -7302
rect 495834 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 496454 -7386
rect 495834 -7654 496454 -7622
rect 505794 75454 506414 82599
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 79174 510134 82599
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 46894 513854 82599
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 516954 50614 517574 82599
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 516954 -3226 517574 14058
rect 516954 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 517574 -3226
rect 516954 -3546 517574 -3462
rect 516954 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 517574 -3546
rect 516954 -7654 517574 -3782
rect 520674 54334 521294 82599
rect 520674 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 521294 54334
rect 520674 54014 521294 54098
rect 520674 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 521294 54014
rect 520674 18334 521294 53778
rect 520674 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 521294 18334
rect 520674 18014 521294 18098
rect 520674 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 521294 18014
rect 520674 -4186 521294 17778
rect 520674 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 521294 -4186
rect 520674 -4506 521294 -4422
rect 520674 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 521294 -4506
rect 520674 -7654 521294 -4742
rect 524394 58054 525014 82599
rect 524394 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 525014 58054
rect 524394 57734 525014 57818
rect 524394 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 525014 57734
rect 524394 22054 525014 57498
rect 524394 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 525014 22054
rect 524394 21734 525014 21818
rect 524394 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 525014 21734
rect 524394 -5146 525014 21498
rect 524394 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 525014 -5146
rect 524394 -5466 525014 -5382
rect 524394 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 525014 -5466
rect 524394 -7654 525014 -5702
rect 528114 61774 528734 82599
rect 528114 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 528734 61774
rect 528114 61454 528734 61538
rect 528114 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 528734 61454
rect 528114 25774 528734 61218
rect 528114 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 528734 25774
rect 528114 25454 528734 25538
rect 528114 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 528734 25454
rect 528114 -6106 528734 25218
rect 528114 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 528734 -6106
rect 528114 -6426 528734 -6342
rect 528114 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 528734 -6426
rect 528114 -7654 528734 -6662
rect 531834 65494 532454 82599
rect 531834 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 532454 65494
rect 531834 65174 532454 65258
rect 531834 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 532454 65174
rect 531834 29494 532454 64938
rect 531834 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 532454 29494
rect 531834 29174 532454 29258
rect 531834 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 532454 29174
rect 531834 -7066 532454 28938
rect 531834 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 532454 -7066
rect 531834 -7386 532454 -7302
rect 531834 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 532454 -7386
rect 531834 -7654 532454 -7622
rect 541794 75454 542414 110898
rect 542678 84421 542738 318003
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 542675 84420 542741 84421
rect 542675 84356 542676 84420
rect 542740 84356 542741 84420
rect 542675 84355 542741 84356
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 51692 546134 78618
rect 549234 406894 549854 442338
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 550487 435454 550807 435486
rect 550487 435218 550529 435454
rect 550765 435218 550807 435454
rect 550487 435134 550807 435218
rect 550487 434898 550529 435134
rect 550765 434898 550807 435134
rect 550487 434866 550807 434898
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 552954 410614 553574 446058
rect 556674 708678 557294 711590
rect 556674 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 557294 708678
rect 556674 708358 557294 708442
rect 556674 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 557294 708358
rect 556674 666334 557294 708122
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 558131 699820 558197 699821
rect 558131 699756 558132 699820
rect 558196 699756 558197 699820
rect 558131 699755 558197 699756
rect 556674 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 557294 666334
rect 556674 666014 557294 666098
rect 556674 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 557294 666014
rect 556674 630334 557294 665778
rect 556674 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 557294 630334
rect 556674 630014 557294 630098
rect 556674 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 557294 630014
rect 556674 594334 557294 629778
rect 556674 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 557294 594334
rect 556674 594014 557294 594098
rect 556674 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 557294 594014
rect 556674 558334 557294 593778
rect 556674 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 557294 558334
rect 556674 558014 557294 558098
rect 556674 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 557294 558014
rect 556674 522334 557294 557778
rect 556674 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 557294 522334
rect 556674 522014 557294 522098
rect 556674 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 557294 522014
rect 556674 486334 557294 521778
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 554707 439174 555027 439206
rect 554707 438938 554749 439174
rect 554985 438938 555027 439174
rect 554707 438854 555027 438938
rect 554707 438618 554749 438854
rect 554985 438618 555027 438854
rect 554707 438586 555027 438618
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 377884 553574 410058
rect 556674 414334 557294 449778
rect 556674 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 557294 414334
rect 556674 414014 557294 414098
rect 556674 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 557294 414014
rect 556674 378243 557294 413778
rect 556674 378007 556706 378243
rect 556942 378007 557026 378243
rect 557262 378007 557294 378243
rect 556674 377884 557294 378007
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 554876 367174 555196 367206
rect 554876 366938 554918 367174
rect 555154 366938 555196 367174
rect 554876 366854 555196 366938
rect 554876 366618 554918 366854
rect 555154 366618 555196 366854
rect 554876 366586 555196 366618
rect 552910 363454 553230 363486
rect 552910 363218 552952 363454
rect 553188 363218 553230 363454
rect 552910 363134 553230 363218
rect 552910 362898 552952 363134
rect 553188 362898 553230 363134
rect 552910 362866 553230 362898
rect 556843 363454 557163 363486
rect 556843 363218 556885 363454
rect 557121 363218 557163 363454
rect 556843 363134 557163 363218
rect 556843 362898 556885 363134
rect 557121 362898 557163 363134
rect 556843 362866 557163 362898
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 552954 338614 553574 360068
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 51692 553574 86058
rect 556674 342334 557294 360068
rect 556674 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 557294 342334
rect 556674 342014 557294 342098
rect 556674 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 557294 342014
rect 556674 306334 557294 341778
rect 558134 321469 558194 699755
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 560394 377884 561014 381498
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 377884 564734 385218
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 558809 367174 559129 367206
rect 558809 366938 558851 367174
rect 559087 366938 559129 367174
rect 558809 366854 559129 366938
rect 558809 366618 558851 366854
rect 559087 366618 559129 366854
rect 558809 366586 559129 366618
rect 562742 367174 563062 367206
rect 562742 366938 562784 367174
rect 563020 366938 563062 367174
rect 562742 366854 563062 366938
rect 562742 366618 562784 366854
rect 563020 366618 563062 366854
rect 562742 366586 563062 366618
rect 566675 367174 566995 367206
rect 566675 366938 566717 367174
rect 566953 366938 566995 367174
rect 566675 366854 566995 366938
rect 566675 366618 566717 366854
rect 566953 366618 566995 366854
rect 566675 366586 566995 366618
rect 560776 363454 561096 363486
rect 560776 363218 560818 363454
rect 561054 363218 561096 363454
rect 560776 363134 561096 363218
rect 560776 362898 560818 363134
rect 561054 362898 561096 363134
rect 560776 362866 561096 362898
rect 564709 363454 565029 363486
rect 564709 363218 564751 363454
rect 564987 363218 565029 363454
rect 564709 363134 565029 363218
rect 564709 362898 564751 363134
rect 564987 362898 565029 363134
rect 564709 362866 565029 362898
rect 560394 346054 561014 360068
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 558131 321468 558197 321469
rect 558131 321404 558132 321468
rect 558196 321404 558197 321468
rect 558131 321403 558197 321404
rect 556674 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 557294 306334
rect 556674 306014 557294 306098
rect 556674 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 557294 306014
rect 556674 270334 557294 305778
rect 556674 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 557294 270334
rect 556674 270014 557294 270098
rect 556674 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 557294 270014
rect 556674 234334 557294 269778
rect 556674 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 557294 234334
rect 556674 234014 557294 234098
rect 556674 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 557294 234014
rect 556674 198334 557294 233778
rect 556674 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 557294 198334
rect 556674 198014 557294 198098
rect 556674 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 557294 198014
rect 556674 162334 557294 197778
rect 556674 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 557294 162334
rect 556674 162014 557294 162098
rect 556674 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 557294 162014
rect 556674 126334 557294 161778
rect 556674 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 557294 126334
rect 556674 126014 557294 126098
rect 556674 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 557294 126014
rect 556674 90334 557294 125778
rect 556674 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 557294 90334
rect 556674 90014 557294 90098
rect 556674 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 557294 90014
rect 556674 54334 557294 89778
rect 556674 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 557294 54334
rect 556674 54014 557294 54098
rect 556674 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 557294 54014
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 545888 43174 546208 43206
rect 545888 42938 545930 43174
rect 546166 42938 546208 43174
rect 545888 42854 546208 42938
rect 545888 42618 545930 42854
rect 546166 42618 546208 42854
rect 545888 42586 546208 42618
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 543416 39454 543736 39486
rect 543416 39218 543458 39454
rect 543694 39218 543736 39454
rect 543416 39134 543736 39218
rect 543416 38898 543458 39134
rect 543694 38898 543736 39134
rect 543416 38866 543736 38898
rect 548361 39454 548681 39486
rect 548361 39218 548403 39454
rect 548639 39218 548681 39454
rect 548361 39134 548681 39218
rect 548361 38898 548403 39134
rect 548639 38898 548681 39134
rect 548361 38866 548681 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 7174 546134 30068
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 10894 549854 46338
rect 550833 43174 551153 43206
rect 550833 42938 550875 43174
rect 551111 42938 551153 43174
rect 550833 42854 551153 42938
rect 550833 42618 550875 42854
rect 551111 42618 551153 42854
rect 550833 42586 551153 42618
rect 555778 43174 556098 43206
rect 555778 42938 555820 43174
rect 556056 42938 556098 43174
rect 555778 42854 556098 42938
rect 555778 42618 555820 42854
rect 556056 42618 556098 42854
rect 555778 42586 556098 42618
rect 553306 39454 553626 39486
rect 553306 39218 553348 39454
rect 553584 39218 553626 39454
rect 553306 39134 553626 39218
rect 553306 38898 553348 39134
rect 553584 38898 553626 39134
rect 553306 38866 553626 38898
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 14614 553574 30068
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552954 -3226 553574 14058
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 18334 557294 53778
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 560394 51692 561014 57498
rect 564114 349774 564734 360068
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 560723 43174 561043 43206
rect 560723 42938 560765 43174
rect 561001 42938 561043 43174
rect 560723 42854 561043 42938
rect 560723 42618 560765 42854
rect 561001 42618 561043 42854
rect 560723 42586 561043 42618
rect 558251 39454 558571 39486
rect 558251 39218 558293 39454
rect 558529 39218 558571 39454
rect 558251 39134 558571 39218
rect 558251 38898 558293 39134
rect 558529 38898 558571 39134
rect 558251 38866 558571 38898
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 556674 -4186 557294 17778
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 22054 561014 30068
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 16706 594098 16942 594334
rect 17026 594098 17262 594334
rect 16706 593778 16942 594014
rect 17026 593778 17262 594014
rect 16706 558098 16942 558334
rect 17026 558098 17262 558334
rect 16706 557778 16942 558014
rect 17026 557778 17262 558014
rect 16706 522098 16942 522334
rect 17026 522098 17262 522334
rect 16706 521778 16942 522014
rect 17026 521778 17262 522014
rect 16706 486098 16942 486334
rect 17026 486098 17262 486334
rect 16706 485778 16942 486014
rect 17026 485778 17262 486014
rect 16706 450098 16942 450334
rect 17026 450098 17262 450334
rect 16706 449778 16942 450014
rect 17026 449778 17262 450014
rect 16706 414098 16942 414334
rect 17026 414098 17262 414334
rect 16706 413778 16942 414014
rect 17026 413778 17262 414014
rect 16706 378098 16942 378334
rect 17026 378098 17262 378334
rect 16706 377778 16942 378014
rect 17026 377778 17262 378014
rect 16706 342098 16942 342334
rect 17026 342098 17262 342334
rect 16706 341778 16942 342014
rect 17026 341778 17262 342014
rect 16706 306098 16942 306334
rect 17026 306098 17262 306334
rect 16706 305778 16942 306014
rect 17026 305778 17262 306014
rect 16706 270098 16942 270334
rect 17026 270098 17262 270334
rect 16706 269778 16942 270014
rect 17026 269778 17262 270014
rect 16706 234098 16942 234334
rect 17026 234098 17262 234334
rect 16706 233778 16942 234014
rect 17026 233778 17262 234014
rect 16706 198098 16942 198334
rect 17026 198098 17262 198334
rect 16706 197778 16942 198014
rect 17026 197778 17262 198014
rect 16706 162098 16942 162334
rect 17026 162098 17262 162334
rect 16706 161778 16942 162014
rect 17026 161778 17262 162014
rect 16706 126098 16942 126334
rect 17026 126098 17262 126334
rect 16706 125778 16942 126014
rect 17026 125778 17262 126014
rect 16706 90098 16942 90334
rect 17026 90098 17262 90334
rect 16706 89778 16942 90014
rect 17026 89778 17262 90014
rect 16706 54098 16942 54334
rect 17026 54098 17262 54334
rect 16706 53778 16942 54014
rect 17026 53778 17262 54014
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 20426 669818 20662 670054
rect 20746 669818 20982 670054
rect 20426 669498 20662 669734
rect 20746 669498 20982 669734
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 27866 677258 28102 677494
rect 28186 677258 28422 677494
rect 27866 676938 28102 677174
rect 28186 676938 28422 677174
rect 24250 651218 24486 651454
rect 24250 650898 24486 651134
rect 20426 633818 20662 634054
rect 20746 633818 20982 634054
rect 20426 633498 20662 633734
rect 20746 633498 20982 633734
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 63866 711322 64102 711558
rect 64186 711322 64422 711558
rect 63866 711002 64102 711238
rect 64186 711002 64422 711238
rect 63866 677258 64102 677494
rect 64186 677258 64422 677494
rect 63866 676938 64102 677174
rect 64186 676938 64422 677174
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 99866 711322 100102 711558
rect 100186 711322 100422 711558
rect 99866 711002 100102 711238
rect 100186 711002 100422 711238
rect 99866 677258 100102 677494
rect 100186 677258 100422 677494
rect 99866 676938 100102 677174
rect 100186 676938 100422 677174
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 135866 711322 136102 711558
rect 136186 711322 136422 711558
rect 135866 711002 136102 711238
rect 136186 711002 136422 711238
rect 135866 677258 136102 677494
rect 136186 677258 136422 677494
rect 135866 676938 136102 677174
rect 136186 676938 136422 677174
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 171866 711322 172102 711558
rect 172186 711322 172422 711558
rect 171866 711002 172102 711238
rect 172186 711002 172422 711238
rect 171866 677258 172102 677494
rect 172186 677258 172422 677494
rect 171866 676938 172102 677174
rect 172186 676938 172422 677174
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 207866 711322 208102 711558
rect 208186 711322 208422 711558
rect 207866 711002 208102 711238
rect 208186 711002 208422 711238
rect 207866 677258 208102 677494
rect 208186 677258 208422 677494
rect 207866 676938 208102 677174
rect 208186 676938 208422 677174
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 243866 711322 244102 711558
rect 244186 711322 244422 711558
rect 243866 711002 244102 711238
rect 244186 711002 244422 711238
rect 243866 677258 244102 677494
rect 244186 677258 244422 677494
rect 243866 676938 244102 677174
rect 244186 676938 244422 677174
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 279866 711322 280102 711558
rect 280186 711322 280422 711558
rect 279866 711002 280102 711238
rect 280186 711002 280422 711238
rect 279866 677258 280102 677494
rect 280186 677258 280422 677494
rect 279866 676938 280102 677174
rect 280186 676938 280422 677174
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 351866 711322 352102 711558
rect 352186 711322 352422 711558
rect 351866 711002 352102 711238
rect 352186 711002 352422 711238
rect 351866 677258 352102 677494
rect 352186 677258 352422 677494
rect 351866 676938 352102 677174
rect 352186 676938 352422 677174
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 39610 654938 39846 655174
rect 39610 654618 39846 654854
rect 70330 654938 70566 655174
rect 70330 654618 70566 654854
rect 101050 654938 101286 655174
rect 101050 654618 101286 654854
rect 131770 654938 132006 655174
rect 131770 654618 132006 654854
rect 162490 654938 162726 655174
rect 162490 654618 162726 654854
rect 193210 654938 193446 655174
rect 193210 654618 193446 654854
rect 223930 654938 224166 655174
rect 223930 654618 224166 654854
rect 254650 654938 254886 655174
rect 254650 654618 254886 654854
rect 285370 654938 285606 655174
rect 285370 654618 285606 654854
rect 316090 654938 316326 655174
rect 316090 654618 316326 654854
rect 346810 654938 347046 655174
rect 346810 654618 347046 654854
rect 54970 651218 55206 651454
rect 54970 650898 55206 651134
rect 85690 651218 85926 651454
rect 85690 650898 85926 651134
rect 116410 651218 116646 651454
rect 116410 650898 116646 651134
rect 147130 651218 147366 651454
rect 147130 650898 147366 651134
rect 177850 651218 178086 651454
rect 177850 650898 178086 651134
rect 208570 651218 208806 651454
rect 208570 650898 208806 651134
rect 239290 651218 239526 651454
rect 239290 650898 239526 651134
rect 270010 651218 270246 651454
rect 270010 650898 270246 651134
rect 300730 651218 300966 651454
rect 300730 650898 300966 651134
rect 331450 651218 331686 651454
rect 331450 650898 331686 651134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 27866 641258 28102 641494
rect 28186 641258 28422 641494
rect 27866 640938 28102 641174
rect 28186 640938 28422 641174
rect 24250 615218 24486 615454
rect 24250 614898 24486 615134
rect 20426 597818 20662 598054
rect 20746 597818 20982 598054
rect 20426 597498 20662 597734
rect 20746 597498 20982 597734
rect 39610 618938 39846 619174
rect 39610 618618 39846 618854
rect 70330 618938 70566 619174
rect 70330 618618 70566 618854
rect 101050 618938 101286 619174
rect 101050 618618 101286 618854
rect 131770 618938 132006 619174
rect 131770 618618 132006 618854
rect 162490 618938 162726 619174
rect 162490 618618 162726 618854
rect 193210 618938 193446 619174
rect 193210 618618 193446 618854
rect 223930 618938 224166 619174
rect 223930 618618 224166 618854
rect 254650 618938 254886 619174
rect 254650 618618 254886 618854
rect 285370 618938 285606 619174
rect 285370 618618 285606 618854
rect 316090 618938 316326 619174
rect 316090 618618 316326 618854
rect 346810 618938 347046 619174
rect 346810 618618 347046 618854
rect 54970 615218 55206 615454
rect 54970 614898 55206 615134
rect 85690 615218 85926 615454
rect 85690 614898 85926 615134
rect 116410 615218 116646 615454
rect 116410 614898 116646 615134
rect 147130 615218 147366 615454
rect 147130 614898 147366 615134
rect 177850 615218 178086 615454
rect 177850 614898 178086 615134
rect 208570 615218 208806 615454
rect 208570 614898 208806 615134
rect 239290 615218 239526 615454
rect 239290 614898 239526 615134
rect 270010 615218 270246 615454
rect 270010 614898 270246 615134
rect 300730 615218 300966 615454
rect 300730 614898 300966 615134
rect 331450 615218 331686 615454
rect 331450 614898 331686 615134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 27866 605258 28102 605494
rect 28186 605258 28422 605494
rect 27866 604938 28102 605174
rect 28186 604938 28422 605174
rect 24250 579218 24486 579454
rect 24250 578898 24486 579134
rect 20426 561818 20662 562054
rect 20746 561818 20982 562054
rect 20426 561498 20662 561734
rect 20746 561498 20982 561734
rect 39610 582938 39846 583174
rect 39610 582618 39846 582854
rect 70330 582938 70566 583174
rect 70330 582618 70566 582854
rect 101050 582938 101286 583174
rect 101050 582618 101286 582854
rect 131770 582938 132006 583174
rect 131770 582618 132006 582854
rect 162490 582938 162726 583174
rect 162490 582618 162726 582854
rect 193210 582938 193446 583174
rect 193210 582618 193446 582854
rect 223930 582938 224166 583174
rect 223930 582618 224166 582854
rect 254650 582938 254886 583174
rect 254650 582618 254886 582854
rect 285370 582938 285606 583174
rect 285370 582618 285606 582854
rect 316090 582938 316326 583174
rect 316090 582618 316326 582854
rect 346810 582938 347046 583174
rect 346810 582618 347046 582854
rect 54970 579218 55206 579454
rect 54970 578898 55206 579134
rect 85690 579218 85926 579454
rect 85690 578898 85926 579134
rect 116410 579218 116646 579454
rect 116410 578898 116646 579134
rect 147130 579218 147366 579454
rect 147130 578898 147366 579134
rect 177850 579218 178086 579454
rect 177850 578898 178086 579134
rect 208570 579218 208806 579454
rect 208570 578898 208806 579134
rect 239290 579218 239526 579454
rect 239290 578898 239526 579134
rect 270010 579218 270246 579454
rect 270010 578898 270246 579134
rect 300730 579218 300966 579454
rect 300730 578898 300966 579134
rect 331450 579218 331686 579454
rect 331450 578898 331686 579134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 27866 569258 28102 569494
rect 28186 569258 28422 569494
rect 27866 568938 28102 569174
rect 28186 568938 28422 569174
rect 24250 543218 24486 543454
rect 24250 542898 24486 543134
rect 20426 525818 20662 526054
rect 20746 525818 20982 526054
rect 20426 525498 20662 525734
rect 20746 525498 20982 525734
rect 39610 546938 39846 547174
rect 39610 546618 39846 546854
rect 70330 546938 70566 547174
rect 70330 546618 70566 546854
rect 101050 546938 101286 547174
rect 101050 546618 101286 546854
rect 131770 546938 132006 547174
rect 131770 546618 132006 546854
rect 162490 546938 162726 547174
rect 162490 546618 162726 546854
rect 193210 546938 193446 547174
rect 193210 546618 193446 546854
rect 223930 546938 224166 547174
rect 223930 546618 224166 546854
rect 254650 546938 254886 547174
rect 254650 546618 254886 546854
rect 285370 546938 285606 547174
rect 285370 546618 285606 546854
rect 316090 546938 316326 547174
rect 316090 546618 316326 546854
rect 346810 546938 347046 547174
rect 346810 546618 347046 546854
rect 54970 543218 55206 543454
rect 54970 542898 55206 543134
rect 85690 543218 85926 543454
rect 85690 542898 85926 543134
rect 116410 543218 116646 543454
rect 116410 542898 116646 543134
rect 147130 543218 147366 543454
rect 147130 542898 147366 543134
rect 177850 543218 178086 543454
rect 177850 542898 178086 543134
rect 208570 543218 208806 543454
rect 208570 542898 208806 543134
rect 239290 543218 239526 543454
rect 239290 542898 239526 543134
rect 270010 543218 270246 543454
rect 270010 542898 270246 543134
rect 300730 543218 300966 543454
rect 300730 542898 300966 543134
rect 331450 543218 331686 543454
rect 331450 542898 331686 543134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 27866 533258 28102 533494
rect 28186 533258 28422 533494
rect 27866 532938 28102 533174
rect 28186 532938 28422 533174
rect 24250 507218 24486 507454
rect 24250 506898 24486 507134
rect 20426 489818 20662 490054
rect 20746 489818 20982 490054
rect 20426 489498 20662 489734
rect 20746 489498 20982 489734
rect 39610 510938 39846 511174
rect 39610 510618 39846 510854
rect 70330 510938 70566 511174
rect 70330 510618 70566 510854
rect 101050 510938 101286 511174
rect 101050 510618 101286 510854
rect 131770 510938 132006 511174
rect 131770 510618 132006 510854
rect 162490 510938 162726 511174
rect 162490 510618 162726 510854
rect 193210 510938 193446 511174
rect 193210 510618 193446 510854
rect 223930 510938 224166 511174
rect 223930 510618 224166 510854
rect 254650 510938 254886 511174
rect 254650 510618 254886 510854
rect 285370 510938 285606 511174
rect 285370 510618 285606 510854
rect 316090 510938 316326 511174
rect 316090 510618 316326 510854
rect 346810 510938 347046 511174
rect 346810 510618 347046 510854
rect 54970 507218 55206 507454
rect 54970 506898 55206 507134
rect 85690 507218 85926 507454
rect 85690 506898 85926 507134
rect 116410 507218 116646 507454
rect 116410 506898 116646 507134
rect 147130 507218 147366 507454
rect 147130 506898 147366 507134
rect 177850 507218 178086 507454
rect 177850 506898 178086 507134
rect 208570 507218 208806 507454
rect 208570 506898 208806 507134
rect 239290 507218 239526 507454
rect 239290 506898 239526 507134
rect 270010 507218 270246 507454
rect 270010 506898 270246 507134
rect 300730 507218 300966 507454
rect 300730 506898 300966 507134
rect 331450 507218 331686 507454
rect 331450 506898 331686 507134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 27866 497258 28102 497494
rect 28186 497258 28422 497494
rect 27866 496938 28102 497174
rect 28186 496938 28422 497174
rect 24250 471218 24486 471454
rect 24250 470898 24486 471134
rect 20426 453818 20662 454054
rect 20746 453818 20982 454054
rect 20426 453498 20662 453734
rect 20746 453498 20982 453734
rect 39610 474938 39846 475174
rect 39610 474618 39846 474854
rect 70330 474938 70566 475174
rect 70330 474618 70566 474854
rect 101050 474938 101286 475174
rect 101050 474618 101286 474854
rect 131770 474938 132006 475174
rect 131770 474618 132006 474854
rect 162490 474938 162726 475174
rect 162490 474618 162726 474854
rect 193210 474938 193446 475174
rect 193210 474618 193446 474854
rect 223930 474938 224166 475174
rect 223930 474618 224166 474854
rect 254650 474938 254886 475174
rect 254650 474618 254886 474854
rect 285370 474938 285606 475174
rect 285370 474618 285606 474854
rect 316090 474938 316326 475174
rect 316090 474618 316326 474854
rect 346810 474938 347046 475174
rect 346810 474618 347046 474854
rect 54970 471218 55206 471454
rect 54970 470898 55206 471134
rect 85690 471218 85926 471454
rect 85690 470898 85926 471134
rect 116410 471218 116646 471454
rect 116410 470898 116646 471134
rect 147130 471218 147366 471454
rect 147130 470898 147366 471134
rect 177850 471218 178086 471454
rect 177850 470898 178086 471134
rect 208570 471218 208806 471454
rect 208570 470898 208806 471134
rect 239290 471218 239526 471454
rect 239290 470898 239526 471134
rect 270010 471218 270246 471454
rect 270010 470898 270246 471134
rect 300730 471218 300966 471454
rect 300730 470898 300966 471134
rect 331450 471218 331686 471454
rect 331450 470898 331686 471134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 27866 461258 28102 461494
rect 28186 461258 28422 461494
rect 27866 460938 28102 461174
rect 28186 460938 28422 461174
rect 24250 435218 24486 435454
rect 24250 434898 24486 435134
rect 20426 417818 20662 418054
rect 20746 417818 20982 418054
rect 20426 417498 20662 417734
rect 20746 417498 20982 417734
rect 39610 438938 39846 439174
rect 39610 438618 39846 438854
rect 70330 438938 70566 439174
rect 70330 438618 70566 438854
rect 101050 438938 101286 439174
rect 101050 438618 101286 438854
rect 131770 438938 132006 439174
rect 131770 438618 132006 438854
rect 162490 438938 162726 439174
rect 162490 438618 162726 438854
rect 193210 438938 193446 439174
rect 193210 438618 193446 438854
rect 223930 438938 224166 439174
rect 223930 438618 224166 438854
rect 254650 438938 254886 439174
rect 254650 438618 254886 438854
rect 285370 438938 285606 439174
rect 285370 438618 285606 438854
rect 316090 438938 316326 439174
rect 316090 438618 316326 438854
rect 346810 438938 347046 439174
rect 346810 438618 347046 438854
rect 54970 435218 55206 435454
rect 54970 434898 55206 435134
rect 85690 435218 85926 435454
rect 85690 434898 85926 435134
rect 116410 435218 116646 435454
rect 116410 434898 116646 435134
rect 147130 435218 147366 435454
rect 147130 434898 147366 435134
rect 177850 435218 178086 435454
rect 177850 434898 178086 435134
rect 208570 435218 208806 435454
rect 208570 434898 208806 435134
rect 239290 435218 239526 435454
rect 239290 434898 239526 435134
rect 270010 435218 270246 435454
rect 270010 434898 270246 435134
rect 300730 435218 300966 435454
rect 300730 434898 300966 435134
rect 331450 435218 331686 435454
rect 331450 434898 331686 435134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 27866 425258 28102 425494
rect 28186 425258 28422 425494
rect 27866 424938 28102 425174
rect 28186 424938 28422 425174
rect 24250 399218 24486 399454
rect 24250 398898 24486 399134
rect 20426 381818 20662 382054
rect 20746 381818 20982 382054
rect 20426 381498 20662 381734
rect 20746 381498 20982 381734
rect 39610 402938 39846 403174
rect 39610 402618 39846 402854
rect 70330 402938 70566 403174
rect 70330 402618 70566 402854
rect 101050 402938 101286 403174
rect 101050 402618 101286 402854
rect 131770 402938 132006 403174
rect 131770 402618 132006 402854
rect 162490 402938 162726 403174
rect 162490 402618 162726 402854
rect 193210 402938 193446 403174
rect 193210 402618 193446 402854
rect 223930 402938 224166 403174
rect 223930 402618 224166 402854
rect 254650 402938 254886 403174
rect 254650 402618 254886 402854
rect 285370 402938 285606 403174
rect 285370 402618 285606 402854
rect 316090 402938 316326 403174
rect 316090 402618 316326 402854
rect 346810 402938 347046 403174
rect 346810 402618 347046 402854
rect 54970 399218 55206 399454
rect 54970 398898 55206 399134
rect 85690 399218 85926 399454
rect 85690 398898 85926 399134
rect 116410 399218 116646 399454
rect 116410 398898 116646 399134
rect 147130 399218 147366 399454
rect 147130 398898 147366 399134
rect 177850 399218 178086 399454
rect 177850 398898 178086 399134
rect 208570 399218 208806 399454
rect 208570 398898 208806 399134
rect 239290 399218 239526 399454
rect 239290 398898 239526 399134
rect 270010 399218 270246 399454
rect 270010 398898 270246 399134
rect 300730 399218 300966 399454
rect 300730 398898 300966 399134
rect 331450 399218 331686 399454
rect 331450 398898 331686 399134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 27866 389258 28102 389494
rect 28186 389258 28422 389494
rect 27866 388938 28102 389174
rect 28186 388938 28422 389174
rect 24250 363218 24486 363454
rect 24250 362898 24486 363134
rect 20426 345818 20662 346054
rect 20746 345818 20982 346054
rect 20426 345498 20662 345734
rect 20746 345498 20982 345734
rect 39610 366938 39846 367174
rect 39610 366618 39846 366854
rect 70330 366938 70566 367174
rect 70330 366618 70566 366854
rect 101050 366938 101286 367174
rect 101050 366618 101286 366854
rect 131770 366938 132006 367174
rect 131770 366618 132006 366854
rect 162490 366938 162726 367174
rect 162490 366618 162726 366854
rect 193210 366938 193446 367174
rect 193210 366618 193446 366854
rect 223930 366938 224166 367174
rect 223930 366618 224166 366854
rect 254650 366938 254886 367174
rect 254650 366618 254886 366854
rect 285370 366938 285606 367174
rect 285370 366618 285606 366854
rect 316090 366938 316326 367174
rect 316090 366618 316326 366854
rect 346810 366938 347046 367174
rect 346810 366618 347046 366854
rect 54970 363218 55206 363454
rect 54970 362898 55206 363134
rect 85690 363218 85926 363454
rect 85690 362898 85926 363134
rect 116410 363218 116646 363454
rect 116410 362898 116646 363134
rect 147130 363218 147366 363454
rect 147130 362898 147366 363134
rect 177850 363218 178086 363454
rect 177850 362898 178086 363134
rect 208570 363218 208806 363454
rect 208570 362898 208806 363134
rect 239290 363218 239526 363454
rect 239290 362898 239526 363134
rect 270010 363218 270246 363454
rect 270010 362898 270246 363134
rect 300730 363218 300966 363454
rect 300730 362898 300966 363134
rect 331450 363218 331686 363454
rect 331450 362898 331686 363134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 27866 353258 28102 353494
rect 28186 353258 28422 353494
rect 27866 352938 28102 353174
rect 28186 352938 28422 353174
rect 24250 327218 24486 327454
rect 24250 326898 24486 327134
rect 20426 309818 20662 310054
rect 20746 309818 20982 310054
rect 20426 309498 20662 309734
rect 20746 309498 20982 309734
rect 39610 330938 39846 331174
rect 39610 330618 39846 330854
rect 70330 330938 70566 331174
rect 70330 330618 70566 330854
rect 101050 330938 101286 331174
rect 101050 330618 101286 330854
rect 131770 330938 132006 331174
rect 131770 330618 132006 330854
rect 162490 330938 162726 331174
rect 162490 330618 162726 330854
rect 193210 330938 193446 331174
rect 193210 330618 193446 330854
rect 223930 330938 224166 331174
rect 223930 330618 224166 330854
rect 254650 330938 254886 331174
rect 254650 330618 254886 330854
rect 285370 330938 285606 331174
rect 285370 330618 285606 330854
rect 316090 330938 316326 331174
rect 316090 330618 316326 330854
rect 346810 330938 347046 331174
rect 346810 330618 347046 330854
rect 54970 327218 55206 327454
rect 54970 326898 55206 327134
rect 85690 327218 85926 327454
rect 85690 326898 85926 327134
rect 116410 327218 116646 327454
rect 116410 326898 116646 327134
rect 147130 327218 147366 327454
rect 147130 326898 147366 327134
rect 177850 327218 178086 327454
rect 177850 326898 178086 327134
rect 208570 327218 208806 327454
rect 208570 326898 208806 327134
rect 239290 327218 239526 327454
rect 239290 326898 239526 327134
rect 270010 327218 270246 327454
rect 270010 326898 270246 327134
rect 300730 327218 300966 327454
rect 300730 326898 300966 327134
rect 331450 327218 331686 327454
rect 331450 326898 331686 327134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 27866 317258 28102 317494
rect 28186 317258 28422 317494
rect 27866 316938 28102 317174
rect 28186 316938 28422 317174
rect 24250 291218 24486 291454
rect 24250 290898 24486 291134
rect 20426 273818 20662 274054
rect 20746 273818 20982 274054
rect 20426 273498 20662 273734
rect 20746 273498 20982 273734
rect 39610 294938 39846 295174
rect 39610 294618 39846 294854
rect 70330 294938 70566 295174
rect 70330 294618 70566 294854
rect 101050 294938 101286 295174
rect 101050 294618 101286 294854
rect 131770 294938 132006 295174
rect 131770 294618 132006 294854
rect 162490 294938 162726 295174
rect 162490 294618 162726 294854
rect 193210 294938 193446 295174
rect 193210 294618 193446 294854
rect 223930 294938 224166 295174
rect 223930 294618 224166 294854
rect 254650 294938 254886 295174
rect 254650 294618 254886 294854
rect 285370 294938 285606 295174
rect 285370 294618 285606 294854
rect 316090 294938 316326 295174
rect 316090 294618 316326 294854
rect 346810 294938 347046 295174
rect 346810 294618 347046 294854
rect 54970 291218 55206 291454
rect 54970 290898 55206 291134
rect 85690 291218 85926 291454
rect 85690 290898 85926 291134
rect 116410 291218 116646 291454
rect 116410 290898 116646 291134
rect 147130 291218 147366 291454
rect 147130 290898 147366 291134
rect 177850 291218 178086 291454
rect 177850 290898 178086 291134
rect 208570 291218 208806 291454
rect 208570 290898 208806 291134
rect 239290 291218 239526 291454
rect 239290 290898 239526 291134
rect 270010 291218 270246 291454
rect 270010 290898 270246 291134
rect 300730 291218 300966 291454
rect 300730 290898 300966 291134
rect 331450 291218 331686 291454
rect 331450 290898 331686 291134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 27866 281258 28102 281494
rect 28186 281258 28422 281494
rect 27866 280938 28102 281174
rect 28186 280938 28422 281174
rect 24250 255218 24486 255454
rect 24250 254898 24486 255134
rect 20426 237818 20662 238054
rect 20746 237818 20982 238054
rect 20426 237498 20662 237734
rect 20746 237498 20982 237734
rect 39610 258938 39846 259174
rect 39610 258618 39846 258854
rect 70330 258938 70566 259174
rect 70330 258618 70566 258854
rect 101050 258938 101286 259174
rect 101050 258618 101286 258854
rect 131770 258938 132006 259174
rect 131770 258618 132006 258854
rect 162490 258938 162726 259174
rect 162490 258618 162726 258854
rect 193210 258938 193446 259174
rect 193210 258618 193446 258854
rect 223930 258938 224166 259174
rect 223930 258618 224166 258854
rect 254650 258938 254886 259174
rect 254650 258618 254886 258854
rect 285370 258938 285606 259174
rect 285370 258618 285606 258854
rect 316090 258938 316326 259174
rect 316090 258618 316326 258854
rect 346810 258938 347046 259174
rect 346810 258618 347046 258854
rect 54970 255218 55206 255454
rect 54970 254898 55206 255134
rect 85690 255218 85926 255454
rect 85690 254898 85926 255134
rect 116410 255218 116646 255454
rect 116410 254898 116646 255134
rect 147130 255218 147366 255454
rect 147130 254898 147366 255134
rect 177850 255218 178086 255454
rect 177850 254898 178086 255134
rect 208570 255218 208806 255454
rect 208570 254898 208806 255134
rect 239290 255218 239526 255454
rect 239290 254898 239526 255134
rect 270010 255218 270246 255454
rect 270010 254898 270246 255134
rect 300730 255218 300966 255454
rect 300730 254898 300966 255134
rect 331450 255218 331686 255454
rect 331450 254898 331686 255134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 27866 245258 28102 245494
rect 28186 245258 28422 245494
rect 27866 244938 28102 245174
rect 28186 244938 28422 245174
rect 24250 219218 24486 219454
rect 24250 218898 24486 219134
rect 20426 201818 20662 202054
rect 20746 201818 20982 202054
rect 20426 201498 20662 201734
rect 20746 201498 20982 201734
rect 39610 222938 39846 223174
rect 39610 222618 39846 222854
rect 70330 222938 70566 223174
rect 70330 222618 70566 222854
rect 101050 222938 101286 223174
rect 101050 222618 101286 222854
rect 131770 222938 132006 223174
rect 131770 222618 132006 222854
rect 162490 222938 162726 223174
rect 162490 222618 162726 222854
rect 193210 222938 193446 223174
rect 193210 222618 193446 222854
rect 223930 222938 224166 223174
rect 223930 222618 224166 222854
rect 254650 222938 254886 223174
rect 254650 222618 254886 222854
rect 285370 222938 285606 223174
rect 285370 222618 285606 222854
rect 316090 222938 316326 223174
rect 316090 222618 316326 222854
rect 346810 222938 347046 223174
rect 346810 222618 347046 222854
rect 54970 219218 55206 219454
rect 54970 218898 55206 219134
rect 85690 219218 85926 219454
rect 85690 218898 85926 219134
rect 116410 219218 116646 219454
rect 116410 218898 116646 219134
rect 147130 219218 147366 219454
rect 147130 218898 147366 219134
rect 177850 219218 178086 219454
rect 177850 218898 178086 219134
rect 208570 219218 208806 219454
rect 208570 218898 208806 219134
rect 239290 219218 239526 219454
rect 239290 218898 239526 219134
rect 270010 219218 270246 219454
rect 270010 218898 270246 219134
rect 300730 219218 300966 219454
rect 300730 218898 300966 219134
rect 331450 219218 331686 219454
rect 331450 218898 331686 219134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 27866 209258 28102 209494
rect 28186 209258 28422 209494
rect 27866 208938 28102 209174
rect 28186 208938 28422 209174
rect 24250 183218 24486 183454
rect 24250 182898 24486 183134
rect 20426 165818 20662 166054
rect 20746 165818 20982 166054
rect 20426 165498 20662 165734
rect 20746 165498 20982 165734
rect 39610 186938 39846 187174
rect 39610 186618 39846 186854
rect 70330 186938 70566 187174
rect 70330 186618 70566 186854
rect 101050 186938 101286 187174
rect 101050 186618 101286 186854
rect 131770 186938 132006 187174
rect 131770 186618 132006 186854
rect 162490 186938 162726 187174
rect 162490 186618 162726 186854
rect 193210 186938 193446 187174
rect 193210 186618 193446 186854
rect 223930 186938 224166 187174
rect 223930 186618 224166 186854
rect 254650 186938 254886 187174
rect 254650 186618 254886 186854
rect 285370 186938 285606 187174
rect 285370 186618 285606 186854
rect 316090 186938 316326 187174
rect 316090 186618 316326 186854
rect 346810 186938 347046 187174
rect 346810 186618 347046 186854
rect 54970 183218 55206 183454
rect 54970 182898 55206 183134
rect 85690 183218 85926 183454
rect 85690 182898 85926 183134
rect 116410 183218 116646 183454
rect 116410 182898 116646 183134
rect 147130 183218 147366 183454
rect 147130 182898 147366 183134
rect 177850 183218 178086 183454
rect 177850 182898 178086 183134
rect 208570 183218 208806 183454
rect 208570 182898 208806 183134
rect 239290 183218 239526 183454
rect 239290 182898 239526 183134
rect 270010 183218 270246 183454
rect 270010 182898 270246 183134
rect 300730 183218 300966 183454
rect 300730 182898 300966 183134
rect 331450 183218 331686 183454
rect 331450 182898 331686 183134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 27866 173258 28102 173494
rect 28186 173258 28422 173494
rect 27866 172938 28102 173174
rect 28186 172938 28422 173174
rect 24250 147218 24486 147454
rect 24250 146898 24486 147134
rect 20426 129818 20662 130054
rect 20746 129818 20982 130054
rect 20426 129498 20662 129734
rect 20746 129498 20982 129734
rect 39610 150938 39846 151174
rect 39610 150618 39846 150854
rect 70330 150938 70566 151174
rect 70330 150618 70566 150854
rect 101050 150938 101286 151174
rect 101050 150618 101286 150854
rect 131770 150938 132006 151174
rect 131770 150618 132006 150854
rect 162490 150938 162726 151174
rect 162490 150618 162726 150854
rect 193210 150938 193446 151174
rect 193210 150618 193446 150854
rect 223930 150938 224166 151174
rect 223930 150618 224166 150854
rect 254650 150938 254886 151174
rect 254650 150618 254886 150854
rect 285370 150938 285606 151174
rect 285370 150618 285606 150854
rect 316090 150938 316326 151174
rect 316090 150618 316326 150854
rect 346810 150938 347046 151174
rect 346810 150618 347046 150854
rect 54970 147218 55206 147454
rect 54970 146898 55206 147134
rect 85690 147218 85926 147454
rect 85690 146898 85926 147134
rect 116410 147218 116646 147454
rect 116410 146898 116646 147134
rect 147130 147218 147366 147454
rect 147130 146898 147366 147134
rect 177850 147218 178086 147454
rect 177850 146898 178086 147134
rect 208570 147218 208806 147454
rect 208570 146898 208806 147134
rect 239290 147218 239526 147454
rect 239290 146898 239526 147134
rect 270010 147218 270246 147454
rect 270010 146898 270246 147134
rect 300730 147218 300966 147454
rect 300730 146898 300966 147134
rect 331450 147218 331686 147454
rect 331450 146898 331686 147134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 27866 137258 28102 137494
rect 28186 137258 28422 137494
rect 27866 136938 28102 137174
rect 28186 136938 28422 137174
rect 24250 111218 24486 111454
rect 24250 110898 24486 111134
rect 20426 93818 20662 94054
rect 20746 93818 20982 94054
rect 20426 93498 20662 93734
rect 20746 93498 20982 93734
rect 39610 114938 39846 115174
rect 39610 114618 39846 114854
rect 70330 114938 70566 115174
rect 70330 114618 70566 114854
rect 101050 114938 101286 115174
rect 101050 114618 101286 114854
rect 131770 114938 132006 115174
rect 131770 114618 132006 114854
rect 162490 114938 162726 115174
rect 162490 114618 162726 114854
rect 193210 114938 193446 115174
rect 193210 114618 193446 114854
rect 223930 114938 224166 115174
rect 223930 114618 224166 114854
rect 254650 114938 254886 115174
rect 254650 114618 254886 114854
rect 285370 114938 285606 115174
rect 285370 114618 285606 114854
rect 316090 114938 316326 115174
rect 316090 114618 316326 114854
rect 346810 114938 347046 115174
rect 346810 114618 347046 114854
rect 54970 111218 55206 111454
rect 54970 110898 55206 111134
rect 85690 111218 85926 111454
rect 85690 110898 85926 111134
rect 116410 111218 116646 111454
rect 116410 110898 116646 111134
rect 147130 111218 147366 111454
rect 147130 110898 147366 111134
rect 177850 111218 178086 111454
rect 177850 110898 178086 111134
rect 208570 111218 208806 111454
rect 208570 110898 208806 111134
rect 239290 111218 239526 111454
rect 239290 110898 239526 111134
rect 270010 111218 270246 111454
rect 270010 110898 270246 111134
rect 300730 111218 300966 111454
rect 300730 110898 300966 111134
rect 331450 111218 331686 111454
rect 331450 110898 331686 111134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 27866 101258 28102 101494
rect 28186 101258 28422 101494
rect 27866 100938 28102 101174
rect 28186 100938 28422 101174
rect 24250 75218 24486 75454
rect 24250 74898 24486 75134
rect 20426 57818 20662 58054
rect 20746 57818 20982 58054
rect 20426 57498 20662 57734
rect 20746 57498 20982 57734
rect 39610 78938 39846 79174
rect 39610 78618 39846 78854
rect 70330 78938 70566 79174
rect 70330 78618 70566 78854
rect 101050 78938 101286 79174
rect 101050 78618 101286 78854
rect 131770 78938 132006 79174
rect 131770 78618 132006 78854
rect 162490 78938 162726 79174
rect 162490 78618 162726 78854
rect 193210 78938 193446 79174
rect 193210 78618 193446 78854
rect 223930 78938 224166 79174
rect 223930 78618 224166 78854
rect 254650 78938 254886 79174
rect 254650 78618 254886 78854
rect 285370 78938 285606 79174
rect 285370 78618 285606 78854
rect 316090 78938 316326 79174
rect 316090 78618 316326 78854
rect 346810 78938 347046 79174
rect 346810 78618 347046 78854
rect 54970 75218 55206 75454
rect 54970 74898 55206 75134
rect 85690 75218 85926 75454
rect 85690 74898 85926 75134
rect 116410 75218 116646 75454
rect 116410 74898 116646 75134
rect 147130 75218 147366 75454
rect 147130 74898 147366 75134
rect 177850 75218 178086 75454
rect 177850 74898 178086 75134
rect 208570 75218 208806 75454
rect 208570 74898 208806 75134
rect 239290 75218 239526 75454
rect 239290 74898 239526 75134
rect 270010 75218 270246 75454
rect 270010 74898 270246 75134
rect 300730 75218 300966 75454
rect 300730 74898 300966 75134
rect 331450 75218 331686 75454
rect 331450 74898 331686 75134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 27866 65258 28102 65494
rect 28186 65258 28422 65494
rect 27866 64938 28102 65174
rect 28186 64938 28422 65174
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 20426 -5382 20662 -5146
rect 20746 -5382 20982 -5146
rect 20426 -5702 20662 -5466
rect 20746 -5702 20982 -5466
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 24146 -6342 24382 -6106
rect 24466 -6342 24702 -6106
rect 24146 -6662 24382 -6426
rect 24466 -6662 24702 -6426
rect 27866 29258 28102 29494
rect 28186 29258 28422 29494
rect 27866 28938 28102 29174
rect 28186 28938 28422 29174
rect 27866 -7302 28102 -7066
rect 28186 -7302 28422 -7066
rect 27866 -7622 28102 -7386
rect 28186 -7622 28422 -7386
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 48986 -3462 49222 -3226
rect 49306 -3462 49542 -3226
rect 48986 -3782 49222 -3546
rect 49306 -3782 49542 -3546
rect 52706 18098 52942 18334
rect 53026 18098 53262 18334
rect 52706 17778 52942 18014
rect 53026 17778 53262 18014
rect 52706 -4422 52942 -4186
rect 53026 -4422 53262 -4186
rect 52706 -4742 52942 -4506
rect 53026 -4742 53262 -4506
rect 56426 21818 56662 22054
rect 56746 21818 56982 22054
rect 56426 21498 56662 21734
rect 56746 21498 56982 21734
rect 56426 -5382 56662 -5146
rect 56746 -5382 56982 -5146
rect 56426 -5702 56662 -5466
rect 56746 -5702 56982 -5466
rect 60146 25538 60382 25774
rect 60466 25538 60702 25774
rect 60146 25218 60382 25454
rect 60466 25218 60702 25454
rect 60146 -6342 60382 -6106
rect 60466 -6342 60702 -6106
rect 60146 -6662 60382 -6426
rect 60466 -6662 60702 -6426
rect 63866 29258 64102 29494
rect 64186 29258 64422 29494
rect 63866 28938 64102 29174
rect 64186 28938 64422 29174
rect 63866 -7302 64102 -7066
rect 64186 -7302 64422 -7066
rect 63866 -7622 64102 -7386
rect 64186 -7622 64422 -7386
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 84986 -3462 85222 -3226
rect 85306 -3462 85542 -3226
rect 84986 -3782 85222 -3546
rect 85306 -3782 85542 -3546
rect 88706 18098 88942 18334
rect 89026 18098 89262 18334
rect 88706 17778 88942 18014
rect 89026 17778 89262 18014
rect 88706 -4422 88942 -4186
rect 89026 -4422 89262 -4186
rect 88706 -4742 88942 -4506
rect 89026 -4742 89262 -4506
rect 92426 21818 92662 22054
rect 92746 21818 92982 22054
rect 92426 21498 92662 21734
rect 92746 21498 92982 21734
rect 92426 -5382 92662 -5146
rect 92746 -5382 92982 -5146
rect 92426 -5702 92662 -5466
rect 92746 -5702 92982 -5466
rect 96146 25538 96382 25774
rect 96466 25538 96702 25774
rect 96146 25218 96382 25454
rect 96466 25218 96702 25454
rect 96146 -6342 96382 -6106
rect 96466 -6342 96702 -6106
rect 96146 -6662 96382 -6426
rect 96466 -6662 96702 -6426
rect 99866 29258 100102 29494
rect 100186 29258 100422 29494
rect 99866 28938 100102 29174
rect 100186 28938 100422 29174
rect 99866 -7302 100102 -7066
rect 100186 -7302 100422 -7066
rect 99866 -7622 100102 -7386
rect 100186 -7622 100422 -7386
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 120986 -3462 121222 -3226
rect 121306 -3462 121542 -3226
rect 120986 -3782 121222 -3546
rect 121306 -3782 121542 -3546
rect 124706 18098 124942 18334
rect 125026 18098 125262 18334
rect 124706 17778 124942 18014
rect 125026 17778 125262 18014
rect 124706 -4422 124942 -4186
rect 125026 -4422 125262 -4186
rect 124706 -4742 124942 -4506
rect 125026 -4742 125262 -4506
rect 128426 21818 128662 22054
rect 128746 21818 128982 22054
rect 128426 21498 128662 21734
rect 128746 21498 128982 21734
rect 128426 -5382 128662 -5146
rect 128746 -5382 128982 -5146
rect 128426 -5702 128662 -5466
rect 128746 -5702 128982 -5466
rect 132146 25538 132382 25774
rect 132466 25538 132702 25774
rect 132146 25218 132382 25454
rect 132466 25218 132702 25454
rect 132146 -6342 132382 -6106
rect 132466 -6342 132702 -6106
rect 132146 -6662 132382 -6426
rect 132466 -6662 132702 -6426
rect 135866 29258 136102 29494
rect 136186 29258 136422 29494
rect 135866 28938 136102 29174
rect 136186 28938 136422 29174
rect 135866 -7302 136102 -7066
rect 136186 -7302 136422 -7066
rect 135866 -7622 136102 -7386
rect 136186 -7622 136422 -7386
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 156986 -3462 157222 -3226
rect 157306 -3462 157542 -3226
rect 156986 -3782 157222 -3546
rect 157306 -3782 157542 -3546
rect 160706 18098 160942 18334
rect 161026 18098 161262 18334
rect 160706 17778 160942 18014
rect 161026 17778 161262 18014
rect 160706 -4422 160942 -4186
rect 161026 -4422 161262 -4186
rect 160706 -4742 160942 -4506
rect 161026 -4742 161262 -4506
rect 164426 21818 164662 22054
rect 164746 21818 164982 22054
rect 164426 21498 164662 21734
rect 164746 21498 164982 21734
rect 164426 -5382 164662 -5146
rect 164746 -5382 164982 -5146
rect 164426 -5702 164662 -5466
rect 164746 -5702 164982 -5466
rect 168146 25538 168382 25774
rect 168466 25538 168702 25774
rect 168146 25218 168382 25454
rect 168466 25218 168702 25454
rect 168146 -6342 168382 -6106
rect 168466 -6342 168702 -6106
rect 168146 -6662 168382 -6426
rect 168466 -6662 168702 -6426
rect 171866 29258 172102 29494
rect 172186 29258 172422 29494
rect 171866 28938 172102 29174
rect 172186 28938 172422 29174
rect 171866 -7302 172102 -7066
rect 172186 -7302 172422 -7066
rect 171866 -7622 172102 -7386
rect 172186 -7622 172422 -7386
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 192986 -3462 193222 -3226
rect 193306 -3462 193542 -3226
rect 192986 -3782 193222 -3546
rect 193306 -3782 193542 -3546
rect 196706 18098 196942 18334
rect 197026 18098 197262 18334
rect 196706 17778 196942 18014
rect 197026 17778 197262 18014
rect 196706 -4422 196942 -4186
rect 197026 -4422 197262 -4186
rect 196706 -4742 196942 -4506
rect 197026 -4742 197262 -4506
rect 200426 21818 200662 22054
rect 200746 21818 200982 22054
rect 200426 21498 200662 21734
rect 200746 21498 200982 21734
rect 200426 -5382 200662 -5146
rect 200746 -5382 200982 -5146
rect 200426 -5702 200662 -5466
rect 200746 -5702 200982 -5466
rect 204146 25538 204382 25774
rect 204466 25538 204702 25774
rect 204146 25218 204382 25454
rect 204466 25218 204702 25454
rect 204146 -6342 204382 -6106
rect 204466 -6342 204702 -6106
rect 204146 -6662 204382 -6426
rect 204466 -6662 204702 -6426
rect 207866 29258 208102 29494
rect 208186 29258 208422 29494
rect 207866 28938 208102 29174
rect 208186 28938 208422 29174
rect 207866 -7302 208102 -7066
rect 208186 -7302 208422 -7066
rect 207866 -7622 208102 -7386
rect 208186 -7622 208422 -7386
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 228986 -3462 229222 -3226
rect 229306 -3462 229542 -3226
rect 228986 -3782 229222 -3546
rect 229306 -3782 229542 -3546
rect 232706 18098 232942 18334
rect 233026 18098 233262 18334
rect 232706 17778 232942 18014
rect 233026 17778 233262 18014
rect 232706 -4422 232942 -4186
rect 233026 -4422 233262 -4186
rect 232706 -4742 232942 -4506
rect 233026 -4742 233262 -4506
rect 236426 21818 236662 22054
rect 236746 21818 236982 22054
rect 236426 21498 236662 21734
rect 236746 21498 236982 21734
rect 236426 -5382 236662 -5146
rect 236746 -5382 236982 -5146
rect 236426 -5702 236662 -5466
rect 236746 -5702 236982 -5466
rect 240146 25538 240382 25774
rect 240466 25538 240702 25774
rect 240146 25218 240382 25454
rect 240466 25218 240702 25454
rect 240146 -6342 240382 -6106
rect 240466 -6342 240702 -6106
rect 240146 -6662 240382 -6426
rect 240466 -6662 240702 -6426
rect 243866 29258 244102 29494
rect 244186 29258 244422 29494
rect 243866 28938 244102 29174
rect 244186 28938 244422 29174
rect 243866 -7302 244102 -7066
rect 244186 -7302 244422 -7066
rect 243866 -7622 244102 -7386
rect 244186 -7622 244422 -7386
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 264986 -3462 265222 -3226
rect 265306 -3462 265542 -3226
rect 264986 -3782 265222 -3546
rect 265306 -3782 265542 -3546
rect 268706 18098 268942 18334
rect 269026 18098 269262 18334
rect 268706 17778 268942 18014
rect 269026 17778 269262 18014
rect 268706 -4422 268942 -4186
rect 269026 -4422 269262 -4186
rect 268706 -4742 268942 -4506
rect 269026 -4742 269262 -4506
rect 272426 21818 272662 22054
rect 272746 21818 272982 22054
rect 272426 21498 272662 21734
rect 272746 21498 272982 21734
rect 272426 -5382 272662 -5146
rect 272746 -5382 272982 -5146
rect 272426 -5702 272662 -5466
rect 272746 -5702 272982 -5466
rect 276146 25538 276382 25774
rect 276466 25538 276702 25774
rect 276146 25218 276382 25454
rect 276466 25218 276702 25454
rect 276146 -6342 276382 -6106
rect 276466 -6342 276702 -6106
rect 276146 -6662 276382 -6426
rect 276466 -6662 276702 -6426
rect 279866 29258 280102 29494
rect 280186 29258 280422 29494
rect 279866 28938 280102 29174
rect 280186 28938 280422 29174
rect 279866 -7302 280102 -7066
rect 280186 -7302 280422 -7066
rect 279866 -7622 280102 -7386
rect 280186 -7622 280422 -7386
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 300986 -3462 301222 -3226
rect 301306 -3462 301542 -3226
rect 300986 -3782 301222 -3546
rect 301306 -3782 301542 -3546
rect 304706 18098 304942 18334
rect 305026 18098 305262 18334
rect 304706 17778 304942 18014
rect 305026 17778 305262 18014
rect 304706 -4422 304942 -4186
rect 305026 -4422 305262 -4186
rect 304706 -4742 304942 -4506
rect 305026 -4742 305262 -4506
rect 308426 21818 308662 22054
rect 308746 21818 308982 22054
rect 308426 21498 308662 21734
rect 308746 21498 308982 21734
rect 308426 -5382 308662 -5146
rect 308746 -5382 308982 -5146
rect 308426 -5702 308662 -5466
rect 308746 -5702 308982 -5466
rect 312146 25538 312382 25774
rect 312466 25538 312702 25774
rect 312146 25218 312382 25454
rect 312466 25218 312702 25454
rect 312146 -6342 312382 -6106
rect 312466 -6342 312702 -6106
rect 312146 -6662 312382 -6426
rect 312466 -6662 312702 -6426
rect 315866 29258 316102 29494
rect 316186 29258 316422 29494
rect 315866 28938 316102 29174
rect 316186 28938 316422 29174
rect 315866 -7302 316102 -7066
rect 316186 -7302 316422 -7066
rect 315866 -7622 316102 -7386
rect 316186 -7622 316422 -7386
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 336986 -3462 337222 -3226
rect 337306 -3462 337542 -3226
rect 336986 -3782 337222 -3546
rect 337306 -3782 337542 -3546
rect 340706 18098 340942 18334
rect 341026 18098 341262 18334
rect 340706 17778 340942 18014
rect 341026 17778 341262 18014
rect 340706 -4422 340942 -4186
rect 341026 -4422 341262 -4186
rect 340706 -4742 340942 -4506
rect 341026 -4742 341262 -4506
rect 344426 21818 344662 22054
rect 344746 21818 344982 22054
rect 344426 21498 344662 21734
rect 344746 21498 344982 21734
rect 344426 -5382 344662 -5146
rect 344746 -5382 344982 -5146
rect 344426 -5702 344662 -5466
rect 344746 -5702 344982 -5466
rect 348146 25538 348382 25774
rect 348466 25538 348702 25774
rect 348146 25218 348382 25454
rect 348466 25218 348702 25454
rect 348146 -6342 348382 -6106
rect 348466 -6342 348702 -6106
rect 348146 -6662 348382 -6426
rect 348466 -6662 348702 -6426
rect 351866 29258 352102 29494
rect 352186 29258 352422 29494
rect 351866 28938 352102 29174
rect 352186 28938 352422 29174
rect 351866 -7302 352102 -7066
rect 352186 -7302 352422 -7066
rect 351866 -7622 352102 -7386
rect 352186 -7622 352422 -7386
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 372986 -3462 373222 -3226
rect 373306 -3462 373542 -3226
rect 372986 -3782 373222 -3546
rect 373306 -3782 373542 -3546
rect 376706 708442 376942 708678
rect 377026 708442 377262 708678
rect 376706 708122 376942 708358
rect 377026 708122 377262 708358
rect 376706 666098 376942 666334
rect 377026 666098 377262 666334
rect 376706 665778 376942 666014
rect 377026 665778 377262 666014
rect 376706 630098 376942 630334
rect 377026 630098 377262 630334
rect 376706 629778 376942 630014
rect 377026 629778 377262 630014
rect 376706 594098 376942 594334
rect 377026 594098 377262 594334
rect 376706 593778 376942 594014
rect 377026 593778 377262 594014
rect 376706 558098 376942 558334
rect 377026 558098 377262 558334
rect 376706 557778 376942 558014
rect 377026 557778 377262 558014
rect 376706 522098 376942 522334
rect 377026 522098 377262 522334
rect 376706 521778 376942 522014
rect 377026 521778 377262 522014
rect 376706 486098 376942 486334
rect 377026 486098 377262 486334
rect 376706 485778 376942 486014
rect 377026 485778 377262 486014
rect 376706 450098 376942 450334
rect 377026 450098 377262 450334
rect 376706 449778 376942 450014
rect 377026 449778 377262 450014
rect 376706 414098 376942 414334
rect 377026 414098 377262 414334
rect 376706 413778 376942 414014
rect 377026 413778 377262 414014
rect 376706 378098 376942 378334
rect 377026 378098 377262 378334
rect 376706 377778 376942 378014
rect 377026 377778 377262 378014
rect 376706 342098 376942 342334
rect 377026 342098 377262 342334
rect 376706 341778 376942 342014
rect 377026 341778 377262 342014
rect 376706 306098 376942 306334
rect 377026 306098 377262 306334
rect 376706 305778 376942 306014
rect 377026 305778 377262 306014
rect 376706 270098 376942 270334
rect 377026 270098 377262 270334
rect 376706 269778 376942 270014
rect 377026 269778 377262 270014
rect 376706 234098 376942 234334
rect 377026 234098 377262 234334
rect 376706 233778 376942 234014
rect 377026 233778 377262 234014
rect 376706 198098 376942 198334
rect 377026 198098 377262 198334
rect 376706 197778 376942 198014
rect 377026 197778 377262 198014
rect 376706 162098 376942 162334
rect 377026 162098 377262 162334
rect 376706 161778 376942 162014
rect 377026 161778 377262 162014
rect 376706 126098 376942 126334
rect 377026 126098 377262 126334
rect 376706 125778 376942 126014
rect 377026 125778 377262 126014
rect 376706 90098 376942 90334
rect 377026 90098 377262 90334
rect 376706 89778 376942 90014
rect 377026 89778 377262 90014
rect 376706 54098 376942 54334
rect 377026 54098 377262 54334
rect 376706 53778 376942 54014
rect 377026 53778 377262 54014
rect 376706 18098 376942 18334
rect 377026 18098 377262 18334
rect 376706 17778 376942 18014
rect 377026 17778 377262 18014
rect 376706 -4422 376942 -4186
rect 377026 -4422 377262 -4186
rect 376706 -4742 376942 -4506
rect 377026 -4742 377262 -4506
rect 380426 709402 380662 709638
rect 380746 709402 380982 709638
rect 380426 709082 380662 709318
rect 380746 709082 380982 709318
rect 380426 669818 380662 670054
rect 380746 669818 380982 670054
rect 380426 669498 380662 669734
rect 380746 669498 380982 669734
rect 380426 633818 380662 634054
rect 380746 633818 380982 634054
rect 380426 633498 380662 633734
rect 380746 633498 380982 633734
rect 380426 597818 380662 598054
rect 380746 597818 380982 598054
rect 380426 597498 380662 597734
rect 380746 597498 380982 597734
rect 380426 561818 380662 562054
rect 380746 561818 380982 562054
rect 380426 561498 380662 561734
rect 380746 561498 380982 561734
rect 380426 525818 380662 526054
rect 380746 525818 380982 526054
rect 380426 525498 380662 525734
rect 380746 525498 380982 525734
rect 380426 489818 380662 490054
rect 380746 489818 380982 490054
rect 380426 489498 380662 489734
rect 380746 489498 380982 489734
rect 380426 453818 380662 454054
rect 380746 453818 380982 454054
rect 380426 453498 380662 453734
rect 380746 453498 380982 453734
rect 380426 417818 380662 418054
rect 380746 417818 380982 418054
rect 380426 417498 380662 417734
rect 380746 417498 380982 417734
rect 380426 381818 380662 382054
rect 380746 381818 380982 382054
rect 380426 381498 380662 381734
rect 380746 381498 380982 381734
rect 380426 345818 380662 346054
rect 380746 345818 380982 346054
rect 380426 345498 380662 345734
rect 380746 345498 380982 345734
rect 380426 309818 380662 310054
rect 380746 309818 380982 310054
rect 380426 309498 380662 309734
rect 380746 309498 380982 309734
rect 380426 273818 380662 274054
rect 380746 273818 380982 274054
rect 380426 273498 380662 273734
rect 380746 273498 380982 273734
rect 380426 237818 380662 238054
rect 380746 237818 380982 238054
rect 380426 237498 380662 237734
rect 380746 237498 380982 237734
rect 380426 201818 380662 202054
rect 380746 201818 380982 202054
rect 380426 201498 380662 201734
rect 380746 201498 380982 201734
rect 380426 165818 380662 166054
rect 380746 165818 380982 166054
rect 380426 165498 380662 165734
rect 380746 165498 380982 165734
rect 380426 129818 380662 130054
rect 380746 129818 380982 130054
rect 380426 129498 380662 129734
rect 380746 129498 380982 129734
rect 380426 93818 380662 94054
rect 380746 93818 380982 94054
rect 380426 93498 380662 93734
rect 380746 93498 380982 93734
rect 380426 57818 380662 58054
rect 380746 57818 380982 58054
rect 380426 57498 380662 57734
rect 380746 57498 380982 57734
rect 380426 21818 380662 22054
rect 380746 21818 380982 22054
rect 380426 21498 380662 21734
rect 380746 21498 380982 21734
rect 380426 -5382 380662 -5146
rect 380746 -5382 380982 -5146
rect 380426 -5702 380662 -5466
rect 380746 -5702 380982 -5466
rect 384146 710362 384382 710598
rect 384466 710362 384702 710598
rect 384146 710042 384382 710278
rect 384466 710042 384702 710278
rect 384146 673538 384382 673774
rect 384466 673538 384702 673774
rect 384146 673218 384382 673454
rect 384466 673218 384702 673454
rect 384146 637538 384382 637774
rect 384466 637538 384702 637774
rect 384146 637218 384382 637454
rect 384466 637218 384702 637454
rect 384146 601538 384382 601774
rect 384466 601538 384702 601774
rect 384146 601218 384382 601454
rect 384466 601218 384702 601454
rect 384146 565538 384382 565774
rect 384466 565538 384702 565774
rect 384146 565218 384382 565454
rect 384466 565218 384702 565454
rect 384146 529538 384382 529774
rect 384466 529538 384702 529774
rect 384146 529218 384382 529454
rect 384466 529218 384702 529454
rect 384146 493538 384382 493774
rect 384466 493538 384702 493774
rect 384146 493218 384382 493454
rect 384466 493218 384702 493454
rect 384146 457538 384382 457774
rect 384466 457538 384702 457774
rect 384146 457218 384382 457454
rect 384466 457218 384702 457454
rect 384146 421538 384382 421774
rect 384466 421538 384702 421774
rect 384146 421218 384382 421454
rect 384466 421218 384702 421454
rect 384146 385538 384382 385774
rect 384466 385538 384702 385774
rect 384146 385218 384382 385454
rect 384466 385218 384702 385454
rect 384146 349538 384382 349774
rect 384466 349538 384702 349774
rect 384146 349218 384382 349454
rect 384466 349218 384702 349454
rect 384146 313538 384382 313774
rect 384466 313538 384702 313774
rect 384146 313218 384382 313454
rect 384466 313218 384702 313454
rect 384146 277538 384382 277774
rect 384466 277538 384702 277774
rect 384146 277218 384382 277454
rect 384466 277218 384702 277454
rect 384146 241538 384382 241774
rect 384466 241538 384702 241774
rect 384146 241218 384382 241454
rect 384466 241218 384702 241454
rect 384146 205538 384382 205774
rect 384466 205538 384702 205774
rect 384146 205218 384382 205454
rect 384466 205218 384702 205454
rect 384146 169538 384382 169774
rect 384466 169538 384702 169774
rect 384146 169218 384382 169454
rect 384466 169218 384702 169454
rect 384146 133538 384382 133774
rect 384466 133538 384702 133774
rect 384146 133218 384382 133454
rect 384466 133218 384702 133454
rect 384146 97538 384382 97774
rect 384466 97538 384702 97774
rect 384146 97218 384382 97454
rect 384466 97218 384702 97454
rect 387866 711322 388102 711558
rect 388186 711322 388422 711558
rect 387866 711002 388102 711238
rect 388186 711002 388422 711238
rect 387866 677258 388102 677494
rect 388186 677258 388422 677494
rect 387866 676938 388102 677174
rect 388186 676938 388422 677174
rect 387866 641258 388102 641494
rect 388186 641258 388422 641494
rect 387866 640938 388102 641174
rect 388186 640938 388422 641174
rect 387866 605258 388102 605494
rect 388186 605258 388422 605494
rect 387866 604938 388102 605174
rect 388186 604938 388422 605174
rect 387866 569258 388102 569494
rect 388186 569258 388422 569494
rect 387866 568938 388102 569174
rect 388186 568938 388422 569174
rect 387866 533258 388102 533494
rect 388186 533258 388422 533494
rect 387866 532938 388102 533174
rect 388186 532938 388422 533174
rect 387866 497258 388102 497494
rect 388186 497258 388422 497494
rect 387866 496938 388102 497174
rect 388186 496938 388422 497174
rect 387866 461258 388102 461494
rect 388186 461258 388422 461494
rect 387866 460938 388102 461174
rect 388186 460938 388422 461174
rect 387866 425258 388102 425494
rect 388186 425258 388422 425494
rect 387866 424938 388102 425174
rect 388186 424938 388422 425174
rect 387866 389258 388102 389494
rect 388186 389258 388422 389494
rect 387866 388938 388102 389174
rect 388186 388938 388422 389174
rect 387866 353258 388102 353494
rect 388186 353258 388422 353494
rect 387866 352938 388102 353174
rect 388186 352938 388422 353174
rect 387866 317258 388102 317494
rect 388186 317258 388422 317494
rect 387866 316938 388102 317174
rect 388186 316938 388422 317174
rect 387866 281258 388102 281494
rect 388186 281258 388422 281494
rect 387866 280938 388102 281174
rect 388186 280938 388422 281174
rect 387866 245258 388102 245494
rect 388186 245258 388422 245494
rect 387866 244938 388102 245174
rect 388186 244938 388422 245174
rect 387866 209258 388102 209494
rect 388186 209258 388422 209494
rect 387866 208938 388102 209174
rect 388186 208938 388422 209174
rect 387866 173258 388102 173494
rect 388186 173258 388422 173494
rect 387866 172938 388102 173174
rect 388186 172938 388422 173174
rect 387866 137258 388102 137494
rect 388186 137258 388422 137494
rect 387866 136938 388102 137174
rect 388186 136938 388422 137174
rect 387866 101258 388102 101494
rect 388186 101258 388422 101494
rect 387866 100938 388102 101174
rect 388186 100938 388422 101174
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 404459 327218 404695 327454
rect 404459 326898 404695 327134
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 407932 330938 408168 331174
rect 407932 330618 408168 330854
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 412706 708442 412942 708678
rect 413026 708442 413262 708678
rect 412706 708122 412942 708358
rect 413026 708122 413262 708358
rect 412706 666098 412942 666334
rect 413026 666098 413262 666334
rect 412706 665778 412942 666014
rect 413026 665778 413262 666014
rect 412706 630098 412942 630334
rect 413026 630098 413262 630334
rect 412706 629778 412942 630014
rect 413026 629778 413262 630014
rect 412706 594098 412942 594334
rect 413026 594098 413262 594334
rect 412706 593778 412942 594014
rect 413026 593778 413262 594014
rect 412706 558098 412942 558334
rect 413026 558098 413262 558334
rect 412706 557778 412942 558014
rect 413026 557778 413262 558014
rect 412706 522098 412942 522334
rect 413026 522098 413262 522334
rect 412706 521778 412942 522014
rect 413026 521778 413262 522014
rect 412706 486098 412942 486334
rect 413026 486098 413262 486334
rect 412706 485778 412942 486014
rect 413026 485778 413262 486014
rect 412706 450098 412942 450334
rect 413026 450098 413262 450334
rect 412706 449778 412942 450014
rect 413026 449778 413262 450014
rect 412706 414098 412942 414334
rect 413026 414098 413262 414334
rect 412706 413778 412942 414014
rect 413026 413778 413262 414014
rect 412706 378098 412942 378334
rect 413026 378098 413262 378334
rect 412706 377778 412942 378014
rect 413026 377778 413262 378014
rect 412706 342098 412942 342334
rect 413026 342098 413262 342334
rect 412706 341778 412942 342014
rect 413026 341778 413262 342014
rect 411405 327218 411641 327454
rect 411405 326898 411641 327134
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 416426 709402 416662 709638
rect 416746 709402 416982 709638
rect 416426 709082 416662 709318
rect 416746 709082 416982 709318
rect 416426 669818 416662 670054
rect 416746 669818 416982 670054
rect 416426 669498 416662 669734
rect 416746 669498 416982 669734
rect 416426 633818 416662 634054
rect 416746 633818 416982 634054
rect 416426 633498 416662 633734
rect 416746 633498 416982 633734
rect 416426 597818 416662 598054
rect 416746 597818 416982 598054
rect 416426 597498 416662 597734
rect 416746 597498 416982 597734
rect 416426 561818 416662 562054
rect 416746 561818 416982 562054
rect 416426 561498 416662 561734
rect 416746 561498 416982 561734
rect 416426 525818 416662 526054
rect 416746 525818 416982 526054
rect 416426 525498 416662 525734
rect 416746 525498 416982 525734
rect 416426 489818 416662 490054
rect 416746 489818 416982 490054
rect 416426 489498 416662 489734
rect 416746 489498 416982 489734
rect 416426 453818 416662 454054
rect 416746 453818 416982 454054
rect 416426 453498 416662 453734
rect 416746 453498 416982 453734
rect 416426 417818 416662 418054
rect 416746 417818 416982 418054
rect 416426 417498 416662 417734
rect 416746 417498 416982 417734
rect 416426 381818 416662 382054
rect 416746 381818 416982 382054
rect 416426 381498 416662 381734
rect 416746 381498 416982 381734
rect 416426 345818 416662 346054
rect 416746 345818 416982 346054
rect 416426 345498 416662 345734
rect 416746 345498 416982 345734
rect 414878 330938 415114 331174
rect 414878 330618 415114 330854
rect 412706 306098 412942 306334
rect 413026 306098 413262 306334
rect 412706 305778 412942 306014
rect 413026 305778 413262 306014
rect 412706 270098 412942 270334
rect 413026 270098 413262 270334
rect 412706 269778 412942 270014
rect 413026 269778 413262 270014
rect 412706 234098 412942 234334
rect 413026 234098 413262 234334
rect 412706 233778 412942 234014
rect 413026 233778 413262 234014
rect 412706 198098 412942 198334
rect 413026 198098 413262 198334
rect 412706 197778 412942 198014
rect 413026 197778 413262 198014
rect 412706 162098 412942 162334
rect 413026 162098 413262 162334
rect 412706 161778 412942 162014
rect 413026 161778 413262 162014
rect 420146 710362 420382 710598
rect 420466 710362 420702 710598
rect 420146 710042 420382 710278
rect 420466 710042 420702 710278
rect 420146 673538 420382 673774
rect 420466 673538 420702 673774
rect 420146 673218 420382 673454
rect 420466 673218 420702 673454
rect 420146 637538 420382 637774
rect 420466 637538 420702 637774
rect 420146 637218 420382 637454
rect 420466 637218 420702 637454
rect 420146 601538 420382 601774
rect 420466 601538 420702 601774
rect 420146 601218 420382 601454
rect 420466 601218 420702 601454
rect 420146 565538 420382 565774
rect 420466 565538 420702 565774
rect 420146 565218 420382 565454
rect 420466 565218 420702 565454
rect 420146 529538 420382 529774
rect 420466 529538 420702 529774
rect 420146 529218 420382 529454
rect 420466 529218 420702 529454
rect 420146 493538 420382 493774
rect 420466 493538 420702 493774
rect 420146 493218 420382 493454
rect 420466 493218 420702 493454
rect 420146 457538 420382 457774
rect 420466 457538 420702 457774
rect 420146 457218 420382 457454
rect 420466 457218 420702 457454
rect 423866 711322 424102 711558
rect 424186 711322 424422 711558
rect 423866 711002 424102 711238
rect 424186 711002 424422 711238
rect 423866 677258 424102 677494
rect 424186 677258 424422 677494
rect 423866 676938 424102 677174
rect 424186 676938 424422 677174
rect 423866 641258 424102 641494
rect 424186 641258 424422 641494
rect 423866 640938 424102 641174
rect 424186 640938 424422 641174
rect 423866 605258 424102 605494
rect 424186 605258 424422 605494
rect 423866 604938 424102 605174
rect 424186 604938 424422 605174
rect 423866 569258 424102 569494
rect 424186 569258 424422 569494
rect 423866 568938 424102 569174
rect 424186 568938 424422 569174
rect 423866 533258 424102 533494
rect 424186 533258 424422 533494
rect 423866 532938 424102 533174
rect 424186 532938 424422 533174
rect 423866 497258 424102 497494
rect 424186 497258 424422 497494
rect 423866 496938 424102 497174
rect 424186 496938 424422 497174
rect 423866 461258 424102 461494
rect 424186 461258 424422 461494
rect 423866 460938 424102 461174
rect 424186 460938 424422 461174
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 426666 438938 426902 439174
rect 426666 438618 426902 438854
rect 432347 438938 432583 439174
rect 432347 438618 432583 438854
rect 438028 438938 438264 439174
rect 438028 438618 438264 438854
rect 443709 438938 443945 439174
rect 443709 438618 443945 438854
rect 423826 435218 424062 435454
rect 423826 434898 424062 435134
rect 429507 435218 429743 435454
rect 429507 434898 429743 435134
rect 435188 435218 435424 435454
rect 435188 434898 435424 435134
rect 440869 435218 441105 435454
rect 440869 434898 441105 435134
rect 420146 421538 420382 421774
rect 420466 421538 420702 421774
rect 420146 421218 420382 421454
rect 420466 421218 420702 421454
rect 420146 385538 420382 385774
rect 420466 385538 420702 385774
rect 420146 385218 420382 385454
rect 420466 385218 420702 385454
rect 420146 349538 420382 349774
rect 420466 349538 420702 349774
rect 420146 349218 420382 349454
rect 420466 349218 420702 349454
rect 418351 327218 418587 327454
rect 418351 326898 418587 327134
rect 416426 309818 416662 310054
rect 416746 309818 416982 310054
rect 416426 309498 416662 309734
rect 416746 309498 416982 309734
rect 416426 273818 416662 274054
rect 416746 273818 416982 274054
rect 416426 273498 416662 273734
rect 416746 273498 416982 273734
rect 416426 237818 416662 238054
rect 416746 237818 416982 238054
rect 416426 237498 416662 237734
rect 416746 237498 416982 237734
rect 416426 201818 416662 202054
rect 416746 201818 416982 202054
rect 416426 201498 416662 201734
rect 416746 201498 416982 201734
rect 416426 165818 416662 166054
rect 416746 165818 416982 166054
rect 416426 165498 416662 165734
rect 416746 165498 416982 165734
rect 423866 389258 424102 389494
rect 424186 389258 424422 389494
rect 423866 388938 424102 389174
rect 424186 388938 424422 389174
rect 423866 353258 424102 353494
rect 424186 353258 424422 353494
rect 423866 352938 424102 353174
rect 424186 352938 424422 353174
rect 420146 313538 420382 313774
rect 420466 313538 420702 313774
rect 420146 313218 420382 313454
rect 420466 313218 420702 313454
rect 420146 277538 420382 277774
rect 420466 277538 420702 277774
rect 420146 277218 420382 277454
rect 420466 277218 420702 277454
rect 420146 241538 420382 241774
rect 420466 241538 420702 241774
rect 420146 241218 420382 241454
rect 420466 241218 420702 241454
rect 420146 205538 420382 205774
rect 420466 205538 420702 205774
rect 420146 205218 420382 205454
rect 420466 205218 420702 205454
rect 420146 169538 420382 169774
rect 420466 169538 420702 169774
rect 420146 169218 420382 169454
rect 420466 169218 420702 169454
rect 421824 330938 422060 331174
rect 421824 330618 422060 330854
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 425297 327218 425533 327454
rect 425297 326898 425533 327134
rect 423866 317258 424102 317494
rect 424186 317258 424422 317494
rect 423866 316938 424102 317174
rect 424186 316938 424422 317174
rect 423866 281258 424102 281494
rect 424186 281258 424422 281494
rect 423866 280938 424102 281174
rect 424186 280938 424422 281174
rect 423866 245258 424102 245494
rect 424186 245258 424422 245494
rect 423866 244938 424102 245174
rect 424186 244938 424422 245174
rect 423866 209258 424102 209494
rect 424186 209258 424422 209494
rect 423866 208938 424102 209174
rect 424186 208938 424422 209174
rect 423866 173258 424102 173494
rect 424186 173258 424422 173494
rect 423866 172938 424102 173174
rect 424186 172938 424422 173174
rect 428770 330938 429006 331174
rect 428770 330618 429006 330854
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 448706 708442 448942 708678
rect 449026 708442 449262 708678
rect 448706 708122 448942 708358
rect 449026 708122 449262 708358
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 452426 709402 452662 709638
rect 452746 709402 452982 709638
rect 452426 709082 452662 709318
rect 452746 709082 452982 709318
rect 448706 666098 448942 666334
rect 449026 666098 449262 666334
rect 448706 665778 448942 666014
rect 449026 665778 449262 666014
rect 448706 630098 448942 630334
rect 449026 630098 449262 630334
rect 448706 629778 448942 630014
rect 449026 629778 449262 630014
rect 448706 594098 448942 594334
rect 449026 594098 449262 594334
rect 448706 593778 448942 594014
rect 449026 593778 449262 594014
rect 448706 558098 448942 558334
rect 449026 558098 449262 558334
rect 448706 557778 448942 558014
rect 449026 557778 449262 558014
rect 448706 522098 448942 522334
rect 449026 522098 449262 522334
rect 448706 521778 448942 522014
rect 449026 521778 449262 522014
rect 448706 486098 448942 486334
rect 449026 486098 449262 486334
rect 448706 485778 448942 486014
rect 449026 485778 449262 486014
rect 448706 450098 448942 450334
rect 449026 450098 449262 450334
rect 448706 449778 448942 450014
rect 449026 449778 449262 450014
rect 448706 414098 448942 414334
rect 449026 414098 449262 414334
rect 448706 413778 448942 414014
rect 449026 413778 449262 414014
rect 448706 378098 448942 378334
rect 449026 378098 449262 378334
rect 448706 377778 448942 378014
rect 449026 377778 449262 378014
rect 448706 342098 448942 342334
rect 449026 342098 449262 342334
rect 448706 341778 448942 342014
rect 449026 341778 449262 342014
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 452426 669818 452662 670054
rect 452746 669818 452982 670054
rect 452426 669498 452662 669734
rect 452746 669498 452982 669734
rect 452426 633818 452662 634054
rect 452746 633818 452982 634054
rect 452426 633498 452662 633734
rect 452746 633498 452982 633734
rect 452426 597818 452662 598054
rect 452746 597818 452982 598054
rect 452426 597498 452662 597734
rect 452746 597498 452982 597734
rect 452426 561818 452662 562054
rect 452746 561818 452982 562054
rect 452426 561498 452662 561734
rect 452746 561498 452982 561734
rect 452426 525818 452662 526054
rect 452746 525818 452982 526054
rect 452426 525498 452662 525734
rect 452746 525498 452982 525734
rect 456146 710362 456382 710598
rect 456466 710362 456702 710598
rect 456146 710042 456382 710278
rect 456466 710042 456702 710278
rect 456146 673538 456382 673774
rect 456466 673538 456702 673774
rect 456146 673218 456382 673454
rect 456466 673218 456702 673454
rect 459866 711322 460102 711558
rect 460186 711322 460422 711558
rect 459866 711002 460102 711238
rect 460186 711002 460422 711238
rect 459866 677258 460102 677494
rect 460186 677258 460422 677494
rect 459866 676938 460102 677174
rect 460186 676938 460422 677174
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 488426 709402 488662 709638
rect 488746 709402 488982 709638
rect 488426 709082 488662 709318
rect 488746 709082 488982 709318
rect 488426 669818 488662 670054
rect 488746 669818 488982 670054
rect 488426 669498 488662 669734
rect 488746 669498 488982 669734
rect 492146 710362 492382 710598
rect 492466 710362 492702 710598
rect 492146 710042 492382 710278
rect 492466 710042 492702 710278
rect 492146 673538 492382 673774
rect 492466 673538 492702 673774
rect 492146 673218 492382 673454
rect 492466 673218 492702 673454
rect 495866 711322 496102 711558
rect 496186 711322 496422 711558
rect 495866 711002 496102 711238
rect 496186 711002 496422 711238
rect 495866 677258 496102 677494
rect 496186 677258 496422 677494
rect 495866 676938 496102 677174
rect 496186 676938 496422 677174
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 520706 708442 520942 708678
rect 521026 708442 521262 708678
rect 520706 708122 520942 708358
rect 521026 708122 521262 708358
rect 520706 666098 520942 666334
rect 521026 666098 521262 666334
rect 520706 665778 520942 666014
rect 521026 665778 521262 666014
rect 456146 637538 456382 637774
rect 456466 637538 456702 637774
rect 456146 637218 456382 637454
rect 456466 637218 456702 637454
rect 456146 601538 456382 601774
rect 456466 601538 456702 601774
rect 456146 601218 456382 601454
rect 456466 601218 456702 601454
rect 456146 565538 456382 565774
rect 456466 565538 456702 565774
rect 456146 565218 456382 565454
rect 456466 565218 456702 565454
rect 456146 529538 456382 529774
rect 456466 529538 456702 529774
rect 456146 529218 456382 529454
rect 456466 529218 456702 529454
rect 453424 510938 453660 511174
rect 453424 510618 453660 510854
rect 455862 510938 456098 511174
rect 455862 510618 456098 510854
rect 458300 510938 458536 511174
rect 458300 510618 458536 510854
rect 452205 507218 452441 507454
rect 452205 506898 452441 507134
rect 454643 507218 454879 507454
rect 454643 506898 454879 507134
rect 457081 507218 457317 507454
rect 457081 506898 457317 507134
rect 452426 489818 452662 490054
rect 452746 489818 452982 490054
rect 452426 489498 452662 489734
rect 452746 489498 452982 489734
rect 452426 453818 452662 454054
rect 452746 453818 452982 454054
rect 452426 453498 452662 453734
rect 452746 453498 452982 453734
rect 452426 417818 452662 418054
rect 452746 417818 452982 418054
rect 452426 417498 452662 417734
rect 452746 417498 452982 417734
rect 452426 381818 452662 382054
rect 452746 381818 452982 382054
rect 452426 381498 452662 381734
rect 452746 381498 452982 381734
rect 456146 493538 456382 493774
rect 456466 493538 456702 493774
rect 456146 493218 456382 493454
rect 456466 493218 456702 493454
rect 456146 457538 456382 457774
rect 456466 457538 456702 457774
rect 456146 457218 456382 457454
rect 456466 457218 456702 457454
rect 479610 654938 479846 655174
rect 479610 654618 479846 654854
rect 510330 654938 510566 655174
rect 510330 654618 510566 654854
rect 464250 651218 464486 651454
rect 464250 650898 464486 651134
rect 494970 651218 495206 651454
rect 494970 650898 495206 651134
rect 520706 630098 520942 630334
rect 521026 630098 521262 630334
rect 520706 629778 520942 630014
rect 521026 629778 521262 630014
rect 479610 618938 479846 619174
rect 479610 618618 479846 618854
rect 510330 618938 510566 619174
rect 510330 618618 510566 618854
rect 464250 615218 464486 615454
rect 464250 614898 464486 615134
rect 494970 615218 495206 615454
rect 494970 614898 495206 615134
rect 459866 569258 460102 569494
rect 460186 569258 460422 569494
rect 459866 568938 460102 569174
rect 460186 568938 460422 569174
rect 459866 533258 460102 533494
rect 460186 533258 460422 533494
rect 459866 532938 460102 533174
rect 460186 532938 460422 533174
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 460738 510938 460974 511174
rect 460738 510618 460974 510854
rect 459519 507218 459755 507454
rect 459519 506898 459755 507134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 459866 497258 460102 497494
rect 460186 497258 460422 497494
rect 459866 496938 460102 497174
rect 460186 496938 460422 497174
rect 459866 461258 460102 461494
rect 460186 461258 460422 461494
rect 459866 460938 460102 461174
rect 460186 460938 460422 461174
rect 456146 421538 456382 421774
rect 456466 421538 456702 421774
rect 456146 421218 456382 421454
rect 456466 421218 456702 421454
rect 456146 385538 456382 385774
rect 456466 385538 456702 385774
rect 456146 385218 456382 385454
rect 456466 385218 456702 385454
rect 454250 363218 454486 363454
rect 454250 362898 454486 363134
rect 452426 345818 452662 346054
rect 452746 345818 452982 346054
rect 452426 345498 452662 345734
rect 452746 345498 452982 345734
rect 448706 306098 448942 306334
rect 449026 306098 449262 306334
rect 448706 305778 448942 306014
rect 449026 305778 449262 306014
rect 448706 270098 448942 270334
rect 449026 270098 449262 270334
rect 448706 269778 448942 270014
rect 449026 269778 449262 270014
rect 448706 234098 448942 234334
rect 449026 234098 449262 234334
rect 448706 233778 448942 234014
rect 449026 233778 449262 234014
rect 448706 198098 448942 198334
rect 449026 198098 449262 198334
rect 448706 197778 448942 198014
rect 449026 197778 449262 198014
rect 448706 162098 448942 162334
rect 449026 162098 449262 162334
rect 448706 161778 448942 162014
rect 449026 161778 449262 162014
rect 429610 150938 429846 151174
rect 429610 150618 429846 150854
rect 414250 147218 414486 147454
rect 414250 146898 414486 147134
rect 444970 147218 445206 147454
rect 444970 146898 445206 147134
rect 412706 126098 412942 126334
rect 413026 126098 413262 126334
rect 412706 125778 412942 126014
rect 413026 125778 413262 126014
rect 416426 93818 416662 94054
rect 416746 93818 416982 94054
rect 416426 93498 416662 93734
rect 416746 93498 416982 93734
rect 420146 97538 420382 97774
rect 420466 97538 420702 97774
rect 420146 97218 420382 97454
rect 420466 97218 420702 97454
rect 423866 101258 424102 101494
rect 424186 101258 424422 101494
rect 423866 100938 424102 101174
rect 424186 100938 424422 101174
rect 448706 126098 448942 126334
rect 449026 126098 449262 126334
rect 448706 125778 448942 126014
rect 449026 125778 449262 126014
rect 456146 349538 456382 349774
rect 456466 349538 456702 349774
rect 456146 349218 456382 349454
rect 456466 349218 456702 349454
rect 454250 327218 454486 327454
rect 454250 326898 454486 327134
rect 452426 309818 452662 310054
rect 452746 309818 452982 310054
rect 452426 309498 452662 309734
rect 452746 309498 452982 309734
rect 452426 273818 452662 274054
rect 452746 273818 452982 274054
rect 452426 273498 452662 273734
rect 452746 273498 452982 273734
rect 452426 237818 452662 238054
rect 452746 237818 452982 238054
rect 452426 237498 452662 237734
rect 452746 237498 452982 237734
rect 452426 201818 452662 202054
rect 452746 201818 452982 202054
rect 452426 201498 452662 201734
rect 452746 201498 452982 201734
rect 452426 165818 452662 166054
rect 452746 165818 452982 166054
rect 452426 165498 452662 165734
rect 452746 165498 452982 165734
rect 452426 129818 452662 130054
rect 452746 129818 452982 130054
rect 452426 129498 452662 129734
rect 452746 129498 452982 129734
rect 452426 93818 452662 94054
rect 452746 93818 452982 94054
rect 452426 93498 452662 93734
rect 452746 93498 452982 93734
rect 456146 313538 456382 313774
rect 456466 313538 456702 313774
rect 456146 313218 456382 313454
rect 456466 313218 456702 313454
rect 456146 277538 456382 277774
rect 456466 277538 456702 277774
rect 456146 277218 456382 277454
rect 456466 277218 456702 277454
rect 456146 241538 456382 241774
rect 456466 241538 456702 241774
rect 456146 241218 456382 241454
rect 456466 241218 456702 241454
rect 456146 205538 456382 205774
rect 456466 205538 456702 205774
rect 456146 205218 456382 205454
rect 456466 205218 456702 205454
rect 456146 169538 456382 169774
rect 456466 169538 456702 169774
rect 456146 169218 456382 169454
rect 456466 169218 456702 169454
rect 456146 133538 456382 133774
rect 456466 133538 456702 133774
rect 456146 133218 456382 133454
rect 456466 133218 456702 133454
rect 456146 97538 456382 97774
rect 456466 97538 456702 97774
rect 456146 97218 456382 97454
rect 456466 97218 456702 97454
rect 459866 425258 460102 425494
rect 460186 425258 460422 425494
rect 459866 424938 460102 425174
rect 460186 424938 460422 425174
rect 459866 389258 460102 389494
rect 460186 389258 460422 389494
rect 459866 388938 460102 389174
rect 460186 388938 460422 389174
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473458 435218 473694 435454
rect 473458 434898 473694 435134
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 475930 438938 476166 439174
rect 475930 438618 476166 438854
rect 478403 435218 478639 435454
rect 478403 434898 478639 435134
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 484706 594098 484942 594334
rect 485026 594098 485262 594334
rect 484706 593778 484942 594014
rect 485026 593778 485262 594014
rect 484706 558098 484942 558334
rect 485026 558098 485262 558334
rect 484706 557778 484942 558014
rect 485026 557778 485262 558014
rect 484706 522098 484942 522334
rect 485026 522098 485262 522334
rect 484706 521778 484942 522014
rect 485026 521778 485262 522014
rect 488426 597818 488662 598054
rect 488746 597818 488982 598054
rect 488426 597498 488662 597734
rect 488746 597498 488982 597734
rect 488426 561818 488662 562054
rect 488746 561818 488982 562054
rect 488426 561498 488662 561734
rect 488746 561498 488982 561734
rect 488426 525818 488662 526054
rect 488746 525818 488982 526054
rect 488426 525498 488662 525734
rect 488746 525498 488982 525734
rect 492146 565538 492382 565774
rect 492466 565538 492702 565774
rect 492146 565218 492382 565454
rect 492466 565218 492702 565454
rect 492146 529538 492382 529774
rect 492466 529538 492702 529774
rect 492146 529218 492382 529454
rect 492466 529218 492702 529454
rect 482205 507218 482441 507454
rect 482205 506898 482441 507134
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 483424 510938 483660 511174
rect 483424 510618 483660 510854
rect 485862 510938 486098 511174
rect 485862 510618 486098 510854
rect 488300 510938 488536 511174
rect 488300 510618 488536 510854
rect 490738 510938 490974 511174
rect 490738 510618 490974 510854
rect 484643 507218 484879 507454
rect 484643 506898 484879 507134
rect 487081 507218 487317 507454
rect 487081 506898 487317 507134
rect 489519 507218 489755 507454
rect 489519 506898 489755 507134
rect 484706 486098 484942 486334
rect 485026 486098 485262 486334
rect 484706 485778 484942 486014
rect 485026 485778 485262 486014
rect 488426 489818 488662 490054
rect 488746 489818 488982 490054
rect 488426 489498 488662 489734
rect 488746 489498 488982 489734
rect 488426 453771 488662 454007
rect 488746 453771 488982 454007
rect 484706 450098 484942 450334
rect 485026 450098 485262 450334
rect 484706 449778 484942 450014
rect 485026 449778 485262 450014
rect 480875 438938 481111 439174
rect 480875 438618 481111 438854
rect 483348 435218 483584 435454
rect 483348 434898 483584 435134
rect 485820 438938 486056 439174
rect 485820 438618 486056 438854
rect 488293 435218 488529 435454
rect 488293 434898 488529 435134
rect 484706 414098 484942 414334
rect 485026 414098 485262 414334
rect 484706 413778 484942 414014
rect 485026 413778 485262 414014
rect 492146 493538 492382 493774
rect 492466 493538 492702 493774
rect 492146 493218 492382 493454
rect 492466 493218 492702 493454
rect 492146 457538 492382 457774
rect 492466 457538 492702 457774
rect 492146 457218 492382 457454
rect 492466 457218 492702 457454
rect 490765 438938 491001 439174
rect 490765 438618 491001 438854
rect 492146 421538 492382 421774
rect 492466 421538 492702 421774
rect 492146 421218 492382 421454
rect 492466 421218 492702 421454
rect 495866 569258 496102 569494
rect 496186 569258 496422 569494
rect 495866 568938 496102 569174
rect 496186 568938 496422 569174
rect 495866 533258 496102 533494
rect 496186 533258 496422 533494
rect 495866 532938 496102 533174
rect 496186 532938 496422 533174
rect 495866 497258 496102 497494
rect 496186 497258 496422 497494
rect 495866 496938 496102 497174
rect 496186 496938 496422 497174
rect 495866 461258 496102 461494
rect 496186 461258 496422 461494
rect 495866 460938 496102 461174
rect 496186 460938 496422 461174
rect 495866 425258 496102 425494
rect 496186 425258 496422 425494
rect 495866 424938 496102 425174
rect 496186 424938 496422 425174
rect 495866 389258 496102 389494
rect 496186 389258 496422 389494
rect 495866 388938 496102 389174
rect 496186 388938 496422 389174
rect 469610 366938 469846 367174
rect 469610 366618 469846 366854
rect 484970 363218 485206 363454
rect 484970 362898 485206 363134
rect 459866 353258 460102 353494
rect 460186 353258 460422 353494
rect 459866 352938 460102 353174
rect 460186 352938 460422 353174
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 500330 366938 500566 367174
rect 500330 366618 500566 366854
rect 495866 353258 496102 353494
rect 496186 353258 496422 353494
rect 495866 352938 496102 353174
rect 496186 352938 496422 353174
rect 469610 330938 469846 331174
rect 469610 330618 469846 330854
rect 484970 327218 485206 327454
rect 484970 326898 485206 327134
rect 459866 317258 460102 317494
rect 460186 317258 460422 317494
rect 459866 316938 460102 317174
rect 460186 316938 460422 317174
rect 459866 281258 460102 281494
rect 460186 281258 460422 281494
rect 459866 280938 460102 281174
rect 460186 280938 460422 281174
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 484706 306098 484942 306334
rect 485026 306098 485262 306334
rect 484706 305778 484942 306014
rect 485026 305778 485262 306014
rect 484706 270098 484942 270334
rect 485026 270098 485262 270334
rect 484706 269778 484942 270014
rect 485026 269778 485262 270014
rect 488426 309818 488662 310054
rect 488746 309818 488982 310054
rect 488426 309498 488662 309734
rect 488746 309498 488982 309734
rect 488426 273818 488662 274054
rect 488746 273818 488982 274054
rect 488426 273498 488662 273734
rect 488746 273498 488982 273734
rect 492146 313538 492382 313774
rect 492466 313538 492702 313774
rect 492146 313218 492382 313454
rect 492466 313218 492702 313454
rect 492146 277538 492382 277774
rect 492466 277538 492702 277774
rect 492146 277218 492382 277454
rect 492466 277218 492702 277454
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 500330 330938 500566 331174
rect 500330 330618 500566 330854
rect 495866 317258 496102 317494
rect 496186 317258 496422 317494
rect 495866 316938 496102 317174
rect 496186 316938 496422 317174
rect 495866 281258 496102 281494
rect 496186 281258 496422 281494
rect 495866 280938 496102 281174
rect 496186 280938 496422 281174
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 520706 594098 520942 594334
rect 521026 594098 521262 594334
rect 520706 593778 520942 594014
rect 521026 593778 521262 594014
rect 520706 558098 520942 558334
rect 521026 558098 521262 558334
rect 520706 557778 520942 558014
rect 521026 557778 521262 558014
rect 520706 522098 520942 522334
rect 521026 522098 521262 522334
rect 520706 521778 520942 522014
rect 521026 521778 521262 522014
rect 520706 486098 520942 486334
rect 521026 486098 521262 486334
rect 520706 485778 520942 486014
rect 521026 485778 521262 486014
rect 520706 450098 520942 450334
rect 521026 450098 521262 450334
rect 520706 449778 520942 450014
rect 521026 449778 521262 450014
rect 520706 414098 520942 414334
rect 521026 414098 521262 414334
rect 520706 413778 520942 414014
rect 521026 413778 521262 414014
rect 520706 378098 520942 378334
rect 521026 378098 521262 378334
rect 520706 377778 520942 378014
rect 521026 377778 521262 378014
rect 520706 342098 520942 342334
rect 521026 342098 521262 342334
rect 520706 341778 520942 342014
rect 521026 341778 521262 342014
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 520706 306098 520942 306334
rect 521026 306098 521262 306334
rect 520706 305778 520942 306014
rect 521026 305778 521262 306014
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 520706 270098 520942 270334
rect 521026 270098 521262 270334
rect 520706 269778 520942 270014
rect 521026 269778 521262 270014
rect 524426 709402 524662 709638
rect 524746 709402 524982 709638
rect 524426 709082 524662 709318
rect 524746 709082 524982 709318
rect 528146 710362 528382 710598
rect 528466 710362 528702 710598
rect 528146 710042 528382 710278
rect 528466 710042 528702 710278
rect 524426 669818 524662 670054
rect 524746 669818 524982 670054
rect 524426 669498 524662 669734
rect 524746 669498 524982 669734
rect 525690 651218 525926 651454
rect 525690 650898 525926 651134
rect 524426 633818 524662 634054
rect 524746 633818 524982 634054
rect 524426 633498 524662 633734
rect 524746 633498 524982 633734
rect 525690 615218 525926 615454
rect 525690 614898 525926 615134
rect 524426 597818 524662 598054
rect 524746 597818 524982 598054
rect 524426 597498 524662 597734
rect 524746 597498 524982 597734
rect 524426 561818 524662 562054
rect 524746 561818 524982 562054
rect 524426 561498 524662 561734
rect 524746 561498 524982 561734
rect 524426 525818 524662 526054
rect 524746 525818 524982 526054
rect 524426 525498 524662 525734
rect 524746 525498 524982 525734
rect 524426 489818 524662 490054
rect 524746 489818 524982 490054
rect 524426 489498 524662 489734
rect 524746 489498 524982 489734
rect 524426 453818 524662 454054
rect 524746 453818 524982 454054
rect 524426 453498 524662 453734
rect 524746 453498 524982 453734
rect 525206 435218 525442 435454
rect 525206 434898 525442 435134
rect 524426 417818 524662 418054
rect 524746 417818 524982 418054
rect 524426 417498 524662 417734
rect 524746 417498 524982 417734
rect 524426 381818 524662 382054
rect 524746 381818 524982 382054
rect 524426 381498 524662 381734
rect 524746 381498 524982 381734
rect 524426 345818 524662 346054
rect 524746 345818 524982 346054
rect 524426 345498 524662 345734
rect 524746 345498 524982 345734
rect 531866 711322 532102 711558
rect 532186 711322 532422 711558
rect 531866 711002 532102 711238
rect 532186 711002 532422 711238
rect 528146 673538 528382 673774
rect 528466 673538 528702 673774
rect 528146 673218 528382 673454
rect 528466 673218 528702 673454
rect 528146 637538 528382 637774
rect 528466 637538 528702 637774
rect 528146 637218 528382 637454
rect 528466 637218 528702 637454
rect 528146 601538 528382 601774
rect 528466 601538 528702 601774
rect 528146 601218 528382 601454
rect 528466 601218 528702 601454
rect 528146 565538 528382 565774
rect 528466 565538 528702 565774
rect 528146 565218 528382 565454
rect 528466 565218 528702 565454
rect 528146 529538 528382 529774
rect 528466 529538 528702 529774
rect 528146 529218 528382 529454
rect 528466 529218 528702 529454
rect 528146 493538 528382 493774
rect 528466 493538 528702 493774
rect 528146 493218 528382 493454
rect 528466 493218 528702 493454
rect 528146 457538 528382 457774
rect 528466 457538 528702 457774
rect 528146 457218 528382 457454
rect 528466 457218 528702 457454
rect 529426 438938 529662 439174
rect 529426 438618 529662 438854
rect 528146 421538 528382 421774
rect 528466 421538 528702 421774
rect 528146 421218 528382 421454
rect 528466 421218 528702 421454
rect 528146 385538 528382 385774
rect 528466 385538 528702 385774
rect 528146 385218 528382 385454
rect 528466 385218 528702 385454
rect 528146 349538 528382 349774
rect 528466 349538 528702 349774
rect 528146 349218 528382 349454
rect 528466 349218 528702 349454
rect 524426 309818 524662 310054
rect 524746 309818 524982 310054
rect 524426 309498 524662 309734
rect 524746 309498 524982 309734
rect 524426 273818 524662 274054
rect 524746 273818 524982 274054
rect 524426 273498 524662 273734
rect 524746 273498 524982 273734
rect 531866 677258 532102 677494
rect 532186 677258 532422 677494
rect 531866 676938 532102 677174
rect 532186 676938 532422 677174
rect 531866 641258 532102 641494
rect 532186 641258 532422 641494
rect 531866 640938 532102 641174
rect 532186 640938 532422 641174
rect 531866 605258 532102 605494
rect 532186 605258 532422 605494
rect 531866 604938 532102 605174
rect 532186 604938 532422 605174
rect 531866 569258 532102 569494
rect 532186 569258 532422 569494
rect 531866 568938 532102 569174
rect 532186 568938 532422 569174
rect 531866 533258 532102 533494
rect 532186 533258 532422 533494
rect 531866 532938 532102 533174
rect 532186 532938 532422 533174
rect 531866 497258 532102 497494
rect 532186 497258 532422 497494
rect 531866 496938 532102 497174
rect 532186 496938 532422 497174
rect 531866 461258 532102 461494
rect 532186 461258 532422 461494
rect 531866 460938 532102 461174
rect 532186 460938 532422 461174
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 537867 438938 538103 439174
rect 537867 438618 538103 438854
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 533647 435218 533883 435454
rect 533647 434898 533883 435134
rect 542088 435218 542324 435454
rect 542088 434898 542324 435134
rect 531866 425258 532102 425494
rect 532186 425258 532422 425494
rect 531866 424938 532102 425174
rect 532186 424938 532422 425174
rect 531866 389258 532102 389494
rect 532186 389258 532422 389494
rect 531866 388938 532102 389174
rect 532186 388938 532422 389174
rect 531866 353258 532102 353494
rect 532186 353258 532422 353494
rect 531866 352938 532102 353174
rect 532186 352938 532422 353174
rect 528146 313538 528382 313774
rect 528466 313538 528702 313774
rect 528146 313218 528382 313454
rect 528466 313218 528702 313454
rect 528146 277538 528382 277774
rect 528466 277538 528702 277774
rect 528146 277218 528382 277454
rect 528466 277218 528702 277454
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 531866 317258 532102 317494
rect 532186 317258 532422 317494
rect 531866 316938 532102 317174
rect 532186 316938 532422 317174
rect 531866 281258 532102 281494
rect 532186 281258 532422 281494
rect 531866 280938 532102 281174
rect 532186 280938 532422 281174
rect 479610 258938 479846 259174
rect 479610 258618 479846 258854
rect 510330 258938 510566 259174
rect 510330 258618 510566 258854
rect 464250 255218 464486 255454
rect 464250 254898 464486 255134
rect 494970 255218 495206 255454
rect 494970 254898 495206 255134
rect 525690 255218 525926 255454
rect 525690 254898 525926 255134
rect 459866 245258 460102 245494
rect 460186 245258 460422 245494
rect 459866 244938 460102 245174
rect 460186 244938 460422 245174
rect 531866 245258 532102 245494
rect 532186 245258 532422 245494
rect 531866 244938 532102 245174
rect 532186 244938 532422 245174
rect 479610 222938 479846 223174
rect 479610 222618 479846 222854
rect 510330 222938 510566 223174
rect 510330 222618 510566 222854
rect 464250 219218 464486 219454
rect 464250 218898 464486 219134
rect 494970 219218 495206 219454
rect 494970 218898 495206 219134
rect 525690 219218 525926 219454
rect 525690 218898 525926 219134
rect 459866 209258 460102 209494
rect 460186 209258 460422 209494
rect 459866 208938 460102 209174
rect 460186 208938 460422 209174
rect 531866 209258 532102 209494
rect 532186 209258 532422 209494
rect 531866 208938 532102 209174
rect 532186 208938 532422 209174
rect 459866 173258 460102 173494
rect 460186 173258 460422 173494
rect 459866 172938 460102 173174
rect 460186 172938 460422 173174
rect 459866 137258 460102 137494
rect 460186 137258 460422 137494
rect 459866 136938 460102 137174
rect 460186 136938 460422 137174
rect 459866 101258 460102 101494
rect 460186 101258 460422 101494
rect 459866 100938 460102 101174
rect 460186 100938 460422 101174
rect 405610 78938 405846 79174
rect 405610 78618 405846 78854
rect 436330 78938 436566 79174
rect 436330 78618 436566 78854
rect 390250 75218 390486 75454
rect 390250 74898 390486 75134
rect 420970 75218 421206 75454
rect 420970 74898 421206 75134
rect 451690 75218 451926 75454
rect 451690 74898 451926 75134
rect 384146 61538 384382 61774
rect 384466 61538 384702 61774
rect 384146 61218 384382 61454
rect 384466 61218 384702 61454
rect 459866 65258 460102 65494
rect 460186 65258 460422 65494
rect 459866 64938 460102 65174
rect 460186 64938 460422 65174
rect 405610 42938 405846 43174
rect 405610 42618 405846 42854
rect 436330 42938 436566 43174
rect 436330 42618 436566 42854
rect 390250 39218 390486 39454
rect 390250 38898 390486 39134
rect 420970 39218 421206 39454
rect 420970 38898 421206 39134
rect 451690 39218 451926 39454
rect 451690 38898 451926 39134
rect 384146 25538 384382 25774
rect 384466 25538 384702 25774
rect 384146 25218 384382 25454
rect 384466 25218 384702 25454
rect 384146 -6342 384382 -6106
rect 384466 -6342 384702 -6106
rect 384146 -6662 384382 -6426
rect 384466 -6662 384702 -6426
rect 387866 29258 388102 29494
rect 388186 29258 388422 29494
rect 387866 28938 388102 29174
rect 388186 28938 388422 29174
rect 387866 -7302 388102 -7066
rect 388186 -7302 388422 -7066
rect 387866 -7622 388102 -7386
rect 388186 -7622 388422 -7386
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 408986 -3462 409222 -3226
rect 409306 -3462 409542 -3226
rect 408986 -3782 409222 -3546
rect 409306 -3782 409542 -3546
rect 412706 18098 412942 18334
rect 413026 18098 413262 18334
rect 412706 17778 412942 18014
rect 413026 17778 413262 18014
rect 412706 -4422 412942 -4186
rect 413026 -4422 413262 -4186
rect 412706 -4742 412942 -4506
rect 413026 -4742 413262 -4506
rect 416426 21818 416662 22054
rect 416746 21818 416982 22054
rect 416426 21498 416662 21734
rect 416746 21498 416982 21734
rect 416426 -5382 416662 -5146
rect 416746 -5382 416982 -5146
rect 416426 -5702 416662 -5466
rect 416746 -5702 416982 -5466
rect 420146 25538 420382 25774
rect 420466 25538 420702 25774
rect 420146 25218 420382 25454
rect 420466 25218 420702 25454
rect 420146 -6342 420382 -6106
rect 420466 -6342 420702 -6106
rect 420146 -6662 420382 -6426
rect 420466 -6662 420702 -6426
rect 423866 29258 424102 29494
rect 424186 29258 424422 29494
rect 423866 28938 424102 29174
rect 424186 28938 424422 29174
rect 423866 -7302 424102 -7066
rect 424186 -7302 424422 -7066
rect 423866 -7622 424102 -7386
rect 424186 -7622 424422 -7386
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 444986 -3462 445222 -3226
rect 445306 -3462 445542 -3226
rect 444986 -3782 445222 -3546
rect 445306 -3782 445542 -3546
rect 448706 18098 448942 18334
rect 449026 18098 449262 18334
rect 448706 17778 448942 18014
rect 449026 17778 449262 18014
rect 448706 -4422 448942 -4186
rect 449026 -4422 449262 -4186
rect 448706 -4742 448942 -4506
rect 449026 -4742 449262 -4506
rect 452426 21818 452662 22054
rect 452746 21818 452982 22054
rect 452426 21498 452662 21734
rect 452746 21498 452982 21734
rect 452426 -5382 452662 -5146
rect 452746 -5382 452982 -5146
rect 452426 -5702 452662 -5466
rect 452746 -5702 452982 -5466
rect 456146 25538 456382 25774
rect 456466 25538 456702 25774
rect 456146 25218 456382 25454
rect 456466 25218 456702 25454
rect 456146 -6342 456382 -6106
rect 456466 -6342 456702 -6106
rect 456146 -6662 456382 -6426
rect 456466 -6662 456702 -6426
rect 459866 29258 460102 29494
rect 460186 29258 460422 29494
rect 459866 28938 460102 29174
rect 460186 28938 460422 29174
rect 459866 -7302 460102 -7066
rect 460186 -7302 460422 -7066
rect 459866 -7622 460102 -7386
rect 460186 -7622 460422 -7386
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 484706 198098 484942 198334
rect 485026 198098 485262 198334
rect 484706 197778 484942 198014
rect 485026 197778 485262 198014
rect 484706 162098 484942 162334
rect 485026 162098 485262 162334
rect 484706 161778 484942 162014
rect 485026 161778 485262 162014
rect 488426 165818 488662 166054
rect 488746 165818 488982 166054
rect 488426 165498 488662 165734
rect 488746 165498 488982 165734
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 520706 198098 520942 198334
rect 521026 198098 521262 198334
rect 520706 197778 520942 198014
rect 521026 197778 521262 198014
rect 520706 162098 520942 162334
rect 521026 162098 521262 162334
rect 520706 161778 520942 162014
rect 521026 161778 521262 162014
rect 524426 165818 524662 166054
rect 524746 165818 524982 166054
rect 524426 165498 524662 165734
rect 524746 165498 524982 165734
rect 531866 173258 532102 173494
rect 532186 173258 532422 173494
rect 531866 172938 532102 173174
rect 532186 172938 532422 173174
rect 546308 438938 546544 439174
rect 546308 438618 546544 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 484706 126098 484942 126334
rect 485026 126098 485262 126334
rect 484706 125778 484942 126014
rect 485026 125778 485262 126014
rect 484250 111218 484486 111454
rect 484250 110898 484486 111134
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 480986 -3462 481222 -3226
rect 481306 -3462 481542 -3226
rect 480986 -3782 481222 -3546
rect 481306 -3782 481542 -3546
rect 499610 114938 499846 115174
rect 499610 114618 499846 114854
rect 530330 114938 530566 115174
rect 530330 114618 530566 114854
rect 514970 111218 515206 111454
rect 514970 110898 515206 111134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 484706 90098 484942 90334
rect 485026 90098 485262 90334
rect 484706 89778 484942 90014
rect 485026 89778 485262 90014
rect 484706 54098 484942 54334
rect 485026 54098 485262 54334
rect 484706 53778 484942 54014
rect 485026 53778 485262 54014
rect 484706 18098 484942 18334
rect 485026 18098 485262 18334
rect 484706 17778 484942 18014
rect 485026 17778 485262 18014
rect 484706 -4422 484942 -4186
rect 485026 -4422 485262 -4186
rect 484706 -4742 484942 -4506
rect 485026 -4742 485262 -4506
rect 488426 57818 488662 58054
rect 488746 57818 488982 58054
rect 488426 57498 488662 57734
rect 488746 57498 488982 57734
rect 488426 21818 488662 22054
rect 488746 21818 488982 22054
rect 488426 21498 488662 21734
rect 488746 21498 488982 21734
rect 488426 -5382 488662 -5146
rect 488746 -5382 488982 -5146
rect 488426 -5702 488662 -5466
rect 488746 -5702 488982 -5466
rect 492146 61538 492382 61774
rect 492466 61538 492702 61774
rect 492146 61218 492382 61454
rect 492466 61218 492702 61454
rect 492146 25538 492382 25774
rect 492466 25538 492702 25774
rect 492146 25218 492382 25454
rect 492466 25218 492702 25454
rect 492146 -6342 492382 -6106
rect 492466 -6342 492702 -6106
rect 492146 -6662 492382 -6426
rect 492466 -6662 492702 -6426
rect 495866 65258 496102 65494
rect 496186 65258 496422 65494
rect 495866 64938 496102 65174
rect 496186 64938 496422 65174
rect 495866 29258 496102 29494
rect 496186 29258 496422 29494
rect 495866 28938 496102 29174
rect 496186 28938 496422 29174
rect 495866 -7302 496102 -7066
rect 496186 -7302 496422 -7066
rect 495866 -7622 496102 -7386
rect 496186 -7622 496422 -7386
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 516986 -3462 517222 -3226
rect 517306 -3462 517542 -3226
rect 516986 -3782 517222 -3546
rect 517306 -3782 517542 -3546
rect 520706 54098 520942 54334
rect 521026 54098 521262 54334
rect 520706 53778 520942 54014
rect 521026 53778 521262 54014
rect 520706 18098 520942 18334
rect 521026 18098 521262 18334
rect 520706 17778 520942 18014
rect 521026 17778 521262 18014
rect 520706 -4422 520942 -4186
rect 521026 -4422 521262 -4186
rect 520706 -4742 520942 -4506
rect 521026 -4742 521262 -4506
rect 524426 57818 524662 58054
rect 524746 57818 524982 58054
rect 524426 57498 524662 57734
rect 524746 57498 524982 57734
rect 524426 21818 524662 22054
rect 524746 21818 524982 22054
rect 524426 21498 524662 21734
rect 524746 21498 524982 21734
rect 524426 -5382 524662 -5146
rect 524746 -5382 524982 -5146
rect 524426 -5702 524662 -5466
rect 524746 -5702 524982 -5466
rect 528146 61538 528382 61774
rect 528466 61538 528702 61774
rect 528146 61218 528382 61454
rect 528466 61218 528702 61454
rect 528146 25538 528382 25774
rect 528466 25538 528702 25774
rect 528146 25218 528382 25454
rect 528466 25218 528702 25454
rect 528146 -6342 528382 -6106
rect 528466 -6342 528702 -6106
rect 528146 -6662 528382 -6426
rect 528466 -6662 528702 -6426
rect 531866 65258 532102 65494
rect 532186 65258 532422 65494
rect 531866 64938 532102 65174
rect 532186 64938 532422 65174
rect 531866 29258 532102 29494
rect 532186 29258 532422 29494
rect 531866 28938 532102 29174
rect 532186 28938 532422 29174
rect 531866 -7302 532102 -7066
rect 532186 -7302 532422 -7066
rect 531866 -7622 532102 -7386
rect 532186 -7622 532422 -7386
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 550529 435218 550765 435454
rect 550529 434898 550765 435134
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 556706 708442 556942 708678
rect 557026 708442 557262 708678
rect 556706 708122 556942 708358
rect 557026 708122 557262 708358
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 556706 666098 556942 666334
rect 557026 666098 557262 666334
rect 556706 665778 556942 666014
rect 557026 665778 557262 666014
rect 556706 630098 556942 630334
rect 557026 630098 557262 630334
rect 556706 629778 556942 630014
rect 557026 629778 557262 630014
rect 556706 594098 556942 594334
rect 557026 594098 557262 594334
rect 556706 593778 556942 594014
rect 557026 593778 557262 594014
rect 556706 558098 556942 558334
rect 557026 558098 557262 558334
rect 556706 557778 556942 558014
rect 557026 557778 557262 558014
rect 556706 522098 556942 522334
rect 557026 522098 557262 522334
rect 556706 521778 556942 522014
rect 557026 521778 557262 522014
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 554749 438938 554985 439174
rect 554749 438618 554985 438854
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 556706 414098 556942 414334
rect 557026 414098 557262 414334
rect 556706 413778 556942 414014
rect 557026 413778 557262 414014
rect 556706 378007 556942 378243
rect 557026 378007 557262 378243
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 554918 366938 555154 367174
rect 554918 366618 555154 366854
rect 552952 363218 553188 363454
rect 552952 362898 553188 363134
rect 556885 363218 557121 363454
rect 556885 362898 557121 363134
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 556706 342098 556942 342334
rect 557026 342098 557262 342334
rect 556706 341778 556942 342014
rect 557026 341778 557262 342014
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 558851 366938 559087 367174
rect 558851 366618 559087 366854
rect 562784 366938 563020 367174
rect 562784 366618 563020 366854
rect 566717 366938 566953 367174
rect 566717 366618 566953 366854
rect 560818 363218 561054 363454
rect 560818 362898 561054 363134
rect 564751 363218 564987 363454
rect 564751 362898 564987 363134
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 556706 306098 556942 306334
rect 557026 306098 557262 306334
rect 556706 305778 556942 306014
rect 557026 305778 557262 306014
rect 556706 270098 556942 270334
rect 557026 270098 557262 270334
rect 556706 269778 556942 270014
rect 557026 269778 557262 270014
rect 556706 234098 556942 234334
rect 557026 234098 557262 234334
rect 556706 233778 556942 234014
rect 557026 233778 557262 234014
rect 556706 198098 556942 198334
rect 557026 198098 557262 198334
rect 556706 197778 556942 198014
rect 557026 197778 557262 198014
rect 556706 162098 556942 162334
rect 557026 162098 557262 162334
rect 556706 161778 556942 162014
rect 557026 161778 557262 162014
rect 556706 126098 556942 126334
rect 557026 126098 557262 126334
rect 556706 125778 556942 126014
rect 557026 125778 557262 126014
rect 556706 90098 556942 90334
rect 557026 90098 557262 90334
rect 556706 89778 556942 90014
rect 557026 89778 557262 90014
rect 556706 54098 556942 54334
rect 557026 54098 557262 54334
rect 556706 53778 556942 54014
rect 557026 53778 557262 54014
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 545930 42938 546166 43174
rect 545930 42618 546166 42854
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 543458 39218 543694 39454
rect 543458 38898 543694 39134
rect 548403 39218 548639 39454
rect 548403 38898 548639 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 550875 42938 551111 43174
rect 550875 42618 551111 42854
rect 555820 42938 556056 43174
rect 555820 42618 556056 42854
rect 553348 39218 553584 39454
rect 553348 38898 553584 39134
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 560765 42938 561001 43174
rect 560765 42618 561001 42854
rect 558293 39218 558529 39454
rect 558293 38898 558529 39134
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 39610 655174
rect 39846 654938 70330 655174
rect 70566 654938 101050 655174
rect 101286 654938 131770 655174
rect 132006 654938 162490 655174
rect 162726 654938 193210 655174
rect 193446 654938 223930 655174
rect 224166 654938 254650 655174
rect 254886 654938 285370 655174
rect 285606 654938 316090 655174
rect 316326 654938 346810 655174
rect 347046 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 479610 655174
rect 479846 654938 510330 655174
rect 510566 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 39610 654854
rect 39846 654618 70330 654854
rect 70566 654618 101050 654854
rect 101286 654618 131770 654854
rect 132006 654618 162490 654854
rect 162726 654618 193210 654854
rect 193446 654618 223930 654854
rect 224166 654618 254650 654854
rect 254886 654618 285370 654854
rect 285606 654618 316090 654854
rect 316326 654618 346810 654854
rect 347046 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 479610 654854
rect 479846 654618 510330 654854
rect 510566 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 24250 651454
rect 24486 651218 54970 651454
rect 55206 651218 85690 651454
rect 85926 651218 116410 651454
rect 116646 651218 147130 651454
rect 147366 651218 177850 651454
rect 178086 651218 208570 651454
rect 208806 651218 239290 651454
rect 239526 651218 270010 651454
rect 270246 651218 300730 651454
rect 300966 651218 331450 651454
rect 331686 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 464250 651454
rect 464486 651218 494970 651454
rect 495206 651218 525690 651454
rect 525926 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 24250 651134
rect 24486 650898 54970 651134
rect 55206 650898 85690 651134
rect 85926 650898 116410 651134
rect 116646 650898 147130 651134
rect 147366 650898 177850 651134
rect 178086 650898 208570 651134
rect 208806 650898 239290 651134
rect 239526 650898 270010 651134
rect 270246 650898 300730 651134
rect 300966 650898 331450 651134
rect 331686 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 464250 651134
rect 464486 650898 494970 651134
rect 495206 650898 525690 651134
rect 525926 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 520706 630334
rect 520942 630098 521026 630334
rect 521262 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 520706 630014
rect 520942 629778 521026 630014
rect 521262 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 39610 619174
rect 39846 618938 70330 619174
rect 70566 618938 101050 619174
rect 101286 618938 131770 619174
rect 132006 618938 162490 619174
rect 162726 618938 193210 619174
rect 193446 618938 223930 619174
rect 224166 618938 254650 619174
rect 254886 618938 285370 619174
rect 285606 618938 316090 619174
rect 316326 618938 346810 619174
rect 347046 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 479610 619174
rect 479846 618938 510330 619174
rect 510566 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 39610 618854
rect 39846 618618 70330 618854
rect 70566 618618 101050 618854
rect 101286 618618 131770 618854
rect 132006 618618 162490 618854
rect 162726 618618 193210 618854
rect 193446 618618 223930 618854
rect 224166 618618 254650 618854
rect 254886 618618 285370 618854
rect 285606 618618 316090 618854
rect 316326 618618 346810 618854
rect 347046 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 479610 618854
rect 479846 618618 510330 618854
rect 510566 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 24250 615454
rect 24486 615218 54970 615454
rect 55206 615218 85690 615454
rect 85926 615218 116410 615454
rect 116646 615218 147130 615454
rect 147366 615218 177850 615454
rect 178086 615218 208570 615454
rect 208806 615218 239290 615454
rect 239526 615218 270010 615454
rect 270246 615218 300730 615454
rect 300966 615218 331450 615454
rect 331686 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 464250 615454
rect 464486 615218 494970 615454
rect 495206 615218 525690 615454
rect 525926 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 24250 615134
rect 24486 614898 54970 615134
rect 55206 614898 85690 615134
rect 85926 614898 116410 615134
rect 116646 614898 147130 615134
rect 147366 614898 177850 615134
rect 178086 614898 208570 615134
rect 208806 614898 239290 615134
rect 239526 614898 270010 615134
rect 270246 614898 300730 615134
rect 300966 614898 331450 615134
rect 331686 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 464250 615134
rect 464486 614898 494970 615134
rect 495206 614898 525690 615134
rect 525926 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 39610 583174
rect 39846 582938 70330 583174
rect 70566 582938 101050 583174
rect 101286 582938 131770 583174
rect 132006 582938 162490 583174
rect 162726 582938 193210 583174
rect 193446 582938 223930 583174
rect 224166 582938 254650 583174
rect 254886 582938 285370 583174
rect 285606 582938 316090 583174
rect 316326 582938 346810 583174
rect 347046 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 39610 582854
rect 39846 582618 70330 582854
rect 70566 582618 101050 582854
rect 101286 582618 131770 582854
rect 132006 582618 162490 582854
rect 162726 582618 193210 582854
rect 193446 582618 223930 582854
rect 224166 582618 254650 582854
rect 254886 582618 285370 582854
rect 285606 582618 316090 582854
rect 316326 582618 346810 582854
rect 347046 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 24250 579454
rect 24486 579218 54970 579454
rect 55206 579218 85690 579454
rect 85926 579218 116410 579454
rect 116646 579218 147130 579454
rect 147366 579218 177850 579454
rect 178086 579218 208570 579454
rect 208806 579218 239290 579454
rect 239526 579218 270010 579454
rect 270246 579218 300730 579454
rect 300966 579218 331450 579454
rect 331686 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 24250 579134
rect 24486 578898 54970 579134
rect 55206 578898 85690 579134
rect 85926 578898 116410 579134
rect 116646 578898 147130 579134
rect 147366 578898 177850 579134
rect 178086 578898 208570 579134
rect 208806 578898 239290 579134
rect 239526 578898 270010 579134
rect 270246 578898 300730 579134
rect 300966 578898 331450 579134
rect 331686 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 39610 547174
rect 39846 546938 70330 547174
rect 70566 546938 101050 547174
rect 101286 546938 131770 547174
rect 132006 546938 162490 547174
rect 162726 546938 193210 547174
rect 193446 546938 223930 547174
rect 224166 546938 254650 547174
rect 254886 546938 285370 547174
rect 285606 546938 316090 547174
rect 316326 546938 346810 547174
rect 347046 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 39610 546854
rect 39846 546618 70330 546854
rect 70566 546618 101050 546854
rect 101286 546618 131770 546854
rect 132006 546618 162490 546854
rect 162726 546618 193210 546854
rect 193446 546618 223930 546854
rect 224166 546618 254650 546854
rect 254886 546618 285370 546854
rect 285606 546618 316090 546854
rect 316326 546618 346810 546854
rect 347046 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 24250 543454
rect 24486 543218 54970 543454
rect 55206 543218 85690 543454
rect 85926 543218 116410 543454
rect 116646 543218 147130 543454
rect 147366 543218 177850 543454
rect 178086 543218 208570 543454
rect 208806 543218 239290 543454
rect 239526 543218 270010 543454
rect 270246 543218 300730 543454
rect 300966 543218 331450 543454
rect 331686 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 24250 543134
rect 24486 542898 54970 543134
rect 55206 542898 85690 543134
rect 85926 542898 116410 543134
rect 116646 542898 147130 543134
rect 147366 542898 177850 543134
rect 178086 542898 208570 543134
rect 208806 542898 239290 543134
rect 239526 542898 270010 543134
rect 270246 542898 300730 543134
rect 300966 542898 331450 543134
rect 331686 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 39610 511174
rect 39846 510938 70330 511174
rect 70566 510938 101050 511174
rect 101286 510938 131770 511174
rect 132006 510938 162490 511174
rect 162726 510938 193210 511174
rect 193446 510938 223930 511174
rect 224166 510938 254650 511174
rect 254886 510938 285370 511174
rect 285606 510938 316090 511174
rect 316326 510938 346810 511174
rect 347046 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 453424 511174
rect 453660 510938 455862 511174
rect 456098 510938 458300 511174
rect 458536 510938 460738 511174
rect 460974 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 483424 511174
rect 483660 510938 485862 511174
rect 486098 510938 488300 511174
rect 488536 510938 490738 511174
rect 490974 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 39610 510854
rect 39846 510618 70330 510854
rect 70566 510618 101050 510854
rect 101286 510618 131770 510854
rect 132006 510618 162490 510854
rect 162726 510618 193210 510854
rect 193446 510618 223930 510854
rect 224166 510618 254650 510854
rect 254886 510618 285370 510854
rect 285606 510618 316090 510854
rect 316326 510618 346810 510854
rect 347046 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 453424 510854
rect 453660 510618 455862 510854
rect 456098 510618 458300 510854
rect 458536 510618 460738 510854
rect 460974 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 483424 510854
rect 483660 510618 485862 510854
rect 486098 510618 488300 510854
rect 488536 510618 490738 510854
rect 490974 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 24250 507454
rect 24486 507218 54970 507454
rect 55206 507218 85690 507454
rect 85926 507218 116410 507454
rect 116646 507218 147130 507454
rect 147366 507218 177850 507454
rect 178086 507218 208570 507454
rect 208806 507218 239290 507454
rect 239526 507218 270010 507454
rect 270246 507218 300730 507454
rect 300966 507218 331450 507454
rect 331686 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 452205 507454
rect 452441 507218 454643 507454
rect 454879 507218 457081 507454
rect 457317 507218 459519 507454
rect 459755 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 482205 507454
rect 482441 507218 484643 507454
rect 484879 507218 487081 507454
rect 487317 507218 489519 507454
rect 489755 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 24250 507134
rect 24486 506898 54970 507134
rect 55206 506898 85690 507134
rect 85926 506898 116410 507134
rect 116646 506898 147130 507134
rect 147366 506898 177850 507134
rect 178086 506898 208570 507134
rect 208806 506898 239290 507134
rect 239526 506898 270010 507134
rect 270246 506898 300730 507134
rect 300966 506898 331450 507134
rect 331686 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 452205 507134
rect 452441 506898 454643 507134
rect 454879 506898 457081 507134
rect 457317 506898 459519 507134
rect 459755 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 482205 507134
rect 482441 506898 484643 507134
rect 484879 506898 487081 507134
rect 487317 506898 489519 507134
rect 489755 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 39610 475174
rect 39846 474938 70330 475174
rect 70566 474938 101050 475174
rect 101286 474938 131770 475174
rect 132006 474938 162490 475174
rect 162726 474938 193210 475174
rect 193446 474938 223930 475174
rect 224166 474938 254650 475174
rect 254886 474938 285370 475174
rect 285606 474938 316090 475174
rect 316326 474938 346810 475174
rect 347046 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 39610 474854
rect 39846 474618 70330 474854
rect 70566 474618 101050 474854
rect 101286 474618 131770 474854
rect 132006 474618 162490 474854
rect 162726 474618 193210 474854
rect 193446 474618 223930 474854
rect 224166 474618 254650 474854
rect 254886 474618 285370 474854
rect 285606 474618 316090 474854
rect 316326 474618 346810 474854
rect 347046 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 24250 471454
rect 24486 471218 54970 471454
rect 55206 471218 85690 471454
rect 85926 471218 116410 471454
rect 116646 471218 147130 471454
rect 147366 471218 177850 471454
rect 178086 471218 208570 471454
rect 208806 471218 239290 471454
rect 239526 471218 270010 471454
rect 270246 471218 300730 471454
rect 300966 471218 331450 471454
rect 331686 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 24250 471134
rect 24486 470898 54970 471134
rect 55206 470898 85690 471134
rect 85926 470898 116410 471134
rect 116646 470898 147130 471134
rect 147366 470898 177850 471134
rect 178086 470898 208570 471134
rect 208806 470898 239290 471134
rect 239526 470898 270010 471134
rect 270246 470898 300730 471134
rect 300966 470898 331450 471134
rect 331686 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 454007 524426 454054
rect 452982 453818 488426 454007
rect -8726 453771 488426 453818
rect 488662 453771 488746 454007
rect 488982 453818 524426 454007
rect 524662 453818 524746 454054
rect 524982 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect 488982 453771 592650 453818
rect -8726 453734 592650 453771
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 39610 439174
rect 39846 438938 70330 439174
rect 70566 438938 101050 439174
rect 101286 438938 131770 439174
rect 132006 438938 162490 439174
rect 162726 438938 193210 439174
rect 193446 438938 223930 439174
rect 224166 438938 254650 439174
rect 254886 438938 285370 439174
rect 285606 438938 316090 439174
rect 316326 438938 346810 439174
rect 347046 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 426666 439174
rect 426902 438938 432347 439174
rect 432583 438938 438028 439174
rect 438264 438938 443709 439174
rect 443945 438938 475930 439174
rect 476166 438938 480875 439174
rect 481111 438938 485820 439174
rect 486056 438938 490765 439174
rect 491001 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 529426 439174
rect 529662 438938 537867 439174
rect 538103 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546308 439174
rect 546544 438938 554749 439174
rect 554985 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 39610 438854
rect 39846 438618 70330 438854
rect 70566 438618 101050 438854
rect 101286 438618 131770 438854
rect 132006 438618 162490 438854
rect 162726 438618 193210 438854
rect 193446 438618 223930 438854
rect 224166 438618 254650 438854
rect 254886 438618 285370 438854
rect 285606 438618 316090 438854
rect 316326 438618 346810 438854
rect 347046 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 426666 438854
rect 426902 438618 432347 438854
rect 432583 438618 438028 438854
rect 438264 438618 443709 438854
rect 443945 438618 475930 438854
rect 476166 438618 480875 438854
rect 481111 438618 485820 438854
rect 486056 438618 490765 438854
rect 491001 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 529426 438854
rect 529662 438618 537867 438854
rect 538103 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546308 438854
rect 546544 438618 554749 438854
rect 554985 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 24250 435454
rect 24486 435218 54970 435454
rect 55206 435218 85690 435454
rect 85926 435218 116410 435454
rect 116646 435218 147130 435454
rect 147366 435218 177850 435454
rect 178086 435218 208570 435454
rect 208806 435218 239290 435454
rect 239526 435218 270010 435454
rect 270246 435218 300730 435454
rect 300966 435218 331450 435454
rect 331686 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 423826 435454
rect 424062 435218 429507 435454
rect 429743 435218 435188 435454
rect 435424 435218 440869 435454
rect 441105 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 473458 435454
rect 473694 435218 478403 435454
rect 478639 435218 483348 435454
rect 483584 435218 488293 435454
rect 488529 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 525206 435454
rect 525442 435218 533647 435454
rect 533883 435218 542088 435454
rect 542324 435218 550529 435454
rect 550765 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 24250 435134
rect 24486 434898 54970 435134
rect 55206 434898 85690 435134
rect 85926 434898 116410 435134
rect 116646 434898 147130 435134
rect 147366 434898 177850 435134
rect 178086 434898 208570 435134
rect 208806 434898 239290 435134
rect 239526 434898 270010 435134
rect 270246 434898 300730 435134
rect 300966 434898 331450 435134
rect 331686 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 423826 435134
rect 424062 434898 429507 435134
rect 429743 434898 435188 435134
rect 435424 434898 440869 435134
rect 441105 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 473458 435134
rect 473694 434898 478403 435134
rect 478639 434898 483348 435134
rect 483584 434898 488293 435134
rect 488529 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 525206 435134
rect 525442 434898 533647 435134
rect 533883 434898 542088 435134
rect 542324 434898 550529 435134
rect 550765 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 39610 403174
rect 39846 402938 70330 403174
rect 70566 402938 101050 403174
rect 101286 402938 131770 403174
rect 132006 402938 162490 403174
rect 162726 402938 193210 403174
rect 193446 402938 223930 403174
rect 224166 402938 254650 403174
rect 254886 402938 285370 403174
rect 285606 402938 316090 403174
rect 316326 402938 346810 403174
rect 347046 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 39610 402854
rect 39846 402618 70330 402854
rect 70566 402618 101050 402854
rect 101286 402618 131770 402854
rect 132006 402618 162490 402854
rect 162726 402618 193210 402854
rect 193446 402618 223930 402854
rect 224166 402618 254650 402854
rect 254886 402618 285370 402854
rect 285606 402618 316090 402854
rect 316326 402618 346810 402854
rect 347046 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 24250 399454
rect 24486 399218 54970 399454
rect 55206 399218 85690 399454
rect 85926 399218 116410 399454
rect 116646 399218 147130 399454
rect 147366 399218 177850 399454
rect 178086 399218 208570 399454
rect 208806 399218 239290 399454
rect 239526 399218 270010 399454
rect 270246 399218 300730 399454
rect 300966 399218 331450 399454
rect 331686 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 24250 399134
rect 24486 398898 54970 399134
rect 55206 398898 85690 399134
rect 85926 398898 116410 399134
rect 116646 398898 147130 399134
rect 147366 398898 177850 399134
rect 178086 398898 208570 399134
rect 208806 398898 239290 399134
rect 239526 398898 270010 399134
rect 270246 398898 300730 399134
rect 300966 398898 331450 399134
rect 331686 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378243 589182 378334
rect 521262 378098 556706 378243
rect -8726 378014 556706 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 378007 556706 378014
rect 556942 378007 557026 378243
rect 557262 378098 589182 378243
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect 557262 378014 592650 378098
rect 557262 378007 589182 378014
rect 521262 377778 589182 378007
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 39610 367174
rect 39846 366938 70330 367174
rect 70566 366938 101050 367174
rect 101286 366938 131770 367174
rect 132006 366938 162490 367174
rect 162726 366938 193210 367174
rect 193446 366938 223930 367174
rect 224166 366938 254650 367174
rect 254886 366938 285370 367174
rect 285606 366938 316090 367174
rect 316326 366938 346810 367174
rect 347046 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 469610 367174
rect 469846 366938 500330 367174
rect 500566 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 554918 367174
rect 555154 366938 558851 367174
rect 559087 366938 562784 367174
rect 563020 366938 566717 367174
rect 566953 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 39610 366854
rect 39846 366618 70330 366854
rect 70566 366618 101050 366854
rect 101286 366618 131770 366854
rect 132006 366618 162490 366854
rect 162726 366618 193210 366854
rect 193446 366618 223930 366854
rect 224166 366618 254650 366854
rect 254886 366618 285370 366854
rect 285606 366618 316090 366854
rect 316326 366618 346810 366854
rect 347046 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 469610 366854
rect 469846 366618 500330 366854
rect 500566 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 554918 366854
rect 555154 366618 558851 366854
rect 559087 366618 562784 366854
rect 563020 366618 566717 366854
rect 566953 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 24250 363454
rect 24486 363218 54970 363454
rect 55206 363218 85690 363454
rect 85926 363218 116410 363454
rect 116646 363218 147130 363454
rect 147366 363218 177850 363454
rect 178086 363218 208570 363454
rect 208806 363218 239290 363454
rect 239526 363218 270010 363454
rect 270246 363218 300730 363454
rect 300966 363218 331450 363454
rect 331686 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 454250 363454
rect 454486 363218 484970 363454
rect 485206 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 552952 363454
rect 553188 363218 556885 363454
rect 557121 363218 560818 363454
rect 561054 363218 564751 363454
rect 564987 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 24250 363134
rect 24486 362898 54970 363134
rect 55206 362898 85690 363134
rect 85926 362898 116410 363134
rect 116646 362898 147130 363134
rect 147366 362898 177850 363134
rect 178086 362898 208570 363134
rect 208806 362898 239290 363134
rect 239526 362898 270010 363134
rect 270246 362898 300730 363134
rect 300966 362898 331450 363134
rect 331686 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 454250 363134
rect 454486 362898 484970 363134
rect 485206 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 552952 363134
rect 553188 362898 556885 363134
rect 557121 362898 560818 363134
rect 561054 362898 564751 363134
rect 564987 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 39610 331174
rect 39846 330938 70330 331174
rect 70566 330938 101050 331174
rect 101286 330938 131770 331174
rect 132006 330938 162490 331174
rect 162726 330938 193210 331174
rect 193446 330938 223930 331174
rect 224166 330938 254650 331174
rect 254886 330938 285370 331174
rect 285606 330938 316090 331174
rect 316326 330938 346810 331174
rect 347046 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 407932 331174
rect 408168 330938 414878 331174
rect 415114 330938 421824 331174
rect 422060 330938 428770 331174
rect 429006 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 469610 331174
rect 469846 330938 500330 331174
rect 500566 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 39610 330854
rect 39846 330618 70330 330854
rect 70566 330618 101050 330854
rect 101286 330618 131770 330854
rect 132006 330618 162490 330854
rect 162726 330618 193210 330854
rect 193446 330618 223930 330854
rect 224166 330618 254650 330854
rect 254886 330618 285370 330854
rect 285606 330618 316090 330854
rect 316326 330618 346810 330854
rect 347046 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 407932 330854
rect 408168 330618 414878 330854
rect 415114 330618 421824 330854
rect 422060 330618 428770 330854
rect 429006 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 469610 330854
rect 469846 330618 500330 330854
rect 500566 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 24250 327454
rect 24486 327218 54970 327454
rect 55206 327218 85690 327454
rect 85926 327218 116410 327454
rect 116646 327218 147130 327454
rect 147366 327218 177850 327454
rect 178086 327218 208570 327454
rect 208806 327218 239290 327454
rect 239526 327218 270010 327454
rect 270246 327218 300730 327454
rect 300966 327218 331450 327454
rect 331686 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 404459 327454
rect 404695 327218 411405 327454
rect 411641 327218 418351 327454
rect 418587 327218 425297 327454
rect 425533 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 454250 327454
rect 454486 327218 484970 327454
rect 485206 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 24250 327134
rect 24486 326898 54970 327134
rect 55206 326898 85690 327134
rect 85926 326898 116410 327134
rect 116646 326898 147130 327134
rect 147366 326898 177850 327134
rect 178086 326898 208570 327134
rect 208806 326898 239290 327134
rect 239526 326898 270010 327134
rect 270246 326898 300730 327134
rect 300966 326898 331450 327134
rect 331686 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 404459 327134
rect 404695 326898 411405 327134
rect 411641 326898 418351 327134
rect 418587 326898 425297 327134
rect 425533 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 454250 327134
rect 454486 326898 484970 327134
rect 485206 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 39610 295174
rect 39846 294938 70330 295174
rect 70566 294938 101050 295174
rect 101286 294938 131770 295174
rect 132006 294938 162490 295174
rect 162726 294938 193210 295174
rect 193446 294938 223930 295174
rect 224166 294938 254650 295174
rect 254886 294938 285370 295174
rect 285606 294938 316090 295174
rect 316326 294938 346810 295174
rect 347046 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 39610 294854
rect 39846 294618 70330 294854
rect 70566 294618 101050 294854
rect 101286 294618 131770 294854
rect 132006 294618 162490 294854
rect 162726 294618 193210 294854
rect 193446 294618 223930 294854
rect 224166 294618 254650 294854
rect 254886 294618 285370 294854
rect 285606 294618 316090 294854
rect 316326 294618 346810 294854
rect 347046 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 24250 291454
rect 24486 291218 54970 291454
rect 55206 291218 85690 291454
rect 85926 291218 116410 291454
rect 116646 291218 147130 291454
rect 147366 291218 177850 291454
rect 178086 291218 208570 291454
rect 208806 291218 239290 291454
rect 239526 291218 270010 291454
rect 270246 291218 300730 291454
rect 300966 291218 331450 291454
rect 331686 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 24250 291134
rect 24486 290898 54970 291134
rect 55206 290898 85690 291134
rect 85926 290898 116410 291134
rect 116646 290898 147130 291134
rect 147366 290898 177850 291134
rect 178086 290898 208570 291134
rect 208806 290898 239290 291134
rect 239526 290898 270010 291134
rect 270246 290898 300730 291134
rect 300966 290898 331450 291134
rect 331686 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 39610 259174
rect 39846 258938 70330 259174
rect 70566 258938 101050 259174
rect 101286 258938 131770 259174
rect 132006 258938 162490 259174
rect 162726 258938 193210 259174
rect 193446 258938 223930 259174
rect 224166 258938 254650 259174
rect 254886 258938 285370 259174
rect 285606 258938 316090 259174
rect 316326 258938 346810 259174
rect 347046 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 479610 259174
rect 479846 258938 510330 259174
rect 510566 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 39610 258854
rect 39846 258618 70330 258854
rect 70566 258618 101050 258854
rect 101286 258618 131770 258854
rect 132006 258618 162490 258854
rect 162726 258618 193210 258854
rect 193446 258618 223930 258854
rect 224166 258618 254650 258854
rect 254886 258618 285370 258854
rect 285606 258618 316090 258854
rect 316326 258618 346810 258854
rect 347046 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 479610 258854
rect 479846 258618 510330 258854
rect 510566 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 24250 255454
rect 24486 255218 54970 255454
rect 55206 255218 85690 255454
rect 85926 255218 116410 255454
rect 116646 255218 147130 255454
rect 147366 255218 177850 255454
rect 178086 255218 208570 255454
rect 208806 255218 239290 255454
rect 239526 255218 270010 255454
rect 270246 255218 300730 255454
rect 300966 255218 331450 255454
rect 331686 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 464250 255454
rect 464486 255218 494970 255454
rect 495206 255218 525690 255454
rect 525926 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 24250 255134
rect 24486 254898 54970 255134
rect 55206 254898 85690 255134
rect 85926 254898 116410 255134
rect 116646 254898 147130 255134
rect 147366 254898 177850 255134
rect 178086 254898 208570 255134
rect 208806 254898 239290 255134
rect 239526 254898 270010 255134
rect 270246 254898 300730 255134
rect 300966 254898 331450 255134
rect 331686 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 464250 255134
rect 464486 254898 494970 255134
rect 495206 254898 525690 255134
rect 525926 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 39610 223174
rect 39846 222938 70330 223174
rect 70566 222938 101050 223174
rect 101286 222938 131770 223174
rect 132006 222938 162490 223174
rect 162726 222938 193210 223174
rect 193446 222938 223930 223174
rect 224166 222938 254650 223174
rect 254886 222938 285370 223174
rect 285606 222938 316090 223174
rect 316326 222938 346810 223174
rect 347046 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 479610 223174
rect 479846 222938 510330 223174
rect 510566 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 39610 222854
rect 39846 222618 70330 222854
rect 70566 222618 101050 222854
rect 101286 222618 131770 222854
rect 132006 222618 162490 222854
rect 162726 222618 193210 222854
rect 193446 222618 223930 222854
rect 224166 222618 254650 222854
rect 254886 222618 285370 222854
rect 285606 222618 316090 222854
rect 316326 222618 346810 222854
rect 347046 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 479610 222854
rect 479846 222618 510330 222854
rect 510566 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 24250 219454
rect 24486 219218 54970 219454
rect 55206 219218 85690 219454
rect 85926 219218 116410 219454
rect 116646 219218 147130 219454
rect 147366 219218 177850 219454
rect 178086 219218 208570 219454
rect 208806 219218 239290 219454
rect 239526 219218 270010 219454
rect 270246 219218 300730 219454
rect 300966 219218 331450 219454
rect 331686 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 464250 219454
rect 464486 219218 494970 219454
rect 495206 219218 525690 219454
rect 525926 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 24250 219134
rect 24486 218898 54970 219134
rect 55206 218898 85690 219134
rect 85926 218898 116410 219134
rect 116646 218898 147130 219134
rect 147366 218898 177850 219134
rect 178086 218898 208570 219134
rect 208806 218898 239290 219134
rect 239526 218898 270010 219134
rect 270246 218898 300730 219134
rect 300966 218898 331450 219134
rect 331686 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 464250 219134
rect 464486 218898 494970 219134
rect 495206 218898 525690 219134
rect 525926 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 39610 187174
rect 39846 186938 70330 187174
rect 70566 186938 101050 187174
rect 101286 186938 131770 187174
rect 132006 186938 162490 187174
rect 162726 186938 193210 187174
rect 193446 186938 223930 187174
rect 224166 186938 254650 187174
rect 254886 186938 285370 187174
rect 285606 186938 316090 187174
rect 316326 186938 346810 187174
rect 347046 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 39610 186854
rect 39846 186618 70330 186854
rect 70566 186618 101050 186854
rect 101286 186618 131770 186854
rect 132006 186618 162490 186854
rect 162726 186618 193210 186854
rect 193446 186618 223930 186854
rect 224166 186618 254650 186854
rect 254886 186618 285370 186854
rect 285606 186618 316090 186854
rect 316326 186618 346810 186854
rect 347046 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 24250 183454
rect 24486 183218 54970 183454
rect 55206 183218 85690 183454
rect 85926 183218 116410 183454
rect 116646 183218 147130 183454
rect 147366 183218 177850 183454
rect 178086 183218 208570 183454
rect 208806 183218 239290 183454
rect 239526 183218 270010 183454
rect 270246 183218 300730 183454
rect 300966 183218 331450 183454
rect 331686 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 24250 183134
rect 24486 182898 54970 183134
rect 55206 182898 85690 183134
rect 85926 182898 116410 183134
rect 116646 182898 147130 183134
rect 147366 182898 177850 183134
rect 178086 182898 208570 183134
rect 208806 182898 239290 183134
rect 239526 182898 270010 183134
rect 270246 182898 300730 183134
rect 300966 182898 331450 183134
rect 331686 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 39610 151174
rect 39846 150938 70330 151174
rect 70566 150938 101050 151174
rect 101286 150938 131770 151174
rect 132006 150938 162490 151174
rect 162726 150938 193210 151174
rect 193446 150938 223930 151174
rect 224166 150938 254650 151174
rect 254886 150938 285370 151174
rect 285606 150938 316090 151174
rect 316326 150938 346810 151174
rect 347046 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 429610 151174
rect 429846 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 39610 150854
rect 39846 150618 70330 150854
rect 70566 150618 101050 150854
rect 101286 150618 131770 150854
rect 132006 150618 162490 150854
rect 162726 150618 193210 150854
rect 193446 150618 223930 150854
rect 224166 150618 254650 150854
rect 254886 150618 285370 150854
rect 285606 150618 316090 150854
rect 316326 150618 346810 150854
rect 347046 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 429610 150854
rect 429846 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 24250 147454
rect 24486 147218 54970 147454
rect 55206 147218 85690 147454
rect 85926 147218 116410 147454
rect 116646 147218 147130 147454
rect 147366 147218 177850 147454
rect 178086 147218 208570 147454
rect 208806 147218 239290 147454
rect 239526 147218 270010 147454
rect 270246 147218 300730 147454
rect 300966 147218 331450 147454
rect 331686 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 414250 147454
rect 414486 147218 444970 147454
rect 445206 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 24250 147134
rect 24486 146898 54970 147134
rect 55206 146898 85690 147134
rect 85926 146898 116410 147134
rect 116646 146898 147130 147134
rect 147366 146898 177850 147134
rect 178086 146898 208570 147134
rect 208806 146898 239290 147134
rect 239526 146898 270010 147134
rect 270246 146898 300730 147134
rect 300966 146898 331450 147134
rect 331686 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 414250 147134
rect 414486 146898 444970 147134
rect 445206 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 39610 115174
rect 39846 114938 70330 115174
rect 70566 114938 101050 115174
rect 101286 114938 131770 115174
rect 132006 114938 162490 115174
rect 162726 114938 193210 115174
rect 193446 114938 223930 115174
rect 224166 114938 254650 115174
rect 254886 114938 285370 115174
rect 285606 114938 316090 115174
rect 316326 114938 346810 115174
rect 347046 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 499610 115174
rect 499846 114938 530330 115174
rect 530566 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 39610 114854
rect 39846 114618 70330 114854
rect 70566 114618 101050 114854
rect 101286 114618 131770 114854
rect 132006 114618 162490 114854
rect 162726 114618 193210 114854
rect 193446 114618 223930 114854
rect 224166 114618 254650 114854
rect 254886 114618 285370 114854
rect 285606 114618 316090 114854
rect 316326 114618 346810 114854
rect 347046 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 499610 114854
rect 499846 114618 530330 114854
rect 530566 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 24250 111454
rect 24486 111218 54970 111454
rect 55206 111218 85690 111454
rect 85926 111218 116410 111454
rect 116646 111218 147130 111454
rect 147366 111218 177850 111454
rect 178086 111218 208570 111454
rect 208806 111218 239290 111454
rect 239526 111218 270010 111454
rect 270246 111218 300730 111454
rect 300966 111218 331450 111454
rect 331686 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 484250 111454
rect 484486 111218 514970 111454
rect 515206 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 24250 111134
rect 24486 110898 54970 111134
rect 55206 110898 85690 111134
rect 85926 110898 116410 111134
rect 116646 110898 147130 111134
rect 147366 110898 177850 111134
rect 178086 110898 208570 111134
rect 208806 110898 239290 111134
rect 239526 110898 270010 111134
rect 270246 110898 300730 111134
rect 300966 110898 331450 111134
rect 331686 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 484250 111134
rect 484486 110898 514970 111134
rect 515206 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 39610 79174
rect 39846 78938 70330 79174
rect 70566 78938 101050 79174
rect 101286 78938 131770 79174
rect 132006 78938 162490 79174
rect 162726 78938 193210 79174
rect 193446 78938 223930 79174
rect 224166 78938 254650 79174
rect 254886 78938 285370 79174
rect 285606 78938 316090 79174
rect 316326 78938 346810 79174
rect 347046 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 405610 79174
rect 405846 78938 436330 79174
rect 436566 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 39610 78854
rect 39846 78618 70330 78854
rect 70566 78618 101050 78854
rect 101286 78618 131770 78854
rect 132006 78618 162490 78854
rect 162726 78618 193210 78854
rect 193446 78618 223930 78854
rect 224166 78618 254650 78854
rect 254886 78618 285370 78854
rect 285606 78618 316090 78854
rect 316326 78618 346810 78854
rect 347046 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 405610 78854
rect 405846 78618 436330 78854
rect 436566 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 24250 75454
rect 24486 75218 54970 75454
rect 55206 75218 85690 75454
rect 85926 75218 116410 75454
rect 116646 75218 147130 75454
rect 147366 75218 177850 75454
rect 178086 75218 208570 75454
rect 208806 75218 239290 75454
rect 239526 75218 270010 75454
rect 270246 75218 300730 75454
rect 300966 75218 331450 75454
rect 331686 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 390250 75454
rect 390486 75218 420970 75454
rect 421206 75218 451690 75454
rect 451926 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 24250 75134
rect 24486 74898 54970 75134
rect 55206 74898 85690 75134
rect 85926 74898 116410 75134
rect 116646 74898 147130 75134
rect 147366 74898 177850 75134
rect 178086 74898 208570 75134
rect 208806 74898 239290 75134
rect 239526 74898 270010 75134
rect 270246 74898 300730 75134
rect 300966 74898 331450 75134
rect 331686 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 390250 75134
rect 390486 74898 420970 75134
rect 421206 74898 451690 75134
rect 451926 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 405610 43174
rect 405846 42938 436330 43174
rect 436566 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545930 43174
rect 546166 42938 550875 43174
rect 551111 42938 555820 43174
rect 556056 42938 560765 43174
rect 561001 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 405610 42854
rect 405846 42618 436330 42854
rect 436566 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545930 42854
rect 546166 42618 550875 42854
rect 551111 42618 555820 42854
rect 556056 42618 560765 42854
rect 561001 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 390250 39454
rect 390486 39218 420970 39454
rect 421206 39218 451690 39454
rect 451926 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 543458 39454
rect 543694 39218 548403 39454
rect 548639 39218 553348 39454
rect 553584 39218 558293 39454
rect 558529 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 390250 39134
rect 390486 38898 420970 39134
rect 421206 38898 451690 39134
rect 451926 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 543458 39134
rect 543694 38898 548403 39134
rect 548639 38898 553348 39134
rect 553584 38898 558293 39134
rect 558529 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use posit_unit  posit_unit
timestamp 0
transform 1 0 460000 0 1 200000
box 0 2128 70000 67504
use multiplexer  proj_multiplexer
timestamp 0
transform 1 0 450000 0 1 322000
box 0 0 60000 64000
use tholin_avalonsemi_5401  tholin_avalonsemi_5401
timestamp 0
transform 1 0 520000 0 1 425000
box 1066 0 36000 36000
use tholin_avalonsemi_tbb1143  tholin_avalonsemi_tbb1143
timestamp 0
transform 1 0 400000 0 1 305000
box 1066 2048 30000 30000
use tt2_tholin_diceroll  tt2_tholin_diceroll
timestamp 0
transform 1 0 470000 0 1 432000
box 1066 0 21043 22000
use tt2_tholin_multiplexed_counter  tt2_tholin_multiplexed_counter
timestamp 0
transform 1 0 550000 0 1 360000
box 842 0 17098 18000
use tt2_tholin_multiplier  tt2_tholin_multiplier
timestamp 0
transform 1 0 450000 0 1 500000
box 0 0 11118 16584
use tt2_tholin_namebadge  tt2_tholin_namebadge
timestamp 0
transform 1 0 420000 0 1 420000
box 1066 0 23987 25000
use tune_player  tune_player
timestamp 0
transform 1 0 540000 0 1 30000
box 0 2128 21043 19632
use wrapped_6502  wrapped_6502
timestamp 0
transform 1 0 410000 0 1 120000
box 1066 1504 40000 40000
use wrapped_MC14500  wrapped_MC14500
timestamp 0
transform 1 0 480000 0 1 500000
box 566 0 12000 18000
use wrapped_as1802  wrapped_as1802
timestamp 0
transform 1 0 480000 0 1 80000
box 1066 2128 60000 60000
use wrapped_as2650  wrapped_as2650
timestamp 0
transform 1 0 460000 0 1 600000
box 0 0 68816 67992
use wrapped_as512512512  wrapped_as512512512
timestamp 0
transform 1 0 20000 0 1 45000
box 1066 2128 340000 637616
use wrapped_vgatest  wrapped_vgatest
timestamp 0
transform 1 0 386000 0 1 30000
box 749 2128 75000 75000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 674393 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 674393 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 674393 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 674393 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 674393 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 674393 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 674393 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 674393 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 674393 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 31919 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 92137 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 31919 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 157249 434414 422599 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 442833 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 201919 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 385580 470414 601103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 669073 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 82599 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 139281 506414 201919 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 259417 506414 601103 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 669073 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 425068 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 460836 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 674393 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 674393 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 674393 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 674393 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 674393 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 674393 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 674393 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 674393 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 674393 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 30068 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 104460 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 31919 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 157249 441854 422599 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 442833 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 201919 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 259417 477854 322287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 385225 477854 601103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 669073 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 82599 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 139281 513854 201919 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 259417 513854 601103 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 669073 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 -7654 53294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 -7654 89294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 -7654 125294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 -7654 161294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 -7654 197294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 -7654 233294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 -7654 269294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 -7654 305294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 -7654 341294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 -7654 377294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 -7654 413294 31919 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 92137 413294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 -7654 449294 31919 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 92137 449294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 -7654 485294 201919 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 259417 485294 322068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 385580 485294 500068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 517884 485294 601103 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 -7654 521294 82599 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 139281 521294 201919 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 259417 521294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 360068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 377884 557294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 -7654 24734 45068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 -7654 60734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 -7654 96734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 -7654 132734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 -7654 168734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 -7654 204734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 -7654 240734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 -7654 276734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 -7654 312734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 -7654 348734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 -7654 384734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 -7654 420734 31919 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 92137 420734 127767 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 157249 420734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 -7654 456734 31919 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 92137 456734 500068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 517884 456734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 -7654 492734 82599 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 259417 492734 322287 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 385225 492734 601103 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 669073 492734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 -7654 528734 82599 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 259417 528734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 360068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 377884 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 -7654 57014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 -7654 93014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 -7654 129014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 -7654 165014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 -7654 201014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 -7654 237014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 -7654 273014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 -7654 309014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 -7654 345014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 -7654 381014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 -7654 417014 31919 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 92137 417014 127767 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 157249 417014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 -7654 453014 31919 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 92137 453014 500068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 517884 453014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 -7654 489014 82599 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 139281 489014 201919 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 259417 489014 322287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 453692 489014 500068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 517884 489014 601103 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 669073 489014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 -7654 525014 82599 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 139281 525014 201919 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 259417 525014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 30068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 51692 561014 360068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 377884 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 -7654 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 -7654 64454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 674393 64454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 -7654 100454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 674393 100454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 -7654 136454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 674393 136454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 -7654 172454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 674393 172454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 -7654 208454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 674393 208454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 -7654 244454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 674393 244454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 -7654 280454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 674393 280454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 -7654 316454 45068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 -7654 352454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 674393 352454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 -7654 388454 31919 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 92137 388454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 -7654 424454 31919 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 92137 424454 127767 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 157249 424454 420068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 444412 424454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 -7654 460454 500068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 517884 460454 601103 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 669073 460454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 -7654 496454 82599 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 259417 496454 601103 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 669073 496454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 -7654 532454 82599 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 139281 532454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 674393 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 674393 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 674393 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 674393 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 674393 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 674393 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 674393 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 674393 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 674393 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 31919 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 92137 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 31919 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 157249 438134 420068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 444412 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 201919 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 453692 474134 601103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 669073 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 82599 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 139281 510134 201919 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 259417 510134 601103 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 669073 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 30068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 51692 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 -7654 49574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 674393 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 -7654 85574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 674393 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 -7654 121574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 674393 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 -7654 157574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 674393 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 -7654 193574 45068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 684676 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 -7654 229574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 674393 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 -7654 265574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 674393 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 -7654 301574 45068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 684676 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 -7654 337574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 674393 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 -7654 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 -7654 409574 31919 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 92137 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 -7654 445574 31919 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 159644 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 -7654 481574 201919 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 259417 481574 322287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 453692 481574 601103 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 669073 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 -7654 517574 82599 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 139281 517574 201919 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 259417 517574 601103 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 669073 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 -7654 553574 30068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 51692 553574 360068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 377884 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 451808 75336 451808 75336 0 vccd1
rlabel via4 333704 46776 333704 46776 0 vccd2
rlabel via4 521144 666216 521144 666216 0 vdda1
rlabel via4 456584 97656 456584 97656 0 vdda2
rlabel via4 452864 93936 452864 93936 0 vssa1
rlabel via4 460304 101376 460304 101376 0 vssa2
rlabel via4 436448 79056 436448 79056 0 vssd1
rlabel via4 481424 122496 481424 122496 0 vssd2
rlabel metal2 422510 446172 422510 446172 0 design_clk
rlabel metal2 411960 159868 411960 159868 0 dsi_all\[0\]
rlabel metal2 448362 161058 448362 161058 0 dsi_all\[10\]
rlabel metal2 447258 172142 447258 172142 0 dsi_all\[11\]
rlabel metal3 449152 332588 449152 332588 0 dsi_all\[12\]
rlabel metal2 447166 332945 447166 332945 0 dsi_all\[13\]
rlabel metal2 447258 333319 447258 333319 0 dsi_all\[14\]
rlabel metal2 447166 334305 447166 334305 0 dsi_all\[15\]
rlabel metal1 445464 334050 445464 334050 0 dsi_all\[16\]
rlabel metal1 445510 335682 445510 335682 0 dsi_all\[17\]
rlabel metal2 447166 336005 447166 336005 0 dsi_all\[18\]
rlabel metal2 447166 337161 447166 337161 0 dsi_all\[19\]
rlabel metal3 449980 503472 449980 503472 0 dsi_all\[1\]
rlabel metal3 448830 338028 448830 338028 0 dsi_all\[20\]
rlabel metal2 447166 338453 447166 338453 0 dsi_all\[21\]
rlabel metal2 447258 338759 447258 338759 0 dsi_all\[22\]
rlabel metal2 431250 322252 431250 322252 0 dsi_all\[23\]
rlabel metal2 371910 327726 371910 327726 0 dsi_all\[24\]
rlabel metal2 444222 338504 444222 338504 0 dsi_all\[25\]
rlabel metal2 447166 341513 447166 341513 0 dsi_all\[26\]
rlabel metal3 449796 342788 449796 342788 0 dsi_all\[27\]
rlabel metal3 450156 505531 450156 505531 0 dsi_all\[2\]
rlabel metal3 450087 326604 450087 326604 0 dsi_all\[3\]
rlabel metal2 425208 159868 425208 159868 0 dsi_all\[4\]
rlabel metal2 428184 159732 428184 159732 0 dsi_all\[5\]
rlabel metal2 431786 159868 431786 159868 0 dsi_all\[6\]
rlabel metal3 450156 329037 450156 329037 0 dsi_all\[7\]
rlabel metal3 448784 329868 448784 329868 0 dsi_all\[8\]
rlabel metal3 448692 330548 448692 330548 0 dsi_all\[9\]
rlabel metal2 451766 121873 451766 121873 0 dso_6502\[0\]
rlabel via2 452594 135133 452594 135133 0 dso_6502\[10\]
rlabel via2 452594 136493 452594 136493 0 dso_6502\[11\]
rlabel via2 452594 137853 452594 137853 0 dso_6502\[12\]
rlabel via2 452594 139213 452594 139213 0 dso_6502\[13\]
rlabel via2 452594 140573 452594 140573 0 dso_6502\[14\]
rlabel via2 452594 141933 452594 141933 0 dso_6502\[15\]
rlabel metal1 476192 275298 476192 275298 0 dso_6502\[16\]
rlabel metal2 451490 144721 451490 144721 0 dso_6502\[17\]
rlabel metal1 476054 311202 476054 311202 0 dso_6502\[18\]
rlabel metal1 475548 271150 475548 271150 0 dso_6502\[19\]
rlabel metal2 451858 123505 451858 123505 0 dso_6502\[1\]
rlabel metal1 474720 309842 474720 309842 0 dso_6502\[20\]
rlabel metal2 452502 150161 452502 150161 0 dso_6502\[21\]
rlabel metal1 473432 308482 473432 308482 0 dso_6502\[22\]
rlabel metal3 451114 152796 451114 152796 0 dso_6502\[23\]
rlabel via2 451950 154173 451950 154173 0 dso_6502\[24\]
rlabel metal3 450884 155516 450884 155516 0 dso_6502\[25\]
rlabel metal2 451766 157097 451766 157097 0 dso_6502\[26\]
rlabel metal1 488934 319022 488934 319022 0 dso_6502\[2\]
rlabel metal1 489210 319090 489210 319090 0 dso_6502\[3\]
rlabel metal2 489210 300487 489210 300487 0 dso_6502\[4\]
rlabel metal1 471454 268498 471454 268498 0 dso_6502\[5\]
rlabel via2 452410 129693 452410 129693 0 dso_6502\[6\]
rlabel via2 452318 131053 452318 131053 0 dso_6502\[7\]
rlabel metal3 450976 132396 450976 132396 0 dso_6502\[8\]
rlabel via2 452594 133773 452594 133773 0 dso_6502\[9\]
rlabel metal2 503785 385900 503785 385900 0 dso_LCD\[0\]
rlabel metal2 504337 385900 504337 385900 0 dso_LCD\[1\]
rlabel metal2 505310 388576 505310 388576 0 dso_LCD\[2\]
rlabel metal2 505809 385900 505809 385900 0 dso_LCD\[3\]
rlabel metal2 506683 385900 506683 385900 0 dso_LCD\[4\]
rlabel metal2 507327 385900 507327 385900 0 dso_LCD\[5\]
rlabel metal2 508109 385900 508109 385900 0 dso_LCD\[6\]
rlabel metal2 508799 385900 508799 385900 0 dso_LCD\[7\]
rlabel metal3 540492 82348 540492 82348 0 dso_as1802\[0\]
rlabel metal3 540630 102748 540630 102748 0 dso_as1802\[10\]
rlabel metal3 539948 104705 539948 104705 0 dso_as1802\[11\]
rlabel metal3 540676 106828 540676 106828 0 dso_as1802\[12\]
rlabel metal1 500112 319090 500112 319090 0 dso_as1802\[13\]
rlabel metal2 500158 310891 500158 310891 0 dso_as1802\[14\]
rlabel via2 539603 113220 539603 113220 0 dso_as1802\[15\]
rlabel metal3 540078 114988 540078 114988 0 dso_as1802\[16\]
rlabel metal3 540722 117028 540722 117028 0 dso_as1802\[17\]
rlabel via2 539787 119612 539787 119612 0 dso_as1802\[18\]
rlabel via2 539741 121380 539741 121380 0 dso_as1802\[19\]
rlabel metal3 541343 84388 541343 84388 0 dso_as1802\[1\]
rlabel metal2 501814 297019 501814 297019 0 dso_as1802\[20\]
rlabel metal3 541075 137836 541075 137836 0 dso_as1802\[21\]
rlabel metal1 541006 138618 541006 138618 0 dso_as1802\[22\]
rlabel metal2 503010 315685 503010 315685 0 dso_as1802\[23\]
rlabel metal2 502826 320834 502826 320834 0 dso_as1802\[24\]
rlabel metal4 538844 137700 538844 137700 0 dso_as1802\[25\]
rlabel metal1 539258 136578 539258 136578 0 dso_as1802\[26\]
rlabel metal3 540584 86428 540584 86428 0 dso_as1802\[2\]
rlabel metal3 541504 88468 541504 88468 0 dso_as1802\[3\]
rlabel metal3 541228 90508 541228 90508 0 dso_as1802\[4\]
rlabel metal3 541274 92548 541274 92548 0 dso_as1802\[5\]
rlabel metal3 541412 94588 541412 94588 0 dso_as1802\[6\]
rlabel via2 539925 97172 539925 97172 0 dso_as1802\[7\]
rlabel metal3 541320 98668 541320 98668 0 dso_as1802\[8\]
rlabel metal3 541458 100708 541458 100708 0 dso_as1802\[9\]
rlabel metal2 463121 385900 463121 385900 0 dso_as2650\[0\]
rlabel metal1 465014 584426 465014 584426 0 dso_as2650\[10\]
rlabel metal2 471263 385900 471263 385900 0 dso_as2650\[11\]
rlabel metal2 472190 387471 472190 387471 0 dso_as2650\[12\]
rlabel metal2 458988 603908 458988 603908 0 dso_as2650\[13\]
rlabel metal3 459471 635460 459471 635460 0 dso_as2650\[14\]
rlabel metal2 468510 494326 468510 494326 0 dso_as2650\[15\]
rlabel metal2 467130 494326 467130 494326 0 dso_as2650\[16\]
rlabel metal2 461702 493782 461702 493782 0 dso_as2650\[17\]
rlabel metal2 462990 493102 462990 493102 0 dso_as2650\[18\]
rlabel metal2 477105 385900 477105 385900 0 dso_as2650\[19\]
rlabel metal2 463903 385900 463903 385900 0 dso_as2650\[1\]
rlabel metal2 464370 492830 464370 492830 0 dso_as2650\[20\]
rlabel metal2 468602 492184 468602 492184 0 dso_as2650\[21\]
rlabel metal3 459617 655724 459617 655724 0 dso_as2650\[22\]
rlabel metal2 480286 387386 480286 387386 0 dso_as2650\[23\]
rlabel metal2 481022 387250 481022 387250 0 dso_as2650\[24\]
rlabel metal2 481758 387216 481758 387216 0 dso_as2650\[25\]
rlabel metal2 482494 387182 482494 387182 0 dso_as2650\[26\]
rlabel metal2 464547 385900 464547 385900 0 dso_as2650\[2\]
rlabel metal2 465375 385900 465375 385900 0 dso_as2650\[3\]
rlabel metal2 466111 385900 466111 385900 0 dso_as2650\[4\]
rlabel metal2 466801 385900 466801 385900 0 dso_as2650\[5\]
rlabel metal2 467583 385900 467583 385900 0 dso_as2650\[6\]
rlabel metal2 468273 385900 468273 385900 0 dso_as2650\[7\]
rlabel metal2 469246 389607 469246 389607 0 dso_as2650\[8\]
rlabel metal2 469745 385900 469745 385900 0 dso_as2650\[9\]
rlabel metal2 409906 367778 409906 367778 0 dso_as512512512\[0\]
rlabel metal2 447258 371909 447258 371909 0 dso_as512512512\[10\]
rlabel metal2 447166 372283 447166 372283 0 dso_as512512512\[11\]
rlabel metal2 447258 373303 447258 373303 0 dso_as512512512\[12\]
rlabel metal2 447166 373677 447166 373677 0 dso_as512512512\[13\]
rlabel metal2 407790 449854 407790 449854 0 dso_as512512512\[14\]
rlabel metal2 406410 455396 406410 455396 0 dso_as512512512\[15\]
rlabel metal2 447258 376023 447258 376023 0 dso_as512512512\[16\]
rlabel metal2 403650 467126 403650 467126 0 dso_as512512512\[17\]
rlabel metal2 447258 377451 447258 377451 0 dso_as512512512\[18\]
rlabel metal2 367770 478856 367770 478856 0 dso_as512512512\[19\]
rlabel metal1 445556 365602 445556 365602 0 dso_as512512512\[1\]
rlabel metal2 447350 378811 447350 378811 0 dso_as512512512\[20\]
rlabel metal2 370530 490552 370530 490552 0 dso_as512512512\[21\]
rlabel metal2 447534 380171 447534 380171 0 dso_as512512512\[22\]
rlabel metal2 371910 502282 371910 502282 0 dso_as512512512\[23\]
rlabel metal2 447258 380783 447258 380783 0 dso_as512512512\[24\]
rlabel metal2 447258 381871 447258 381871 0 dso_as512512512\[25\]
rlabel metal2 447166 382177 447166 382177 0 dso_as512512512\[26\]
rlabel metal2 447258 383231 447258 383231 0 dso_as512512512\[27\]
rlabel metal1 445510 366962 445510 366962 0 dso_as512512512\[2\]
rlabel metal2 447166 366809 447166 366809 0 dso_as512512512\[3\]
rlabel metal1 445464 368390 445464 368390 0 dso_as512512512\[4\]
rlabel metal2 447166 368203 447166 368203 0 dso_as512512512\[5\]
rlabel metal2 447258 369189 447258 369189 0 dso_as512512512\[6\]
rlabel metal2 447166 369563 447166 369563 0 dso_as512512512\[7\]
rlabel metal2 447258 370549 447258 370549 0 dso_as512512512\[8\]
rlabel metal2 447166 370923 447166 370923 0 dso_as512512512\[9\]
rlabel metal2 483421 385900 483421 385900 0 dso_as5401\[0\]
rlabel metal2 490590 387862 490590 387862 0 dso_as5401\[10\]
rlabel metal2 491471 385900 491471 385900 0 dso_as5401\[11\]
rlabel metal2 492253 385900 492253 385900 0 dso_as5401\[12\]
rlabel metal2 492989 385900 492989 385900 0 dso_as5401\[13\]
rlabel metal2 539067 425068 539067 425068 0 dso_as5401\[14\]
rlabel metal2 540355 425068 540355 425068 0 dso_as5401\[15\]
rlabel metal2 541834 422630 541834 422630 0 dso_as5401\[16\]
rlabel metal2 542931 425068 542931 425068 0 dso_as5401\[17\]
rlabel metal2 544219 425068 544219 425068 0 dso_as5401\[18\]
rlabel metal2 545698 424092 545698 424092 0 dso_as5401\[19\]
rlabel metal2 483966 387386 483966 387386 0 dso_as5401\[1\]
rlabel metal2 546795 425068 546795 425068 0 dso_as5401\[20\]
rlabel metal2 498877 385900 498877 385900 0 dso_as5401\[21\]
rlabel metal2 522330 406130 522330 406130 0 dso_as5401\[22\]
rlabel metal2 500349 385900 500349 385900 0 dso_as5401\[23\]
rlabel metal2 500894 387318 500894 387318 0 dso_as5401\[24\]
rlabel metal2 501821 385900 501821 385900 0 dso_as5401\[25\]
rlabel metal2 502366 387420 502366 387420 0 dso_as5401\[26\]
rlabel metal2 484702 387284 484702 387284 0 dso_as5401\[2\]
rlabel metal2 485438 387250 485438 387250 0 dso_as5401\[3\]
rlabel metal2 486319 385900 486319 385900 0 dso_as5401\[4\]
rlabel metal2 486910 389607 486910 389607 0 dso_as5401\[5\]
rlabel metal2 487837 385900 487837 385900 0 dso_as5401\[6\]
rlabel metal2 488382 387182 488382 387182 0 dso_as5401\[7\]
rlabel metal2 489309 385900 489309 385900 0 dso_as5401\[8\]
rlabel metal2 489854 387216 489854 387216 0 dso_as5401\[9\]
rlabel metal2 522330 369172 522330 369172 0 dso_counter\[0\]
rlabel metal2 565294 360009 565294 360009 0 dso_counter\[10\]
rlabel via1 566766 360077 566766 360077 0 dso_counter\[11\]
rlabel metal2 547262 369206 547262 369206 0 dso_counter\[1\]
rlabel metal3 511282 379780 511282 379780 0 dso_counter\[2\]
rlabel metal3 511650 380324 511650 380324 0 dso_counter\[3\]
rlabel metal3 511604 380868 511604 380868 0 dso_counter\[4\]
rlabel metal2 547170 370396 547170 370396 0 dso_counter\[5\]
rlabel metal2 544410 367268 544410 367268 0 dso_counter\[6\]
rlabel metal3 511236 382500 511236 382500 0 dso_counter\[7\]
rlabel metal3 511650 383044 511650 383044 0 dso_counter\[8\]
rlabel metal2 519754 370804 519754 370804 0 dso_counter\[9\]
rlabel metal2 456734 387522 456734 387522 0 dso_diceroll\[0\]
rlabel metal2 457661 385900 457661 385900 0 dso_diceroll\[1\]
rlabel metal2 458397 385900 458397 385900 0 dso_diceroll\[2\]
rlabel metal2 459133 385900 459133 385900 0 dso_diceroll\[3\]
rlabel metal1 481620 429182 481620 429182 0 dso_diceroll\[4\]
rlabel metal1 484334 429182 484334 429182 0 dso_diceroll\[5\]
rlabel metal2 461150 387420 461150 387420 0 dso_diceroll\[6\]
rlabel metal2 462031 385900 462031 385900 0 dso_diceroll\[7\]
rlabel metal3 449060 352308 449060 352308 0 dso_mc14500\[0\]
rlabel metal3 449152 352988 449152 352988 0 dso_mc14500\[1\]
rlabel metal3 448876 353668 448876 353668 0 dso_mc14500\[2\]
rlabel metal3 448784 354348 448784 354348 0 dso_mc14500\[3\]
rlabel metal2 485224 500140 485224 500140 0 dso_mc14500\[4\]
rlabel metal2 486190 500140 486190 500140 0 dso_mc14500\[5\]
rlabel metal2 487478 500140 487478 500140 0 dso_mc14500\[6\]
rlabel metal2 489102 500140 489102 500140 0 dso_mc14500\[7\]
rlabel metal3 449888 357748 449888 357748 0 dso_mc14500\[8\]
rlabel metal2 450701 500140 450701 500140 0 dso_multiplier\[0\]
rlabel metal2 451773 385900 451773 385900 0 dso_multiplier\[1\]
rlabel metal2 452463 385900 452463 385900 0 dso_multiplier\[2\]
rlabel metal2 453054 387522 453054 387522 0 dso_multiplier\[3\]
rlabel metal2 453889 385900 453889 385900 0 dso_multiplier\[4\]
rlabel metal2 454717 385900 454717 385900 0 dso_multiplier\[5\]
rlabel metal2 455262 389607 455262 389607 0 dso_multiplier\[6\]
rlabel metal2 461058 498552 461058 498552 0 dso_multiplier\[7\]
rlabel metal3 529828 209047 529828 209047 0 dso_posit\[0\]
rlabel metal1 488106 319090 488106 319090 0 dso_posit\[1\]
rlabel metal3 530602 243644 530602 243644 0 dso_posit\[2\]
rlabel metal2 488290 310279 488290 310279 0 dso_posit\[3\]
rlabel metal1 445556 358870 445556 358870 0 dso_tbb1143\[0\]
rlabel metal2 447166 359295 447166 359295 0 dso_tbb1143\[1\]
rlabel metal2 447166 360349 447166 360349 0 dso_tbb1143\[2\]
rlabel metal2 447258 360723 447258 360723 0 dso_tbb1143\[3\]
rlabel metal1 444774 361658 444774 361658 0 dso_tbb1143\[4\]
rlabel metal2 447166 362049 447166 362049 0 dso_tbb1143\[5\]
rlabel metal2 447166 363103 447166 363103 0 dso_tbb1143\[6\]
rlabel metal2 447258 363409 447258 363409 0 dso_tbb1143\[7\]
rlabel metal2 504489 322116 504489 322116 0 dso_tune
rlabel metal2 580198 6715 580198 6715 0 io_in[0]
rlabel metal2 580198 457453 580198 457453 0 io_in[10]
rlabel metal2 519662 416670 519662 416670 0 io_in[11]
rlabel metal2 579922 563703 579922 563703 0 io_in[12]
rlabel metal2 580198 617185 580198 617185 0 io_in[13]
rlabel metal3 581954 670684 581954 670684 0 io_in[14]
rlabel metal3 558923 699788 558923 699788 0 io_in[15]
rlabel metal1 446154 422926 446154 422926 0 io_in[16]
rlabel metal1 444958 387770 444958 387770 0 io_in[17]
rlabel metal2 365010 702178 365010 702178 0 io_in[18]
rlabel metal2 300150 697112 300150 697112 0 io_in[19]
rlabel metal2 580198 46597 580198 46597 0 io_in[1]
rlabel metal2 235198 702076 235198 702076 0 io_in[20]
rlabel metal1 309764 700366 309764 700366 0 io_in[21]
rlabel metal4 444268 510680 444268 510680 0 io_in[22]
rlabel metal2 40526 701940 40526 701940 0 io_in[23]
rlabel metal3 224127 684284 224127 684284 0 io_in[24]
rlabel metal3 1740 632060 1740 632060 0 io_in[25]
rlabel metal3 1786 579972 1786 579972 0 io_in[26]
rlabel metal3 2154 527884 2154 527884 0 io_in[27]
rlabel metal3 2016 475660 2016 475660 0 io_in[28]
rlabel metal3 1924 423572 1924 423572 0 io_in[29]
rlabel metal2 580198 86547 580198 86547 0 io_in[2]
rlabel metal3 2108 371348 2108 371348 0 io_in[30]
rlabel metal2 366942 117742 366942 117742 0 io_in[31]
rlabel metal3 1924 267172 1924 267172 0 io_in[32]
rlabel metal3 2062 214948 2062 214948 0 io_in[33]
rlabel metal3 2200 162860 2200 162860 0 io_in[34]
rlabel metal3 1855 110636 1855 110636 0 io_in[35]
rlabel metal3 1740 71604 1740 71604 0 io_in[36]
rlabel metal3 1602 32436 1602 32436 0 io_in[37]
rlabel metal2 580198 126463 580198 126463 0 io_in[3]
rlabel metal2 580198 166413 580198 166413 0 io_in[4]
rlabel metal2 579830 206329 579830 206329 0 io_in[5]
rlabel via2 580198 245565 580198 245565 0 io_in[6]
rlabel metal2 461610 308244 461610 308244 0 io_in[7]
rlabel metal3 582184 351900 582184 351900 0 io_in[8]
rlabel metal3 582138 404940 582138 404940 0 io_in[9]
rlabel metal2 566490 173502 566490 173502 0 io_oeb[0]
rlabel metal2 580198 484517 580198 484517 0 io_oeb[10]
rlabel metal3 582000 537812 582000 537812 0 io_oeb[11]
rlabel metal2 519570 455226 519570 455226 0 io_oeb[12]
rlabel metal2 580198 643569 580198 643569 0 io_oeb[13]
rlabel metal2 580198 697085 580198 697085 0 io_oeb[14]
rlabel metal3 526769 699788 526769 699788 0 io_oeb[15]
rlabel metal2 447810 528530 447810 528530 0 io_oeb[16]
rlabel metal2 445050 511666 445050 511666 0 io_oeb[17]
rlabel metal2 332534 702144 332534 702144 0 io_oeb[18]
rlabel metal2 267674 694426 267674 694426 0 io_oeb[19]
rlabel metal2 544410 190128 544410 190128 0 io_oeb[1]
rlabel metal2 446614 511462 446614 511462 0 io_oeb[20]
rlabel metal2 137862 702025 137862 702025 0 io_oeb[21]
rlabel metal2 445326 502180 445326 502180 0 io_oeb[22]
rlabel metal2 445234 503285 445234 503285 0 io_oeb[23]
rlabel metal3 1924 658172 1924 658172 0 io_oeb[24]
rlabel metal3 1855 606084 1855 606084 0 io_oeb[25]
rlabel metal3 2200 553860 2200 553860 0 io_oeb[26]
rlabel metal3 2062 501772 2062 501772 0 io_oeb[27]
rlabel metal3 1878 449548 1878 449548 0 io_oeb[28]
rlabel metal1 5290 57902 5290 57902 0 io_oeb[29]
rlabel metal2 579830 112965 579830 112965 0 io_oeb[2]
rlabel metal3 1970 345372 1970 345372 0 io_oeb[30]
rlabel metal3 1832 293148 1832 293148 0 io_oeb[31]
rlabel metal3 2016 241060 2016 241060 0 io_oeb[32]
rlabel metal3 2154 188836 2154 188836 0 io_oeb[33]
rlabel metal3 1786 136748 1786 136748 0 io_oeb[34]
rlabel metal2 21344 55284 21344 55284 0 io_oeb[35]
rlabel metal3 1924 45492 1924 45492 0 io_oeb[36]
rlabel metal3 1878 6460 1878 6460 0 io_oeb[37]
rlabel metal2 580198 152915 580198 152915 0 io_oeb[3]
rlabel metal2 580198 192831 580198 192831 0 io_oeb[4]
rlabel metal2 580198 232781 580198 232781 0 io_oeb[5]
rlabel metal2 579922 272697 579922 272697 0 io_oeb[6]
rlabel metal2 580198 324445 580198 324445 0 io_oeb[7]
rlabel metal2 580198 378301 580198 378301 0 io_oeb[8]
rlabel metal2 579646 431103 579646 431103 0 io_oeb[9]
rlabel metal2 580014 20213 580014 20213 0 io_out[0]
rlabel metal2 580014 471019 580014 471019 0 io_out[10]
rlabel metal3 582046 524484 582046 524484 0 io_out[11]
rlabel metal2 579646 577269 579646 577269 0 io_out[12]
rlabel metal2 580198 630751 580198 630751 0 io_out[13]
rlabel metal2 502274 320246 502274 320246 0 io_out[14]
rlabel metal2 543490 701957 543490 701957 0 io_out[15]
rlabel metal1 445372 419526 445372 419526 0 io_out[16]
rlabel metal2 413678 519836 413678 519836 0 io_out[17]
rlabel metal2 348818 695752 348818 695752 0 io_out[18]
rlabel metal2 283866 697809 283866 697809 0 io_out[19]
rlabel metal2 580198 60163 580198 60163 0 io_out[1]
rlabel metal2 219006 702110 219006 702110 0 io_out[20]
rlabel metal2 154146 702008 154146 702008 0 io_out[21]
rlabel metal2 89194 694392 89194 694392 0 io_out[22]
rlabel metal2 24334 696449 24334 696449 0 io_out[23]
rlabel metal3 2039 671228 2039 671228 0 io_out[24]
rlabel metal3 1947 619140 1947 619140 0 io_out[25]
rlabel metal3 1832 566916 1832 566916 0 io_out[26]
rlabel metal3 2108 514828 2108 514828 0 io_out[27]
rlabel metal3 1970 462604 1970 462604 0 io_out[28]
rlabel metal3 2154 410516 2154 410516 0 io_out[29]
rlabel metal2 580198 100079 580198 100079 0 io_out[2]
rlabel metal1 4140 307734 4140 307734 0 io_out[30]
rlabel metal2 20930 59959 20930 59959 0 io_out[31]
rlabel metal3 1970 254116 1970 254116 0 io_out[32]
rlabel metal3 2108 201892 2108 201892 0 io_out[33]
rlabel metal3 1832 149804 1832 149804 0 io_out[34]
rlabel metal3 1947 97580 1947 97580 0 io_out[35]
rlabel metal3 1878 58548 1878 58548 0 io_out[36]
rlabel metal3 1878 19380 1878 19380 0 io_out[37]
rlabel via2 580198 139349 580198 139349 0 io_out[3]
rlabel metal2 580198 179265 580198 179265 0 io_out[4]
rlabel metal3 581908 219028 581908 219028 0 io_out[5]
rlabel metal2 468786 292905 468786 292905 0 io_out[6]
rlabel metal2 580198 312647 580198 312647 0 io_out[7]
rlabel metal2 580198 364735 580198 364735 0 io_out[8]
rlabel metal3 582092 418268 582092 418268 0 io_out[9]
rlabel metal1 487830 319226 487830 319226 0 oeb_6502
rlabel via2 539373 137700 539373 137700 0 oeb_as1802
rlabel metal2 462622 386978 462622 386978 0 oeb_as2650
rlabel via2 447166 383605 447166 383605 0 oeb_as512512512
rlabel metal2 503293 385900 503293 385900 0 oeb_as5401
rlabel metal3 449980 358428 449980 358428 0 oeb_mc14500
rlabel metal2 448346 159868 448346 159868 0 rst_6502
rlabel metal2 427478 446070 427478 446070 0 rst_LCD
rlabel metal3 449060 345508 449060 345508 0 rst_as1802
rlabel metal3 449221 346188 449221 346188 0 rst_as2650
rlabel metal2 447166 347633 447166 347633 0 rst_as512512512
rlabel metal3 449566 346868 449566 346868 0 rst_as5401
rlabel metal3 449750 348228 449750 348228 0 rst_counter
rlabel metal3 449198 348908 449198 348908 0 rst_diceroll
rlabel metal3 449244 349588 449244 349588 0 rst_mc14500
rlabel metal3 449980 350268 449980 350268 0 rst_posit
rlabel metal2 405957 334900 405957 334900 0 rst_tbb1143
rlabel metal3 448738 351628 448738 351628 0 rst_tune
rlabel metal2 598 1843 598 1843 0 wb_clk_i
rlabel metal2 1702 1911 1702 1911 0 wb_rst_i
rlabel metal2 2898 1979 2898 1979 0 wbs_ack_o
rlabel metal4 509036 312492 509036 312492 0 wbs_adr_i[0]
rlabel metal1 214912 44914 214912 44914 0 wbs_adr_i[10]
rlabel metal1 215280 44982 215280 44982 0 wbs_adr_i[11]
rlabel metal1 217166 45050 217166 45050 0 wbs_adr_i[12]
rlabel metal2 58466 22736 58466 22736 0 wbs_adr_i[13]
rlabel metal2 62054 22770 62054 22770 0 wbs_adr_i[14]
rlabel metal1 222502 45254 222502 45254 0 wbs_adr_i[15]
rlabel metal1 222870 44778 222870 44778 0 wbs_adr_i[16]
rlabel metal1 224526 44710 224526 44710 0 wbs_adr_i[17]
rlabel metal2 76222 22498 76222 22498 0 wbs_adr_i[18]
rlabel metal2 79718 21240 79718 21240 0 wbs_adr_i[19]
rlabel metal1 194304 42058 194304 42058 0 wbs_adr_i[1]
rlabel metal2 83306 21274 83306 21274 0 wbs_adr_i[20]
rlabel metal2 373474 171428 373474 171428 0 wbs_adr_i[21]
rlabel metal2 373566 171496 373566 171496 0 wbs_adr_i[22]
rlabel metal2 93978 21376 93978 21376 0 wbs_adr_i[23]
rlabel metal2 97474 21410 97474 21410 0 wbs_adr_i[24]
rlabel metal2 101062 21444 101062 21444 0 wbs_adr_i[25]
rlabel metal2 370806 171530 370806 171530 0 wbs_adr_i[26]
rlabel metal2 368046 171428 368046 171428 0 wbs_adr_i[27]
rlabel metal2 368230 171530 368230 171530 0 wbs_adr_i[28]
rlabel metal2 115230 21172 115230 21172 0 wbs_adr_i[29]
rlabel metal2 17066 1775 17066 1775 0 wbs_adr_i[2]
rlabel metal2 118818 20186 118818 20186 0 wbs_adr_i[30]
rlabel metal2 122314 19812 122314 19812 0 wbs_adr_i[31]
rlabel metal2 21850 1962 21850 1962 0 wbs_adr_i[3]
rlabel metal1 194488 39406 194488 39406 0 wbs_adr_i[4]
rlabel metal2 30130 2030 30130 2030 0 wbs_adr_i[5]
rlabel metal2 507702 309536 507702 309536 0 wbs_adr_i[6]
rlabel metal2 37214 19948 37214 19948 0 wbs_adr_i[7]
rlabel metal2 40710 19982 40710 19982 0 wbs_adr_i[8]
rlabel metal2 44298 1996 44298 1996 0 wbs_adr_i[9]
rlabel metal2 4094 19846 4094 19846 0 wbs_cyc_i
rlabel metal2 8786 2183 8786 2183 0 wbs_dat_i[0]
rlabel metal1 206448 39678 206448 39678 0 wbs_dat_i[10]
rlabel metal2 366574 168708 366574 168708 0 wbs_dat_i[11]
rlabel metal2 56074 20084 56074 20084 0 wbs_dat_i[12]
rlabel metal2 59662 20118 59662 20118 0 wbs_dat_i[13]
rlabel metal2 63250 20152 63250 20152 0 wbs_dat_i[14]
rlabel metal2 370714 165648 370714 165648 0 wbs_dat_i[15]
rlabel metal2 369334 165886 369334 165886 0 wbs_dat_i[16]
rlabel metal2 372278 165750 372278 165750 0 wbs_dat_i[17]
rlabel metal2 77418 18554 77418 18554 0 wbs_dat_i[18]
rlabel metal2 80914 18588 80914 18588 0 wbs_dat_i[19]
rlabel metal2 372002 149192 372002 149192 0 wbs_dat_i[1]
rlabel metal1 229632 36890 229632 36890 0 wbs_dat_i[20]
rlabel metal1 231426 37026 231426 37026 0 wbs_dat_i[21]
rlabel metal2 520582 328406 520582 328406 0 wbs_dat_i[22]
rlabel metal2 95174 18724 95174 18724 0 wbs_dat_i[23]
rlabel metal2 98670 18758 98670 18758 0 wbs_dat_i[24]
rlabel metal2 102258 18792 102258 18792 0 wbs_dat_i[25]
rlabel metal2 520398 330242 520398 330242 0 wbs_dat_i[26]
rlabel metal1 447994 292230 447994 292230 0 wbs_dat_i[27]
rlabel metal1 446246 292298 446246 292298 0 wbs_dat_i[28]
rlabel metal2 116426 17364 116426 17364 0 wbs_dat_i[29]
rlabel metal2 18262 17092 18262 17092 0 wbs_dat_i[2]
rlabel metal2 119922 17398 119922 17398 0 wbs_dat_i[30]
rlabel metal1 447534 386546 447534 386546 0 wbs_dat_i[31]
rlabel metal2 23046 17058 23046 17058 0 wbs_dat_i[3]
rlabel metal2 384330 148002 384330 148002 0 wbs_dat_i[4]
rlabel metal2 386078 163166 386078 163166 0 wbs_dat_i[5]
rlabel metal2 519754 314568 519754 314568 0 wbs_dat_i[6]
rlabel metal2 38410 2064 38410 2064 0 wbs_dat_i[7]
rlabel metal2 41906 17194 41906 17194 0 wbs_dat_i[8]
rlabel metal2 45494 17228 45494 17228 0 wbs_dat_i[9]
rlabel metal2 385802 154105 385802 154105 0 wbs_dat_o[0]
rlabel metal2 507334 305422 507334 305422 0 wbs_dat_o[10]
rlabel metal2 365010 152728 365010 152728 0 wbs_dat_o[11]
rlabel metal2 57270 15732 57270 15732 0 wbs_dat_o[12]
rlabel metal2 60858 15766 60858 15766 0 wbs_dat_o[13]
rlabel metal2 64354 15800 64354 15800 0 wbs_dat_o[14]
rlabel metal2 521962 320586 521962 320586 0 wbs_dat_o[15]
rlabel metal1 449052 289646 449052 289646 0 wbs_dat_o[16]
rlabel metal2 75026 2200 75026 2200 0 wbs_dat_o[17]
rlabel metal2 78614 15902 78614 15902 0 wbs_dat_o[18]
rlabel metal2 82110 2234 82110 2234 0 wbs_dat_o[19]
rlabel metal2 385894 160004 385894 160004 0 wbs_dat_o[1]
rlabel metal2 384790 160616 384790 160616 0 wbs_dat_o[20]
rlabel metal2 89194 1860 89194 1860 0 wbs_dat_o[21]
rlabel metal2 521870 326298 521870 326298 0 wbs_dat_o[22]
rlabel metal2 96278 16004 96278 16004 0 wbs_dat_o[23]
rlabel metal2 99866 15664 99866 15664 0 wbs_dat_o[24]
rlabel metal2 103362 1826 103362 1826 0 wbs_dat_o[25]
rlabel metal2 365286 157522 365286 157522 0 wbs_dat_o[26]
rlabel metal2 110538 1792 110538 1792 0 wbs_dat_o[27]
rlabel metal2 114034 14576 114034 14576 0 wbs_dat_o[28]
rlabel metal2 117622 14644 117622 14644 0 wbs_dat_o[29]
rlabel metal2 19458 14372 19458 14372 0 wbs_dat_o[2]
rlabel metal2 121118 14610 121118 14610 0 wbs_dat_o[30]
rlabel metal1 443486 386478 443486 386478 0 wbs_dat_o[31]
rlabel metal2 24242 1894 24242 1894 0 wbs_dat_o[3]
rlabel metal2 520766 310658 520766 310658 0 wbs_dat_o[4]
rlabel metal1 443578 307054 443578 307054 0 wbs_dat_o[5]
rlabel metal2 36018 14508 36018 14508 0 wbs_dat_o[6]
rlabel metal2 39606 2098 39606 2098 0 wbs_dat_o[7]
rlabel metal2 43102 14304 43102 14304 0 wbs_dat_o[8]
rlabel metal2 46690 2132 46690 2132 0 wbs_dat_o[9]
rlabel metal2 5290 14338 5290 14338 0 wbs_stb_i
rlabel metal2 6486 1792 6486 1792 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
