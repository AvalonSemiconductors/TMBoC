magic
tech sky130B
magscale 1 2
timestamp 1683540956
<< viali >>
rect 11989 22117 12023 22151
rect 12357 22049 12391 22083
rect 12449 22049 12483 22083
rect 2053 21981 2087 22015
rect 4537 21981 4571 22015
rect 4804 21981 4838 22015
rect 12173 21981 12207 22015
rect 13001 21981 13035 22015
rect 13645 21981 13679 22015
rect 20453 21981 20487 22015
rect 20637 21981 20671 22015
rect 22477 21981 22511 22015
rect 2320 21913 2354 21947
rect 7113 21913 7147 21947
rect 7665 21913 7699 21947
rect 13185 21913 13219 21947
rect 17049 21913 17083 21947
rect 17601 21913 17635 21947
rect 22661 21913 22695 21947
rect 3433 21845 3467 21879
rect 5917 21845 5951 21879
rect 7757 21845 7791 21879
rect 14289 21845 14323 21879
rect 15025 21845 15059 21879
rect 15669 21845 15703 21879
rect 17693 21845 17727 21879
rect 20545 21845 20579 21879
rect 18613 21641 18647 21675
rect 19257 21641 19291 21675
rect 21097 21641 21131 21675
rect 22385 21641 22419 21675
rect 3902 21573 3936 21607
rect 6828 21573 6862 21607
rect 8668 21573 8702 21607
rect 15945 21573 15979 21607
rect 20729 21573 20763 21607
rect 4169 21505 4203 21539
rect 5742 21505 5776 21539
rect 6009 21505 6043 21539
rect 12357 21505 12391 21539
rect 12449 21505 12483 21539
rect 12541 21505 12575 21539
rect 12725 21505 12759 21539
rect 13185 21505 13219 21539
rect 14197 21505 14231 21539
rect 14657 21505 14691 21539
rect 14841 21505 14875 21539
rect 17785 21505 17819 21539
rect 17877 21505 17911 21539
rect 17969 21505 18003 21539
rect 18153 21505 18187 21539
rect 20269 21505 20303 21539
rect 20913 21505 20947 21539
rect 6561 21437 6595 21471
rect 8401 21437 8435 21471
rect 13921 21437 13955 21471
rect 17509 21437 17543 21471
rect 18797 21437 18831 21471
rect 18889 21437 18923 21471
rect 20085 21437 20119 21471
rect 12173 21369 12207 21403
rect 16313 21369 16347 21403
rect 2789 21301 2823 21335
rect 4629 21301 4663 21335
rect 7941 21301 7975 21335
rect 9781 21301 9815 21335
rect 14749 21301 14783 21335
rect 15761 21301 15795 21335
rect 15945 21301 15979 21335
rect 16957 21301 16991 21335
rect 12081 21097 12115 21131
rect 14749 21097 14783 21131
rect 15393 21097 15427 21131
rect 17141 21097 17175 21131
rect 19441 21097 19475 21131
rect 9137 21029 9171 21063
rect 13185 21029 13219 21063
rect 17417 21029 17451 21063
rect 11437 20961 11471 20995
rect 22661 20961 22695 20995
rect 1961 20893 1995 20927
rect 7205 20893 7239 20927
rect 10517 20893 10551 20927
rect 11345 20893 11379 20927
rect 12173 20893 12207 20927
rect 12633 20893 12667 20927
rect 12909 20893 12943 20927
rect 13185 20893 13219 20927
rect 14565 20893 14599 20927
rect 14749 20893 14783 20927
rect 15485 20893 15519 20927
rect 15577 20893 15611 20927
rect 15853 20893 15887 20927
rect 16221 20893 16255 20927
rect 17325 20893 17359 20927
rect 17509 20893 17543 20927
rect 17601 20893 17635 20927
rect 17785 20893 17819 20927
rect 18429 20893 18463 20927
rect 18613 20893 18647 20927
rect 19625 20893 19659 20927
rect 19717 20893 19751 20927
rect 19901 20893 19935 20927
rect 19993 20893 20027 20927
rect 20453 20893 20487 20927
rect 22569 20893 22603 20927
rect 2228 20825 2262 20859
rect 6960 20825 6994 20859
rect 10272 20825 10306 20859
rect 13461 20825 13495 20859
rect 18521 20825 18555 20859
rect 20729 20825 20763 20859
rect 21925 20825 21959 20859
rect 3341 20757 3375 20791
rect 5825 20757 5859 20791
rect 8493 20757 8527 20791
rect 14933 20757 14967 20791
rect 3065 20553 3099 20587
rect 11069 20553 11103 20587
rect 20085 20553 20119 20587
rect 20729 20553 20763 20587
rect 22661 20553 22695 20587
rect 13553 20485 13587 20519
rect 22109 20485 22143 20519
rect 4353 20417 4387 20451
rect 8484 20417 8518 20451
rect 10057 20417 10091 20451
rect 12541 20417 12575 20451
rect 13737 20417 13771 20451
rect 13829 20417 13863 20451
rect 14289 20417 14323 20451
rect 14473 20417 14507 20451
rect 15117 20417 15151 20451
rect 15301 20417 15335 20451
rect 15393 20417 15427 20451
rect 19993 20417 20027 20451
rect 20177 20417 20211 20451
rect 22017 20417 22051 20451
rect 22661 20417 22695 20451
rect 22845 20417 22879 20451
rect 8217 20349 8251 20383
rect 12633 20349 12667 20383
rect 12817 20349 12851 20383
rect 14381 20349 14415 20383
rect 15209 20349 15243 20383
rect 9597 20281 9631 20315
rect 13553 20281 13587 20315
rect 16037 20281 16071 20315
rect 19349 20281 19383 20315
rect 12173 20213 12207 20247
rect 14933 20213 14967 20247
rect 11437 20009 11471 20043
rect 11989 20009 12023 20043
rect 13277 20009 13311 20043
rect 15577 20009 15611 20043
rect 19441 20009 19475 20043
rect 12265 19941 12299 19975
rect 3433 19873 3467 19907
rect 12357 19873 12391 19907
rect 12449 19873 12483 19907
rect 15117 19873 15151 19907
rect 6745 19805 6779 19839
rect 7205 19805 7239 19839
rect 9137 19805 9171 19839
rect 9413 19805 9447 19839
rect 12173 19805 12207 19839
rect 12633 19805 12667 19839
rect 13461 19805 13495 19839
rect 14381 19805 14415 19839
rect 14565 19805 14599 19839
rect 19625 19805 19659 19839
rect 19901 19805 19935 19839
rect 3166 19737 3200 19771
rect 6478 19737 6512 19771
rect 7472 19737 7506 19771
rect 2053 19669 2087 19703
rect 5365 19669 5399 19703
rect 8585 19669 8619 19703
rect 10517 19669 10551 19703
rect 14473 19669 14507 19703
rect 19809 19669 19843 19703
rect 9597 19465 9631 19499
rect 13001 19465 13035 19499
rect 17049 19465 17083 19499
rect 18153 19465 18187 19499
rect 4629 19397 4663 19431
rect 22201 19397 22235 19431
rect 2973 19329 3007 19363
rect 8217 19329 8251 19363
rect 8484 19329 8518 19363
rect 12633 19329 12667 19363
rect 14473 19329 14507 19363
rect 18337 19329 18371 19363
rect 19533 19329 19567 19363
rect 19717 19329 19751 19363
rect 19809 19329 19843 19363
rect 22017 19329 22051 19363
rect 3249 19261 3283 19295
rect 10149 19261 10183 19295
rect 12540 19261 12574 19295
rect 12725 19261 12759 19295
rect 12825 19261 12859 19295
rect 14749 19261 14783 19295
rect 15393 19261 15427 19295
rect 17233 19261 17267 19295
rect 17325 19261 17359 19295
rect 17417 19261 17451 19295
rect 17509 19261 17543 19295
rect 18521 19261 18555 19295
rect 13553 19193 13587 19227
rect 14657 19193 14691 19227
rect 14565 19125 14599 19159
rect 15853 19125 15887 19159
rect 19349 19125 19383 19159
rect 22293 19125 22327 19159
rect 5825 18921 5859 18955
rect 7665 18921 7699 18955
rect 14289 18921 14323 18955
rect 16589 18921 16623 18955
rect 18889 18921 18923 18955
rect 19441 18921 19475 18955
rect 2053 18785 2087 18819
rect 12909 18785 12943 18819
rect 13001 18785 13035 18819
rect 16405 18785 16439 18819
rect 6377 18717 6411 18751
rect 9137 18717 9171 18751
rect 12817 18717 12851 18751
rect 13093 18717 13127 18751
rect 14473 18717 14507 18751
rect 14933 18717 14967 18751
rect 16865 18717 16899 18751
rect 18245 18717 18279 18751
rect 18393 18717 18427 18751
rect 18613 18717 18647 18751
rect 18751 18717 18785 18751
rect 19717 18717 19751 18751
rect 19809 18717 19843 18751
rect 19901 18717 19935 18751
rect 20085 18717 20119 18751
rect 20545 18717 20579 18751
rect 2320 18649 2354 18683
rect 9404 18649 9438 18683
rect 14565 18649 14599 18683
rect 14657 18649 14691 18683
rect 14775 18649 14809 18683
rect 18521 18649 18555 18683
rect 3433 18581 3467 18615
rect 10517 18581 10551 18615
rect 13277 18581 13311 18615
rect 15393 18581 15427 18615
rect 16773 18581 16807 18615
rect 9137 18377 9171 18411
rect 12081 18377 12115 18411
rect 13737 18377 13771 18411
rect 14105 18377 14139 18411
rect 15209 18377 15243 18411
rect 16957 18377 16991 18411
rect 18981 18377 19015 18411
rect 19533 18377 19567 18411
rect 3332 18309 3366 18343
rect 14565 18309 14599 18343
rect 14657 18309 14691 18343
rect 7849 18241 7883 18275
rect 12265 18241 12299 18275
rect 12357 18241 12391 18275
rect 12633 18241 12667 18275
rect 13185 18241 13219 18275
rect 13645 18241 13679 18275
rect 13921 18241 13955 18275
rect 14933 18241 14967 18275
rect 16865 18241 16899 18275
rect 17233 18241 17267 18275
rect 18061 18241 18095 18275
rect 19717 18241 19751 18275
rect 19901 18241 19935 18275
rect 19993 18241 20027 18275
rect 3065 18173 3099 18207
rect 12541 18173 12575 18207
rect 15025 18173 15059 18207
rect 17417 18173 17451 18207
rect 18337 18173 18371 18207
rect 4445 18037 4479 18071
rect 15669 18037 15703 18071
rect 16313 18037 16347 18071
rect 17877 18037 17911 18071
rect 18245 18037 18279 18071
rect 11713 17833 11747 17867
rect 13185 17833 13219 17867
rect 17509 17833 17543 17867
rect 21465 17833 21499 17867
rect 22661 17833 22695 17867
rect 12725 17765 12759 17799
rect 16773 17765 16807 17799
rect 13553 17697 13587 17731
rect 14841 17697 14875 17731
rect 17601 17697 17635 17731
rect 7113 17629 7147 17663
rect 9137 17629 9171 17663
rect 11161 17629 11195 17663
rect 11621 17629 11655 17663
rect 12265 17629 12299 17663
rect 12357 17629 12391 17663
rect 12541 17629 12575 17663
rect 13369 17629 13403 17663
rect 13461 17629 13495 17663
rect 13645 17629 13679 17663
rect 15025 17629 15059 17663
rect 15669 17629 15703 17663
rect 15945 17629 15979 17663
rect 16589 17629 16623 17663
rect 16865 17629 16899 17663
rect 17693 17629 17727 17663
rect 22017 17629 22051 17663
rect 22201 17629 22235 17663
rect 22293 17629 22327 17663
rect 22385 17629 22419 17663
rect 6868 17561 6902 17595
rect 9404 17561 9438 17595
rect 16405 17561 16439 17595
rect 5733 17493 5767 17527
rect 8401 17493 8435 17527
rect 10517 17493 10551 17527
rect 15485 17493 15519 17527
rect 15853 17493 15887 17527
rect 17325 17493 17359 17527
rect 12357 17289 12391 17323
rect 16221 17289 16255 17323
rect 19349 17289 19383 17323
rect 19993 17289 20027 17323
rect 13921 17221 13955 17255
rect 14841 17221 14875 17255
rect 17141 17221 17175 17255
rect 2973 17153 3007 17187
rect 6828 17153 6862 17187
rect 8760 17153 8794 17187
rect 13004 17153 13038 17187
rect 13093 17153 13127 17187
rect 13277 17153 13311 17187
rect 13369 17153 13403 17187
rect 13829 17153 13863 17187
rect 14013 17153 14047 17187
rect 14705 17153 14739 17187
rect 14933 17153 14967 17187
rect 15116 17153 15150 17187
rect 15202 17153 15236 17187
rect 16129 17153 16163 17187
rect 16313 17153 16347 17187
rect 17049 17153 17083 17187
rect 17233 17153 17267 17187
rect 19257 17153 19291 17187
rect 19533 17153 19567 17187
rect 19717 17153 19751 17187
rect 20913 17153 20947 17187
rect 22201 17153 22235 17187
rect 22385 17153 22419 17187
rect 22477 17153 22511 17187
rect 3249 17085 3283 17119
rect 6561 17085 6595 17119
rect 8493 17085 8527 17119
rect 19625 17085 19659 17119
rect 20637 17085 20671 17119
rect 20729 17017 20763 17051
rect 4537 16949 4571 16983
rect 7941 16949 7975 16983
rect 9873 16949 9907 16983
rect 12817 16949 12851 16983
rect 14565 16949 14599 16983
rect 20821 16949 20855 16983
rect 22017 16949 22051 16983
rect 22109 16745 22143 16779
rect 22293 16745 22327 16779
rect 11345 16677 11379 16711
rect 15945 16677 15979 16711
rect 18889 16677 18923 16711
rect 19717 16677 19751 16711
rect 20637 16677 20671 16711
rect 5365 16609 5399 16643
rect 8309 16609 8343 16643
rect 9137 16609 9171 16643
rect 9413 16609 9447 16643
rect 12541 16609 12575 16643
rect 12633 16609 12667 16643
rect 12725 16609 12759 16643
rect 12817 16609 12851 16643
rect 13369 16609 13403 16643
rect 17141 16609 17175 16643
rect 17233 16609 17267 16643
rect 19901 16609 19935 16643
rect 3433 16541 3467 16575
rect 5109 16541 5143 16575
rect 8033 16541 8067 16575
rect 17417 16541 17451 16575
rect 17509 16541 17543 16575
rect 18153 16541 18187 16575
rect 19625 16541 19659 16575
rect 19809 16541 19843 16575
rect 20085 16507 20119 16541
rect 3188 16473 3222 16507
rect 6653 16473 6687 16507
rect 10793 16473 10827 16507
rect 14841 16473 14875 16507
rect 15485 16473 15519 16507
rect 17049 16473 17083 16507
rect 21925 16473 21959 16507
rect 2053 16405 2087 16439
rect 3985 16405 4019 16439
rect 12357 16405 12391 16439
rect 14381 16405 14415 16439
rect 18061 16405 18095 16439
rect 19441 16405 19475 16439
rect 22125 16405 22159 16439
rect 9137 16201 9171 16235
rect 15393 16201 15427 16235
rect 18337 16201 18371 16235
rect 20729 16201 20763 16235
rect 22385 16201 22419 16235
rect 4353 16133 4387 16167
rect 7849 16133 7883 16167
rect 12265 16065 12299 16099
rect 12633 16065 12667 16099
rect 15577 16065 15611 16099
rect 15669 16065 15703 16099
rect 15945 16065 15979 16099
rect 17325 16065 17359 16099
rect 17601 16065 17635 16099
rect 18521 16065 18555 16099
rect 20177 16065 20211 16099
rect 20269 16065 20303 16099
rect 20453 16065 20487 16099
rect 20545 16065 20579 16099
rect 22109 16065 22143 16099
rect 22937 16065 22971 16099
rect 14565 15997 14599 16031
rect 19073 15997 19107 16031
rect 3065 15861 3099 15895
rect 13921 15861 13955 15895
rect 15853 15861 15887 15895
rect 17417 15861 17451 15895
rect 17785 15861 17819 15895
rect 19717 15861 19751 15895
rect 13185 15657 13219 15691
rect 17049 15657 17083 15691
rect 18889 15657 18923 15691
rect 21833 15657 21867 15691
rect 14473 15589 14507 15623
rect 19441 15589 19475 15623
rect 6745 15521 6779 15555
rect 9137 15521 9171 15555
rect 12357 15521 12391 15555
rect 13553 15521 13587 15555
rect 15025 15521 15059 15555
rect 15945 15521 15979 15555
rect 17693 15521 17727 15555
rect 18797 15521 18831 15555
rect 2421 15453 2455 15487
rect 5641 15453 5675 15487
rect 9404 15453 9438 15487
rect 12265 15453 12299 15487
rect 12541 15453 12575 15487
rect 13369 15453 13403 15487
rect 13461 15453 13495 15487
rect 13645 15453 13679 15487
rect 15669 15453 15703 15487
rect 17233 15453 17267 15487
rect 18889 15453 18923 15487
rect 19625 15453 19659 15487
rect 19717 15453 19751 15487
rect 19901 15453 19935 15487
rect 19993 15453 20027 15487
rect 21373 15453 21407 15487
rect 22017 15453 22051 15487
rect 22293 15453 22327 15487
rect 5273 15385 5307 15419
rect 7012 15385 7046 15419
rect 11805 15385 11839 15419
rect 14841 15385 14875 15419
rect 17325 15385 17359 15419
rect 17417 15385 17451 15419
rect 17555 15385 17589 15419
rect 21097 15385 21131 15419
rect 2237 15317 2271 15351
rect 8125 15317 8159 15351
rect 10517 15317 10551 15351
rect 11161 15317 11195 15351
rect 12725 15317 12759 15351
rect 14933 15317 14967 15351
rect 18521 15317 18555 15351
rect 22201 15317 22235 15351
rect 2421 15113 2455 15147
rect 14841 15113 14875 15147
rect 16865 15113 16899 15147
rect 22569 15113 22603 15147
rect 2145 15045 2179 15079
rect 5641 15045 5675 15079
rect 6745 15045 6779 15079
rect 7297 15045 7331 15079
rect 9404 15045 9438 15079
rect 13553 15045 13587 15079
rect 14565 15045 14599 15079
rect 1869 14977 1903 15011
rect 2053 14977 2087 15011
rect 2237 14977 2271 15011
rect 6561 14977 6595 15011
rect 6837 14977 6871 15011
rect 9137 14977 9171 15011
rect 11805 14977 11839 15011
rect 12909 14977 12943 15011
rect 13277 14977 13311 15011
rect 14289 14977 14323 15011
rect 14473 14977 14507 15011
rect 14657 14977 14691 15011
rect 15945 14977 15979 15011
rect 16037 14977 16071 15011
rect 16221 14977 16255 15011
rect 16313 14977 16347 15011
rect 17233 14977 17267 15011
rect 17325 14977 17359 15011
rect 18245 14977 18279 15011
rect 18429 14977 18463 15011
rect 19257 14977 19291 15011
rect 19441 14977 19475 15011
rect 21465 14977 21499 15011
rect 22293 14977 22327 15011
rect 22845 14977 22879 15011
rect 3065 14909 3099 14943
rect 3341 14909 3375 14943
rect 12081 14909 12115 14943
rect 13369 14909 13403 14943
rect 17049 14909 17083 14943
rect 17141 14909 17175 14943
rect 19625 14909 19659 14943
rect 22017 14909 22051 14943
rect 22661 14909 22695 14943
rect 4629 14841 4663 14875
rect 18337 14841 18371 14875
rect 5733 14773 5767 14807
rect 6561 14773 6595 14807
rect 10517 14773 10551 14807
rect 15761 14773 15795 14807
rect 20913 14773 20947 14807
rect 2329 14569 2363 14603
rect 5089 14569 5123 14603
rect 6101 14569 6135 14603
rect 9137 14569 9171 14603
rect 13645 14569 13679 14603
rect 14565 14569 14599 14603
rect 15669 14569 15703 14603
rect 20085 14569 20119 14603
rect 22293 14569 22327 14603
rect 10425 14501 10459 14535
rect 11621 14433 11655 14467
rect 12725 14433 12759 14467
rect 14933 14433 14967 14467
rect 1777 14365 1811 14399
rect 2145 14365 2179 14399
rect 3433 14365 3467 14399
rect 4169 14365 4203 14399
rect 4537 14365 4571 14399
rect 5273 14365 5307 14399
rect 5365 14365 5399 14399
rect 5641 14365 5675 14399
rect 6285 14365 6319 14399
rect 6653 14365 6687 14399
rect 7849 14365 7883 14399
rect 7941 14365 7975 14399
rect 8125 14365 8159 14399
rect 8227 14375 8261 14409
rect 9321 14365 9355 14399
rect 9689 14365 9723 14399
rect 10701 14365 10735 14399
rect 11713 14365 11747 14399
rect 11989 14365 12023 14399
rect 12081 14365 12115 14399
rect 14749 14365 14783 14399
rect 15669 14365 15703 14399
rect 15945 14365 15979 14399
rect 19441 14365 19475 14399
rect 19533 14365 19567 14399
rect 19901 14365 19935 14399
rect 21649 14365 21683 14399
rect 21742 14365 21776 14399
rect 22017 14365 22051 14399
rect 22155 14365 22189 14399
rect 22937 14365 22971 14399
rect 1961 14297 1995 14331
rect 2053 14297 2087 14331
rect 3157 14297 3191 14331
rect 4261 14297 4295 14331
rect 4353 14297 4387 14331
rect 5457 14297 5491 14331
rect 6377 14297 6411 14331
rect 6469 14297 6503 14331
rect 9413 14297 9447 14331
rect 9505 14297 9539 14331
rect 10885 14297 10919 14331
rect 10977 14297 11011 14331
rect 15761 14297 15795 14331
rect 19717 14297 19751 14331
rect 19809 14297 19843 14331
rect 21925 14297 21959 14331
rect 3985 14229 4019 14263
rect 7665 14229 7699 14263
rect 18613 14229 18647 14263
rect 20913 14229 20947 14263
rect 22845 14229 22879 14263
rect 2145 14025 2179 14059
rect 2881 14025 2915 14059
rect 4721 14025 4755 14059
rect 5273 14025 5307 14059
rect 5733 14025 5767 14059
rect 7205 14025 7239 14059
rect 8217 14025 8251 14059
rect 11805 14025 11839 14059
rect 12909 14025 12943 14059
rect 13645 14025 13679 14059
rect 20453 14025 20487 14059
rect 22109 14025 22143 14059
rect 5641 13957 5675 13991
rect 6745 13957 6779 13991
rect 2421 13889 2455 13923
rect 3994 13889 4028 13923
rect 4261 13889 4295 13923
rect 8309 13889 8343 13923
rect 8861 13889 8895 13923
rect 11713 13889 11747 13923
rect 11897 13889 11931 13923
rect 14013 13889 14047 13923
rect 14381 13889 14415 13923
rect 15669 13889 15703 13923
rect 17049 13889 17083 13923
rect 17141 13889 17175 13923
rect 17325 13889 17359 13923
rect 17417 13889 17451 13923
rect 19809 13889 19843 13923
rect 19993 13889 20027 13923
rect 20085 13889 20119 13923
rect 20177 13889 20211 13923
rect 21097 13889 21131 13923
rect 21281 13889 21315 13923
rect 22017 13889 22051 13923
rect 2145 13821 2179 13855
rect 5825 13821 5859 13855
rect 11161 13821 11195 13855
rect 13921 13821 13955 13855
rect 14289 13821 14323 13855
rect 15025 13821 15059 13855
rect 21465 13821 21499 13855
rect 7113 13753 7147 13787
rect 16221 13753 16255 13787
rect 16865 13753 16899 13787
rect 22477 13753 22511 13787
rect 2329 13685 2363 13719
rect 22293 13685 22327 13719
rect 22385 13685 22419 13719
rect 22753 13685 22787 13719
rect 4169 13481 4203 13515
rect 6101 13481 6135 13515
rect 6837 13481 6871 13515
rect 7481 13481 7515 13515
rect 12817 13481 12851 13515
rect 14841 13481 14875 13515
rect 15301 13481 15335 13515
rect 16865 13481 16899 13515
rect 19993 13481 20027 13515
rect 22937 13481 22971 13515
rect 4721 13413 4755 13447
rect 8033 13413 8067 13447
rect 12725 13413 12759 13447
rect 1869 13345 1903 13379
rect 5273 13345 5307 13379
rect 11989 13345 12023 13379
rect 13553 13345 13587 13379
rect 19717 13345 19751 13379
rect 21189 13345 21223 13379
rect 1685 13277 1719 13311
rect 2053 13277 2087 13311
rect 2973 13277 3007 13311
rect 3249 13277 3283 13311
rect 4077 13277 4111 13311
rect 4261 13277 4295 13311
rect 5089 13277 5123 13311
rect 5181 13277 5215 13311
rect 7389 13277 7423 13311
rect 7573 13277 7607 13311
rect 8217 13277 8251 13311
rect 8309 13277 8343 13311
rect 8585 13277 8619 13311
rect 9137 13277 9171 13311
rect 10731 13277 10765 13311
rect 10885 13277 10919 13311
rect 11345 13277 11379 13311
rect 11621 13277 11655 13311
rect 11805 13277 11839 13311
rect 12541 13277 12575 13311
rect 12817 13277 12851 13311
rect 13277 13277 13311 13311
rect 14565 13277 14599 13311
rect 16405 13277 16439 13311
rect 16497 13277 16531 13311
rect 16681 13277 16715 13311
rect 19533 13277 19567 13311
rect 19625 13277 19659 13311
rect 19809 13277 19843 13311
rect 21005 13277 21039 13311
rect 21925 13277 21959 13311
rect 22293 13277 22327 13311
rect 3065 13209 3099 13243
rect 6285 13209 6319 13243
rect 8401 13209 8435 13243
rect 9965 13209 9999 13243
rect 14289 13209 14323 13243
rect 14473 13209 14507 13243
rect 1777 13141 1811 13175
rect 1961 13141 1995 13175
rect 3433 13141 3467 13175
rect 5917 13141 5951 13175
rect 6085 13141 6119 13175
rect 10517 13141 10551 13175
rect 14657 13141 14691 13175
rect 15945 13141 15979 13175
rect 4353 12937 4387 12971
rect 5381 12937 5415 12971
rect 12925 12937 12959 12971
rect 13553 12937 13587 12971
rect 13921 12937 13955 12971
rect 14749 12937 14783 12971
rect 18337 12937 18371 12971
rect 22017 12937 22051 12971
rect 5181 12869 5215 12903
rect 7021 12869 7055 12903
rect 11713 12869 11747 12903
rect 12725 12869 12759 12903
rect 14013 12869 14047 12903
rect 15485 12869 15519 12903
rect 22385 12869 22419 12903
rect 15715 12835 15749 12869
rect 2237 12801 2271 12835
rect 2789 12801 2823 12835
rect 2973 12801 3007 12835
rect 3065 12801 3099 12835
rect 4537 12801 4571 12835
rect 4721 12801 4755 12835
rect 6745 12801 6779 12835
rect 6837 12801 6871 12835
rect 9045 12801 9079 12835
rect 9229 12801 9263 12835
rect 10149 12801 10183 12835
rect 10241 12801 10275 12835
rect 10425 12801 10459 12835
rect 11897 12801 11931 12835
rect 11989 12801 12023 12835
rect 13829 12801 13863 12835
rect 14197 12801 14231 12835
rect 14289 12801 14323 12835
rect 14749 12801 14783 12835
rect 14933 12801 14967 12835
rect 16865 12801 16899 12835
rect 16958 12801 16992 12835
rect 17141 12801 17175 12835
rect 17233 12801 17267 12835
rect 17371 12801 17405 12835
rect 18613 12801 18647 12835
rect 22201 12801 22235 12835
rect 22477 12801 22511 12835
rect 10885 12733 10919 12767
rect 18521 12733 18555 12767
rect 18705 12733 18739 12767
rect 18797 12733 18831 12767
rect 2789 12665 2823 12699
rect 5549 12665 5583 12699
rect 7021 12665 7055 12699
rect 12173 12665 12207 12699
rect 13093 12665 13127 12699
rect 19349 12665 19383 12699
rect 2145 12597 2179 12631
rect 5365 12597 5399 12631
rect 9321 12597 9355 12631
rect 11713 12597 11747 12631
rect 12909 12597 12943 12631
rect 15669 12597 15703 12631
rect 15853 12597 15887 12631
rect 17509 12597 17543 12631
rect 22937 12597 22971 12631
rect 1777 12393 1811 12427
rect 1869 12393 1903 12427
rect 2421 12393 2455 12427
rect 2605 12393 2639 12427
rect 7573 12393 7607 12427
rect 8125 12393 8159 12427
rect 13645 12393 13679 12427
rect 18153 12393 18187 12427
rect 19717 12393 19751 12427
rect 4445 12325 4479 12359
rect 16037 12325 16071 12359
rect 1961 12257 1995 12291
rect 11897 12257 11931 12291
rect 14841 12257 14875 12291
rect 15761 12257 15795 12291
rect 17141 12257 17175 12291
rect 17693 12257 17727 12291
rect 17785 12257 17819 12291
rect 17877 12257 17911 12291
rect 21097 12257 21131 12291
rect 21741 12257 21775 12291
rect 1685 12189 1719 12223
rect 4077 12189 4111 12223
rect 4231 12189 4265 12223
rect 6929 12189 6963 12223
rect 7389 12189 7423 12223
rect 7573 12189 7607 12223
rect 8033 12189 8067 12223
rect 8309 12189 8343 12223
rect 8401 12189 8435 12223
rect 9137 12189 9171 12223
rect 9689 12189 9723 12223
rect 11989 12189 12023 12223
rect 12173 12189 12207 12223
rect 13093 12189 13127 12223
rect 13277 12189 13311 12223
rect 13461 12189 13495 12223
rect 14289 12189 14323 12223
rect 14473 12189 14507 12223
rect 15577 12189 15611 12223
rect 15669 12189 15703 12223
rect 15853 12189 15887 12223
rect 16497 12189 16531 12223
rect 16681 12189 16715 12223
rect 16773 12189 16807 12223
rect 16865 12189 16899 12223
rect 17969 12189 18003 12223
rect 19901 12189 19935 12223
rect 19993 12189 20027 12223
rect 20085 12189 20119 12223
rect 20177 12189 20211 12223
rect 20361 12189 20395 12223
rect 21281 12189 21315 12223
rect 21465 12189 21499 12223
rect 21583 12189 21617 12223
rect 22293 12189 22327 12223
rect 22385 12189 22419 12223
rect 23029 12189 23063 12223
rect 23213 12189 23247 12223
rect 2789 12121 2823 12155
rect 10701 12121 10735 12155
rect 10885 12121 10919 12155
rect 12633 12121 12667 12155
rect 13369 12121 13403 12155
rect 21373 12121 21407 12155
rect 22569 12121 22603 12155
rect 2579 12053 2613 12087
rect 4905 12053 4939 12087
rect 6377 12053 6411 12087
rect 8585 12053 8619 12087
rect 9229 12053 9263 12087
rect 10517 12053 10551 12087
rect 23121 12053 23155 12087
rect 4353 11849 4387 11883
rect 6561 11849 6595 11883
rect 8585 11849 8619 11883
rect 12633 11849 12667 11883
rect 15209 11849 15243 11883
rect 15577 11849 15611 11883
rect 17417 11849 17451 11883
rect 20729 11849 20763 11883
rect 22201 11849 22235 11883
rect 5181 11781 5215 11815
rect 6837 11781 6871 11815
rect 8953 11781 8987 11815
rect 13553 11781 13587 11815
rect 13921 11781 13955 11815
rect 14381 11781 14415 11815
rect 15301 11781 15335 11815
rect 22753 11781 22787 11815
rect 3939 11713 3973 11747
rect 5365 11713 5399 11747
rect 5457 11713 5491 11747
rect 5549 11713 5583 11747
rect 5687 11713 5721 11747
rect 6745 11713 6779 11747
rect 6929 11713 6963 11747
rect 7047 11713 7081 11747
rect 8769 11713 8803 11747
rect 8861 11713 8895 11747
rect 9071 11713 9105 11747
rect 10057 11713 10091 11747
rect 10609 11713 10643 11747
rect 13461 11713 13495 11747
rect 15393 11713 15427 11747
rect 16865 11713 16899 11747
rect 16957 11713 16991 11747
rect 17141 11713 17175 11747
rect 17233 11713 17267 11747
rect 20913 11713 20947 11747
rect 21097 11713 21131 11747
rect 22109 11713 22143 11747
rect 22293 11713 22327 11747
rect 3709 11645 3743 11679
rect 3801 11645 3835 11679
rect 4077 11645 4111 11679
rect 4169 11645 4203 11679
rect 5825 11645 5859 11679
rect 7205 11645 7239 11679
rect 9229 11645 9263 11679
rect 9965 11645 9999 11679
rect 13369 11645 13403 11679
rect 17877 11645 17911 11679
rect 8033 11577 8067 11611
rect 15025 11577 15059 11611
rect 19349 11577 19383 11611
rect 9781 11509 9815 11543
rect 16221 11509 16255 11543
rect 18521 11509 18555 11543
rect 20913 11509 20947 11543
rect 1869 11305 1903 11339
rect 11805 11305 11839 11339
rect 12633 11305 12667 11339
rect 13185 11305 13219 11339
rect 14381 11305 14415 11339
rect 14841 11305 14875 11339
rect 16865 11305 16899 11339
rect 18521 11305 18555 11339
rect 20085 11305 20119 11339
rect 22937 11305 22971 11339
rect 4537 11237 4571 11271
rect 4261 11169 4295 11203
rect 9321 11169 9355 11203
rect 15945 11169 15979 11203
rect 18429 11169 18463 11203
rect 18613 11169 18647 11203
rect 21925 11169 21959 11203
rect 1593 11101 1627 11135
rect 2145 11101 2179 11135
rect 2697 11101 2731 11135
rect 2973 11101 3007 11135
rect 4169 11101 4203 11135
rect 7481 11101 7515 11135
rect 8217 11101 8251 11135
rect 9597 11101 9631 11135
rect 12081 11101 12115 11135
rect 15117 11101 15151 11135
rect 15209 11101 15243 11135
rect 15301 11101 15335 11135
rect 15485 11101 15519 11135
rect 16129 11101 16163 11135
rect 16313 11101 16347 11135
rect 17049 11101 17083 11135
rect 17141 11101 17175 11135
rect 17325 11101 17359 11135
rect 17417 11101 17451 11135
rect 18705 11101 18739 11135
rect 19717 11101 19751 11135
rect 19809 11101 19843 11135
rect 22385 11101 22419 11135
rect 22477 11101 22511 11135
rect 22661 11101 22695 11135
rect 22753 11101 22787 11135
rect 10149 11033 10183 11067
rect 11621 11033 11655 11067
rect 11805 11033 11839 11067
rect 13737 11033 13771 11067
rect 19533 11033 19567 11067
rect 19901 11033 19935 11067
rect 17877 10965 17911 10999
rect 1777 10761 1811 10795
rect 5457 10761 5491 10795
rect 6745 10761 6779 10795
rect 8953 10761 8987 10795
rect 12817 10761 12851 10795
rect 14749 10761 14783 10795
rect 18337 10761 18371 10795
rect 21373 10761 21407 10795
rect 2237 10693 2271 10727
rect 3065 10693 3099 10727
rect 14381 10693 14415 10727
rect 14473 10693 14507 10727
rect 17509 10693 17543 10727
rect 1961 10625 1995 10659
rect 2697 10625 2731 10659
rect 2973 10625 3007 10659
rect 4537 10625 4571 10659
rect 5641 10625 5675 10659
rect 5733 10625 5767 10659
rect 6929 10625 6963 10659
rect 7113 10625 7147 10659
rect 7757 10625 7791 10659
rect 7941 10625 7975 10659
rect 8953 10625 8987 10659
rect 9137 10625 9171 10659
rect 9873 10625 9907 10659
rect 11897 10625 11931 10659
rect 11989 10625 12023 10659
rect 12081 10625 12115 10659
rect 12265 10625 12299 10659
rect 14105 10625 14139 10659
rect 14253 10625 14287 10659
rect 14570 10625 14604 10659
rect 15577 10625 15611 10659
rect 15669 10625 15703 10659
rect 15853 10625 15887 10659
rect 15945 10625 15979 10659
rect 16865 10625 16899 10659
rect 17049 10625 17083 10659
rect 17141 10625 17175 10659
rect 17234 10625 17268 10659
rect 18521 10625 18555 10659
rect 18613 10625 18647 10659
rect 18889 10625 18923 10659
rect 22385 10625 22419 10659
rect 2053 10557 2087 10591
rect 4261 10557 4295 10591
rect 5825 10557 5859 10591
rect 5917 10557 5951 10591
rect 7021 10557 7055 10591
rect 7205 10557 7239 10591
rect 9689 10557 9723 10591
rect 13093 10557 13127 10591
rect 22109 10557 22143 10591
rect 22201 10557 22235 10591
rect 22293 10557 22327 10591
rect 11713 10489 11747 10523
rect 13185 10489 13219 10523
rect 13645 10489 13679 10523
rect 2237 10421 2271 10455
rect 3617 10421 3651 10455
rect 7757 10421 7791 10455
rect 10057 10421 10091 10455
rect 10609 10421 10643 10455
rect 11069 10421 11103 10455
rect 13277 10421 13311 10455
rect 15393 10421 15427 10455
rect 18797 10421 18831 10455
rect 19441 10421 19475 10455
rect 22569 10421 22603 10455
rect 4537 10217 4571 10251
rect 6193 10217 6227 10251
rect 8585 10217 8619 10251
rect 15485 10217 15519 10251
rect 15669 10217 15703 10251
rect 21649 10217 21683 10251
rect 3249 10149 3283 10183
rect 5457 10149 5491 10183
rect 13277 10149 13311 10183
rect 17417 10149 17451 10183
rect 19901 10149 19935 10183
rect 2237 10081 2271 10115
rect 9689 10081 9723 10115
rect 15025 10081 15059 10115
rect 1961 10013 1995 10047
rect 2145 10013 2179 10047
rect 2973 10013 3007 10047
rect 3249 10013 3283 10047
rect 4077 10013 4111 10047
rect 4169 10013 4203 10047
rect 4261 10013 4295 10047
rect 4353 10013 4387 10047
rect 4997 10013 5031 10047
rect 6929 10013 6963 10047
rect 7389 10013 7423 10047
rect 9229 10013 9263 10047
rect 11713 10013 11747 10047
rect 11989 10013 12023 10047
rect 14289 10013 14323 10047
rect 14381 10013 14415 10047
rect 14565 10013 14599 10047
rect 16405 10013 16439 10047
rect 16589 10013 16623 10047
rect 18061 10013 18095 10047
rect 18245 10013 18279 10047
rect 18337 10013 18371 10047
rect 18429 10013 18463 10047
rect 18521 10013 18555 10047
rect 20085 10013 20119 10047
rect 20545 10013 20579 10047
rect 21005 10013 21039 10047
rect 21189 10013 21223 10047
rect 21281 10013 21315 10047
rect 21373 10013 21407 10047
rect 6009 9945 6043 9979
rect 6209 9945 6243 9979
rect 15637 9945 15671 9979
rect 15853 9945 15887 9979
rect 16957 9945 16991 9979
rect 18705 9945 18739 9979
rect 6377 9877 6411 9911
rect 9413 9877 9447 9911
rect 10241 9877 10275 9911
rect 2237 9673 2271 9707
rect 3157 9673 3191 9707
rect 7021 9673 7055 9707
rect 8217 9673 8251 9707
rect 14289 9673 14323 9707
rect 4905 9605 4939 9639
rect 5181 9605 5215 9639
rect 8309 9605 8343 9639
rect 13737 9605 13771 9639
rect 15945 9605 15979 9639
rect 17601 9605 17635 9639
rect 18061 9605 18095 9639
rect 20361 9605 20395 9639
rect 2148 9537 2182 9571
rect 2421 9537 2455 9571
rect 3065 9537 3099 9571
rect 3249 9537 3283 9571
rect 3893 9537 3927 9571
rect 5089 9537 5123 9571
rect 5273 9537 5307 9571
rect 5411 9537 5445 9571
rect 7205 9537 7239 9571
rect 7297 9537 7331 9571
rect 7425 9537 7459 9571
rect 9137 9537 9171 9571
rect 9321 9537 9355 9571
rect 9413 9537 9447 9571
rect 9505 9537 9539 9571
rect 10241 9537 10275 9571
rect 11713 9537 11747 9571
rect 11897 9537 11931 9571
rect 12909 9537 12943 9571
rect 13093 9537 13127 9571
rect 13277 9537 13311 9571
rect 14289 9537 14323 9571
rect 14473 9537 14507 9571
rect 15025 9537 15059 9571
rect 15117 9537 15151 9571
rect 16865 9537 16899 9571
rect 18245 9537 18279 9571
rect 18429 9537 18463 9571
rect 19073 9537 19107 9571
rect 19349 9537 19383 9571
rect 20085 9537 20119 9571
rect 20269 9537 20303 9571
rect 20821 9537 20855 9571
rect 22017 9537 22051 9571
rect 22109 9537 22143 9571
rect 22293 9537 22327 9571
rect 5549 9469 5583 9503
rect 8033 9469 8067 9503
rect 9781 9469 9815 9503
rect 10333 9469 10367 9503
rect 17233 9469 17267 9503
rect 19165 9469 19199 9503
rect 8677 9401 8711 9435
rect 15393 9401 15427 9435
rect 19533 9401 19567 9435
rect 1685 9333 1719 9367
rect 2605 9333 2639 9367
rect 4353 9333 4387 9367
rect 10333 9333 10367 9367
rect 10609 9333 10643 9367
rect 11805 9333 11839 9367
rect 15025 9333 15059 9367
rect 17003 9333 17037 9367
rect 17141 9333 17175 9367
rect 22477 9333 22511 9367
rect 5181 9129 5215 9163
rect 7021 9129 7055 9163
rect 20085 9129 20119 9163
rect 22109 9129 22143 9163
rect 5273 9061 5307 9095
rect 11529 9061 11563 9095
rect 18797 9061 18831 9095
rect 19533 9061 19567 9095
rect 23213 9061 23247 9095
rect 6745 8993 6779 9027
rect 6837 8993 6871 9027
rect 11069 8993 11103 9027
rect 14565 8993 14599 9027
rect 15485 8993 15519 9027
rect 16865 8993 16899 9027
rect 21281 8993 21315 9027
rect 1869 8925 1903 8959
rect 2053 8925 2087 8959
rect 2973 8925 3007 8959
rect 3985 8925 4019 8959
rect 5365 8925 5399 8959
rect 6561 8925 6595 8959
rect 6653 8925 6687 8959
rect 9137 8925 9171 8959
rect 10057 8925 10091 8959
rect 11713 8925 11747 8959
rect 11805 8925 11839 8959
rect 11989 8925 12023 8959
rect 12081 8925 12115 8959
rect 12541 8925 12575 8959
rect 13185 8925 13219 8959
rect 13277 8925 13311 8959
rect 13461 8925 13495 8959
rect 13553 8925 13587 8959
rect 14473 8925 14507 8959
rect 14749 8925 14783 8959
rect 14933 8925 14967 8959
rect 16589 8925 16623 8959
rect 18153 8925 18187 8959
rect 20269 8925 20303 8959
rect 20361 8925 20395 8959
rect 20545 8925 20579 8959
rect 20637 8925 20671 8959
rect 21189 8925 21223 8959
rect 21373 8925 21407 8959
rect 21465 8925 21499 8959
rect 22385 8925 22419 8959
rect 22477 8925 22511 8959
rect 22569 8925 22603 8959
rect 22753 8925 22787 8959
rect 2697 8857 2731 8891
rect 4261 8857 4295 8891
rect 5089 8857 5123 8891
rect 9597 8857 9631 8891
rect 1961 8789 1995 8823
rect 12633 8789 12667 8823
rect 13737 8789 13771 8823
rect 16037 8789 16071 8823
rect 17877 8789 17911 8823
rect 21649 8789 21683 8823
rect 3525 8585 3559 8619
rect 9321 8585 9355 8619
rect 11713 8585 11747 8619
rect 13093 8585 13127 8619
rect 15485 8585 15519 8619
rect 15577 8585 15611 8619
rect 16221 8585 16255 8619
rect 16865 8585 16899 8619
rect 19349 8585 19383 8619
rect 20085 8585 20119 8619
rect 22017 8585 22051 8619
rect 4261 8517 4295 8551
rect 5181 8517 5215 8551
rect 6745 8517 6779 8551
rect 7297 8517 7331 8551
rect 12357 8517 12391 8551
rect 15209 8517 15243 8551
rect 15761 8517 15795 8551
rect 20453 8517 20487 8551
rect 21005 8517 21039 8551
rect 2329 8449 2363 8483
rect 2421 8449 2455 8483
rect 3065 8449 3099 8483
rect 3341 8449 3375 8483
rect 4169 8449 4203 8483
rect 4629 8449 4663 8483
rect 6857 8449 6891 8483
rect 7941 8449 7975 8483
rect 8401 8449 8435 8483
rect 9873 8449 9907 8483
rect 10241 8449 10275 8483
rect 10977 8449 11011 8483
rect 12265 8449 12299 8483
rect 12541 8449 12575 8483
rect 13553 8449 13587 8483
rect 13737 8449 13771 8483
rect 14013 8449 14047 8483
rect 14105 8449 14139 8483
rect 15393 8449 15427 8483
rect 17417 8449 17451 8483
rect 17601 8449 17635 8483
rect 18153 8449 18187 8483
rect 18337 8449 18371 8483
rect 19257 8449 19291 8483
rect 19441 8449 19475 8483
rect 20269 8449 20303 8483
rect 20545 8449 20579 8483
rect 22201 8449 22235 8483
rect 22293 8449 22327 8483
rect 22477 8449 22511 8483
rect 22661 8449 22695 8483
rect 3249 8381 3283 8415
rect 8033 8381 8067 8415
rect 10425 8381 10459 8415
rect 11069 8381 11103 8415
rect 14749 8381 14783 8415
rect 22385 8381 22419 8415
rect 2605 8313 2639 8347
rect 5733 8313 5767 8347
rect 9965 8313 9999 8347
rect 12541 8313 12575 8347
rect 18613 8313 18647 8347
rect 2145 8245 2179 8279
rect 3065 8245 3099 8279
rect 6561 8245 6595 8279
rect 7757 8245 7791 8279
rect 8309 8245 8343 8279
rect 2237 8041 2271 8075
rect 4629 8041 4663 8075
rect 7757 8041 7791 8075
rect 8125 8041 8159 8075
rect 11621 8041 11655 8075
rect 12633 8041 12667 8075
rect 12817 8041 12851 8075
rect 13737 8041 13771 8075
rect 14565 8041 14599 8075
rect 15853 8041 15887 8075
rect 16037 8041 16071 8075
rect 18429 8041 18463 8075
rect 18613 8041 18647 8075
rect 20821 8041 20855 8075
rect 22753 8041 22787 8075
rect 4077 7973 4111 8007
rect 11069 7973 11103 8007
rect 4813 7905 4847 7939
rect 7849 7905 7883 7939
rect 11875 7905 11909 7939
rect 13001 7905 13035 7939
rect 16497 7905 16531 7939
rect 17877 7905 17911 7939
rect 2145 7837 2179 7871
rect 2329 7837 2363 7871
rect 3249 7837 3283 7871
rect 4537 7837 4571 7871
rect 5273 7837 5307 7871
rect 6285 7837 6319 7871
rect 6929 7837 6963 7871
rect 7757 7837 7791 7871
rect 9137 7837 9171 7871
rect 9413 7837 9447 7871
rect 9505 7837 9539 7871
rect 10333 7837 10367 7871
rect 10425 7837 10459 7871
rect 10701 7837 10735 7871
rect 10793 7837 10827 7871
rect 11792 7837 11826 7871
rect 11989 7837 12023 7871
rect 12081 7837 12115 7871
rect 12817 7837 12851 7871
rect 14473 7837 14507 7871
rect 14657 7837 14691 7871
rect 16865 7837 16899 7871
rect 17049 7837 17083 7871
rect 17233 7837 17267 7871
rect 17417 7837 17451 7871
rect 19441 7837 19475 7871
rect 19625 7837 19659 7871
rect 20085 7837 20119 7871
rect 20821 7837 20855 7871
rect 21097 7837 21131 7871
rect 22109 7837 22143 7871
rect 18567 7803 18601 7837
rect 2973 7769 3007 7803
rect 5549 7769 5583 7803
rect 6745 7769 6779 7803
rect 9321 7769 9355 7803
rect 13093 7769 13127 7803
rect 15669 7769 15703 7803
rect 18797 7769 18831 7803
rect 21005 7769 21039 7803
rect 4813 7701 4847 7735
rect 9689 7701 9723 7735
rect 10609 7701 10643 7735
rect 15117 7701 15151 7735
rect 15869 7701 15903 7735
rect 22201 7701 22235 7735
rect 8401 7497 8435 7531
rect 9505 7497 9539 7531
rect 10241 7497 10275 7531
rect 12081 7497 12115 7531
rect 15117 7497 15151 7531
rect 15209 7497 15243 7531
rect 21465 7497 21499 7531
rect 11161 7429 11195 7463
rect 14381 7429 14415 7463
rect 14933 7429 14967 7463
rect 15485 7429 15519 7463
rect 17601 7429 17635 7463
rect 1960 7361 1994 7395
rect 2053 7361 2087 7395
rect 2789 7361 2823 7395
rect 2973 7361 3007 7395
rect 3893 7361 3927 7395
rect 4813 7361 4847 7395
rect 5457 7361 5491 7395
rect 5549 7361 5583 7395
rect 5917 7361 5951 7395
rect 7021 7361 7055 7395
rect 8033 7361 8067 7395
rect 8125 7361 8159 7395
rect 8861 7361 8895 7395
rect 9045 7361 9079 7395
rect 9137 7361 9171 7395
rect 9229 7361 9263 7395
rect 10149 7361 10183 7395
rect 10333 7361 10367 7395
rect 11989 7361 12023 7395
rect 14289 7361 14323 7395
rect 15301 7361 15335 7395
rect 16865 7361 16899 7395
rect 17012 7361 17046 7395
rect 18797 7361 18831 7395
rect 19441 7361 19475 7395
rect 22385 7361 22419 7395
rect 22569 7361 22603 7395
rect 22661 7361 22695 7395
rect 22753 7361 22787 7395
rect 2605 7293 2639 7327
rect 3617 7293 3651 7327
rect 4629 7293 4663 7327
rect 6929 7293 6963 7327
rect 17233 7293 17267 7327
rect 20085 7293 20119 7327
rect 17141 7225 17175 7259
rect 1869 7157 1903 7191
rect 5273 7157 5307 7191
rect 5825 7157 5859 7191
rect 6653 7157 6687 7191
rect 7021 7157 7055 7191
rect 8125 7157 8159 7191
rect 12725 7157 12759 7191
rect 15945 7157 15979 7191
rect 23029 7157 23063 7191
rect 2329 6953 2363 6987
rect 8585 6953 8619 6987
rect 13277 6953 13311 6987
rect 16681 6953 16715 6987
rect 13645 6885 13679 6919
rect 4721 6817 4755 6851
rect 6101 6817 6135 6851
rect 7481 6817 7515 6851
rect 9965 6817 9999 6851
rect 10241 6817 10275 6851
rect 10333 6817 10367 6851
rect 10425 6817 10459 6851
rect 17325 6817 17359 6851
rect 17785 6817 17819 6851
rect 19901 6817 19935 6851
rect 21741 6817 21775 6851
rect 22201 6817 22235 6851
rect 22661 6817 22695 6851
rect 1961 6749 1995 6783
rect 2329 6749 2363 6783
rect 3065 6749 3099 6783
rect 3249 6749 3283 6783
rect 3341 6749 3375 6783
rect 4261 6749 4295 6783
rect 5641 6749 5675 6783
rect 5825 6749 5859 6783
rect 6193 6749 6227 6783
rect 7941 6749 7975 6783
rect 8034 6749 8068 6783
rect 8309 6749 8343 6783
rect 8406 6749 8440 6783
rect 10149 6749 10183 6783
rect 11621 6749 11655 6783
rect 11897 6749 11931 6783
rect 13461 6749 13495 6783
rect 13737 6749 13771 6783
rect 15117 6749 15151 6783
rect 15301 6749 15335 6783
rect 17509 6749 17543 6783
rect 18889 6749 18923 6783
rect 19441 6749 19475 6783
rect 19625 6749 19659 6783
rect 19993 6749 20027 6783
rect 21097 6749 21131 6783
rect 21281 6749 21315 6783
rect 21373 6749 21407 6783
rect 21465 6749 21499 6783
rect 22385 6749 22419 6783
rect 22477 6749 22511 6783
rect 22753 6749 22787 6783
rect 4169 6681 4203 6715
rect 4629 6681 4663 6715
rect 6837 6681 6871 6715
rect 8217 6681 8251 6715
rect 18337 6681 18371 6715
rect 2513 6613 2547 6647
rect 9505 6613 9539 6647
rect 11437 6613 11471 6647
rect 11805 6613 11839 6647
rect 15209 6613 15243 6647
rect 20361 6613 20395 6647
rect 3433 6409 3467 6443
rect 18981 6409 19015 6443
rect 21465 6409 21499 6443
rect 23029 6409 23063 6443
rect 12265 6341 12299 6375
rect 12475 6341 12509 6375
rect 13185 6341 13219 6375
rect 18061 6341 18095 6375
rect 20453 6341 20487 6375
rect 22937 6341 22971 6375
rect 2237 6273 2271 6307
rect 2421 6273 2455 6307
rect 2697 6273 2731 6307
rect 2973 6273 3007 6307
rect 3065 6273 3099 6307
rect 4169 6273 4203 6307
rect 4629 6273 4663 6307
rect 4905 6273 4939 6307
rect 5365 6273 5399 6307
rect 6561 6273 6595 6307
rect 6745 6273 6779 6307
rect 7389 6273 7423 6307
rect 7941 6273 7975 6307
rect 8309 6273 8343 6307
rect 8401 6273 8435 6307
rect 8953 6273 8987 6307
rect 12173 6273 12207 6307
rect 12357 6273 12391 6307
rect 12633 6273 12667 6307
rect 13829 6273 13863 6307
rect 15485 6273 15519 6307
rect 16865 6273 16899 6307
rect 17049 6273 17083 6307
rect 17417 6273 17451 6307
rect 18521 6273 18555 6307
rect 18797 6273 18831 6307
rect 19717 6273 19751 6307
rect 19993 6273 20027 6307
rect 21097 6273 21131 6307
rect 21281 6273 21315 6307
rect 22017 6273 22051 6307
rect 22293 6273 22327 6307
rect 23213 6273 23247 6307
rect 9137 6205 9171 6239
rect 14105 6205 14139 6239
rect 14749 6205 14783 6239
rect 15393 6205 15427 6239
rect 15761 6205 15795 6239
rect 15853 6205 15887 6239
rect 17325 6205 17359 6239
rect 19809 6205 19843 6239
rect 21005 6205 21039 6239
rect 23305 6205 23339 6239
rect 4721 6137 4755 6171
rect 11989 6137 12023 6171
rect 18613 6137 18647 6171
rect 4077 6069 4111 6103
rect 6009 6069 6043 6103
rect 6561 6069 6595 6103
rect 13645 6069 13679 6103
rect 14013 6069 14047 6103
rect 15209 6069 15243 6103
rect 23121 6069 23155 6103
rect 2145 5865 2179 5899
rect 3985 5865 4019 5899
rect 9229 5865 9263 5899
rect 11713 5865 11747 5899
rect 13369 5865 13403 5899
rect 14841 5865 14875 5899
rect 16405 5865 16439 5899
rect 21281 5865 21315 5899
rect 21925 5865 21959 5899
rect 3341 5797 3375 5831
rect 12357 5797 12391 5831
rect 20177 5797 20211 5831
rect 2329 5729 2363 5763
rect 8033 5729 8067 5763
rect 8125 5729 8159 5763
rect 8217 5729 8251 5763
rect 8401 5729 8435 5763
rect 10149 5729 10183 5763
rect 12725 5729 12759 5763
rect 12817 5729 12851 5763
rect 17509 5729 17543 5763
rect 18245 5729 18279 5763
rect 19533 5729 19567 5763
rect 20637 5729 20671 5763
rect 22293 5729 22327 5763
rect 22937 5729 22971 5763
rect 2421 5661 2455 5695
rect 3249 5661 3283 5695
rect 4169 5661 4203 5695
rect 4813 5661 4847 5695
rect 5181 5661 5215 5695
rect 6009 5661 6043 5695
rect 7021 5661 7055 5695
rect 7941 5661 7975 5695
rect 10333 5661 10367 5695
rect 10609 5661 10643 5695
rect 11069 5661 11103 5695
rect 11253 5661 11287 5695
rect 11345 5661 11379 5695
rect 11437 5661 11471 5695
rect 12541 5661 12575 5695
rect 12633 5661 12667 5695
rect 13369 5661 13403 5695
rect 13553 5661 13587 5695
rect 15117 5661 15151 5695
rect 15577 5661 15611 5695
rect 16589 5661 16623 5695
rect 17049 5661 17083 5695
rect 17233 5661 17267 5695
rect 17601 5661 17635 5695
rect 20085 5661 20119 5695
rect 20361 5661 20395 5695
rect 22109 5661 22143 5695
rect 22753 5661 22787 5695
rect 2145 5593 2179 5627
rect 4353 5593 4387 5627
rect 6653 5593 6687 5627
rect 7205 5593 7239 5627
rect 15025 5593 15059 5627
rect 1685 5525 1719 5559
rect 2605 5525 2639 5559
rect 5759 5525 5793 5559
rect 6837 5525 6871 5559
rect 6929 5525 6963 5559
rect 10517 5525 10551 5559
rect 2605 5321 2639 5355
rect 12449 5321 12483 5355
rect 14381 5321 14415 5355
rect 15025 5321 15059 5355
rect 16221 5321 16255 5355
rect 17141 5321 17175 5355
rect 19257 5321 19291 5355
rect 20453 5321 20487 5355
rect 21189 5321 21223 5355
rect 22293 5321 22327 5355
rect 10977 5253 11011 5287
rect 15301 5253 15335 5287
rect 15393 5253 15427 5287
rect 17293 5253 17327 5287
rect 17509 5253 17543 5287
rect 23029 5253 23063 5287
rect 2053 5185 2087 5219
rect 2145 5185 2179 5219
rect 2329 5185 2363 5219
rect 2421 5185 2455 5219
rect 3249 5185 3283 5219
rect 4169 5185 4203 5219
rect 5549 5185 5583 5219
rect 6561 5185 6595 5219
rect 6745 5185 6779 5219
rect 8033 5185 8067 5219
rect 8677 5185 8711 5219
rect 9413 5185 9447 5219
rect 9689 5185 9723 5219
rect 9781 5185 9815 5219
rect 9965 5185 9999 5219
rect 10425 5185 10459 5219
rect 10517 5185 10551 5219
rect 10701 5185 10735 5219
rect 10793 5185 10827 5219
rect 12633 5185 12667 5219
rect 12725 5185 12759 5219
rect 12817 5185 12851 5219
rect 13001 5185 13035 5219
rect 15163 5185 15197 5219
rect 15576 5185 15610 5219
rect 15669 5185 15703 5219
rect 18153 5185 18187 5219
rect 18245 5185 18279 5219
rect 18429 5185 18463 5219
rect 19625 5185 19659 5219
rect 20545 5185 20579 5219
rect 21097 5185 21131 5219
rect 21281 5185 21315 5219
rect 22753 5185 22787 5219
rect 3525 5117 3559 5151
rect 4997 5117 5031 5151
rect 5733 5117 5767 5151
rect 7757 5117 7791 5151
rect 9597 5117 9631 5151
rect 19717 5117 19751 5151
rect 8493 5049 8527 5083
rect 18613 5049 18647 5083
rect 6653 4981 6687 5015
rect 9229 4981 9263 5015
rect 13553 4981 13587 5015
rect 17325 4981 17359 5015
rect 5733 4777 5767 4811
rect 9413 4777 9447 4811
rect 11161 4777 11195 4811
rect 12081 4777 12115 4811
rect 15025 4777 15059 4811
rect 15577 4777 15611 4811
rect 17325 4777 17359 4811
rect 19809 4777 19843 4811
rect 20269 4777 20303 4811
rect 20821 4777 20855 4811
rect 16405 4709 16439 4743
rect 4813 4641 4847 4675
rect 9597 4641 9631 4675
rect 10057 4641 10091 4675
rect 18889 4641 18923 4675
rect 22661 4641 22695 4675
rect 2421 4573 2455 4607
rect 3341 4573 3375 4607
rect 4261 4573 4295 4607
rect 4353 4573 4387 4607
rect 5365 4573 5399 4607
rect 5549 4573 5583 4607
rect 6929 4573 6963 4607
rect 7021 4573 7055 4607
rect 7297 4573 7331 4607
rect 7481 4573 7515 4607
rect 7941 4573 7975 4607
rect 8125 4573 8159 4607
rect 9689 4573 9723 4607
rect 12265 4573 12299 4607
rect 12541 4573 12575 4607
rect 14565 4573 14599 4607
rect 14841 4573 14875 4607
rect 15761 4573 15795 4607
rect 15945 4573 15979 4607
rect 17509 4573 17543 4607
rect 17877 4573 17911 4607
rect 19625 4573 19659 4607
rect 22753 4573 22787 4607
rect 22937 4573 22971 4607
rect 2145 4505 2179 4539
rect 3065 4505 3099 4539
rect 4077 4505 4111 4539
rect 4445 4505 4479 4539
rect 5273 4505 5307 4539
rect 6285 4505 6319 4539
rect 9965 4505 9999 4539
rect 12449 4505 12483 4539
rect 17601 4505 17635 4539
rect 17693 4505 17727 4539
rect 19441 4505 19475 4539
rect 8033 4437 8067 4471
rect 10609 4437 10643 4471
rect 14657 4437 14691 4471
rect 6745 4233 6779 4267
rect 6837 4233 6871 4267
rect 13645 4233 13679 4267
rect 17969 4233 18003 4267
rect 22661 4233 22695 4267
rect 3709 4165 3743 4199
rect 6653 4165 6687 4199
rect 1961 4097 1995 4131
rect 2053 4097 2087 4131
rect 2145 4097 2179 4131
rect 2789 4097 2823 4131
rect 3893 4097 3927 4131
rect 4445 4097 4479 4131
rect 4629 4097 4663 4131
rect 5457 4097 5491 4131
rect 5641 4097 5675 4131
rect 6009 4097 6043 4131
rect 7389 4097 7423 4131
rect 8125 4097 8159 4131
rect 8309 4097 8343 4131
rect 8769 4097 8803 4131
rect 9045 4097 9079 4131
rect 9229 4097 9263 4131
rect 14289 4097 14323 4131
rect 15209 4097 15243 4131
rect 15945 4097 15979 4131
rect 16037 4097 16071 4131
rect 16129 4100 16163 4134
rect 16313 4097 16347 4131
rect 16865 4097 16899 4131
rect 18521 4097 18555 4131
rect 18981 4097 19015 4131
rect 19165 4097 19199 4131
rect 19349 4097 19383 4131
rect 19533 4097 19567 4131
rect 19809 4097 19843 4131
rect 22569 4097 22603 4131
rect 22753 4097 22787 4131
rect 2697 4029 2731 4063
rect 4905 4029 4939 4063
rect 7205 4029 7239 4063
rect 1777 3893 1811 3927
rect 2973 3893 3007 3927
rect 8125 3893 8159 3927
rect 8861 3893 8895 3927
rect 9689 3893 9723 3927
rect 10333 3893 10367 3927
rect 10977 3893 11011 3927
rect 11713 3893 11747 3927
rect 12265 3893 12299 3927
rect 15669 3893 15703 3927
rect 2513 3689 2547 3723
rect 8585 3689 8619 3723
rect 13093 3689 13127 3723
rect 17969 3689 18003 3723
rect 3065 3621 3099 3655
rect 6101 3621 6135 3655
rect 10885 3621 10919 3655
rect 2605 3553 2639 3587
rect 6745 3553 6779 3587
rect 7941 3553 7975 3587
rect 10425 3553 10459 3587
rect 11161 3553 11195 3587
rect 12817 3553 12851 3587
rect 14933 3553 14967 3587
rect 20085 3553 20119 3587
rect 22385 3553 22419 3587
rect 2329 3485 2363 3519
rect 3340 3485 3374 3519
rect 3426 3485 3460 3519
rect 4445 3485 4479 3519
rect 4905 3485 4939 3519
rect 5181 3485 5215 3519
rect 5273 3485 5307 3519
rect 5641 3485 5675 3519
rect 6561 3485 6595 3519
rect 7849 3485 7883 3519
rect 8033 3485 8067 3519
rect 9321 3485 9355 3519
rect 9965 3485 9999 3519
rect 10241 3485 10275 3519
rect 11069 3485 11103 3519
rect 11529 3485 11563 3519
rect 12909 3485 12943 3519
rect 13553 3485 13587 3519
rect 13737 3485 13771 3519
rect 14289 3485 14323 3519
rect 14473 3485 14507 3519
rect 15577 3485 15611 3519
rect 16221 3485 16255 3519
rect 18889 3485 18923 3519
rect 19809 3485 19843 3519
rect 22845 3485 22879 3519
rect 1685 3417 1719 3451
rect 4169 3417 4203 3451
rect 11437 3417 11471 3451
rect 14381 3417 14415 3451
rect 2145 3349 2179 3383
rect 10057 3349 10091 3383
rect 11345 3349 11379 3383
rect 12449 3349 12483 3383
rect 13645 3349 13679 3383
rect 16865 3349 16899 3383
rect 17417 3349 17451 3383
rect 19515 3349 19549 3383
rect 19993 3349 20027 3383
rect 20637 3349 20671 3383
rect 5457 3145 5491 3179
rect 9597 3145 9631 3179
rect 11897 3145 11931 3179
rect 13185 3145 13219 3179
rect 16865 3145 16899 3179
rect 20821 3145 20855 3179
rect 4445 3077 4479 3111
rect 10149 3077 10183 3111
rect 16037 3077 16071 3111
rect 20637 3077 20671 3111
rect 2237 3009 2271 3043
rect 2420 3009 2454 3043
rect 2513 3009 2547 3043
rect 2789 3009 2823 3043
rect 3801 3009 3835 3043
rect 3985 3009 4019 3043
rect 4077 3009 4111 3043
rect 4261 3009 4295 3043
rect 5089 3009 5123 3043
rect 5641 3009 5675 3043
rect 6561 3009 6595 3043
rect 7389 3009 7423 3043
rect 8401 3009 8435 3043
rect 8861 3009 8895 3043
rect 9045 3009 9079 3043
rect 9321 3009 9355 3043
rect 12265 3009 12299 3043
rect 13277 3009 13311 3043
rect 13461 3009 13495 3043
rect 14197 3009 14231 3043
rect 14565 3009 14599 3043
rect 14933 3009 14967 3043
rect 15669 3009 15703 3043
rect 15853 3009 15887 3043
rect 17049 3009 17083 3043
rect 17141 3009 17175 3043
rect 17233 3009 17267 3043
rect 17351 3009 17385 3043
rect 17509 3009 17543 3043
rect 18429 3009 18463 3043
rect 18797 3009 18831 3043
rect 19257 3009 19291 3043
rect 19349 3009 19383 3043
rect 19809 3009 19843 3043
rect 20453 3009 20487 3043
rect 2605 2941 2639 2975
rect 5181 2941 5215 2975
rect 7481 2941 7515 2975
rect 8125 2941 8159 2975
rect 11713 2941 11747 2975
rect 12173 2941 12207 2975
rect 2973 2873 3007 2907
rect 4169 2873 4203 2907
rect 7665 2873 7699 2907
rect 9229 2873 9263 2907
rect 13001 2873 13035 2907
rect 18061 2873 18095 2907
rect 21281 2873 21315 2907
rect 1777 2805 1811 2839
rect 8217 2805 8251 2839
rect 8309 2805 8343 2839
rect 9137 2805 9171 2839
rect 10609 2805 10643 2839
rect 22017 2805 22051 2839
rect 22661 2805 22695 2839
rect 4905 2601 4939 2635
rect 8401 2601 8435 2635
rect 9137 2601 9171 2635
rect 12081 2601 12115 2635
rect 15853 2601 15887 2635
rect 16957 2601 16991 2635
rect 4537 2533 4571 2567
rect 4629 2533 4663 2567
rect 15485 2533 15519 2567
rect 7757 2465 7791 2499
rect 8125 2465 8159 2499
rect 8217 2465 8251 2499
rect 11161 2465 11195 2499
rect 15393 2465 15427 2499
rect 17877 2465 17911 2499
rect 2513 2397 2547 2431
rect 3433 2397 3467 2431
rect 4445 2397 4479 2431
rect 4721 2397 4755 2431
rect 5917 2397 5951 2431
rect 7021 2397 7055 2431
rect 9873 2397 9907 2431
rect 10517 2397 10551 2431
rect 11713 2397 11747 2431
rect 11897 2397 11931 2431
rect 12541 2397 12575 2431
rect 13185 2397 13219 2431
rect 14289 2397 14323 2431
rect 15669 2397 15703 2431
rect 17141 2397 17175 2431
rect 17417 2397 17451 2431
rect 18521 2397 18555 2431
rect 19441 2397 19475 2431
rect 20085 2397 20119 2431
rect 20729 2397 20763 2431
rect 22017 2397 22051 2431
rect 22661 2397 22695 2431
rect 2237 2329 2271 2363
rect 3157 2329 3191 2363
rect 5641 2329 5675 2363
rect 6745 2329 6779 2363
rect 17325 2329 17359 2363
<< metal1 >>
rect 1104 22330 23828 22352
rect 1104 22278 3790 22330
rect 3842 22278 3854 22330
rect 3906 22278 3918 22330
rect 3970 22278 3982 22330
rect 4034 22278 4046 22330
rect 4098 22278 9471 22330
rect 9523 22278 9535 22330
rect 9587 22278 9599 22330
rect 9651 22278 9663 22330
rect 9715 22278 9727 22330
rect 9779 22278 15152 22330
rect 15204 22278 15216 22330
rect 15268 22278 15280 22330
rect 15332 22278 15344 22330
rect 15396 22278 15408 22330
rect 15460 22278 20833 22330
rect 20885 22278 20897 22330
rect 20949 22278 20961 22330
rect 21013 22278 21025 22330
rect 21077 22278 21089 22330
rect 21141 22278 23828 22330
rect 1104 22256 23828 22278
rect 11977 22151 12035 22157
rect 11977 22117 11989 22151
rect 12023 22148 12035 22151
rect 12710 22148 12716 22160
rect 12023 22120 12716 22148
rect 12023 22117 12035 22120
rect 11977 22111 12035 22117
rect 12710 22108 12716 22120
rect 12768 22108 12774 22160
rect 12066 22040 12072 22092
rect 12124 22080 12130 22092
rect 12345 22083 12403 22089
rect 12345 22080 12357 22083
rect 12124 22052 12357 22080
rect 12124 22040 12130 22052
rect 12345 22049 12357 22052
rect 12391 22049 12403 22083
rect 12345 22043 12403 22049
rect 12437 22083 12495 22089
rect 12437 22049 12449 22083
rect 12483 22080 12495 22083
rect 15654 22080 15660 22092
rect 12483 22052 15660 22080
rect 12483 22049 12495 22052
rect 12437 22043 12495 22049
rect 15654 22040 15660 22052
rect 15712 22040 15718 22092
rect 2038 21972 2044 22024
rect 2096 21972 2102 22024
rect 4522 21972 4528 22024
rect 4580 21972 4586 22024
rect 4792 22015 4850 22021
rect 4792 21981 4804 22015
rect 4838 22012 4850 22015
rect 11974 22012 11980 22024
rect 4838 21984 11980 22012
rect 4838 21981 4850 21984
rect 4792 21975 4850 21981
rect 11974 21972 11980 21984
rect 12032 21972 12038 22024
rect 12161 22015 12219 22021
rect 12161 21981 12173 22015
rect 12207 21981 12219 22015
rect 12161 21975 12219 21981
rect 2308 21947 2366 21953
rect 2308 21913 2320 21947
rect 2354 21944 2366 21947
rect 2590 21944 2596 21956
rect 2354 21916 2596 21944
rect 2354 21913 2366 21916
rect 2308 21907 2366 21913
rect 2590 21904 2596 21916
rect 2648 21904 2654 21956
rect 7101 21947 7159 21953
rect 7101 21913 7113 21947
rect 7147 21944 7159 21947
rect 7466 21944 7472 21956
rect 7147 21916 7472 21944
rect 7147 21913 7159 21916
rect 7101 21907 7159 21913
rect 7466 21904 7472 21916
rect 7524 21944 7530 21956
rect 7653 21947 7711 21953
rect 7653 21944 7665 21947
rect 7524 21916 7665 21944
rect 7524 21904 7530 21916
rect 7653 21913 7665 21916
rect 7699 21913 7711 21947
rect 12176 21944 12204 21975
rect 12526 21972 12532 22024
rect 12584 22012 12590 22024
rect 12989 22015 13047 22021
rect 12989 22012 13001 22015
rect 12584 21984 13001 22012
rect 12584 21972 12590 21984
rect 12989 21981 13001 21984
rect 13035 22012 13047 22015
rect 13633 22015 13691 22021
rect 13633 22012 13645 22015
rect 13035 21984 13645 22012
rect 13035 21981 13047 21984
rect 12989 21975 13047 21981
rect 13633 21981 13645 21984
rect 13679 21981 13691 22015
rect 13633 21975 13691 21981
rect 20438 21972 20444 22024
rect 20496 21972 20502 22024
rect 20625 22015 20683 22021
rect 20625 21981 20637 22015
rect 20671 22012 20683 22015
rect 20714 22012 20720 22024
rect 20671 21984 20720 22012
rect 20671 21981 20683 21984
rect 20625 21975 20683 21981
rect 20714 21972 20720 21984
rect 20772 22012 20778 22024
rect 22465 22015 22523 22021
rect 22465 22012 22477 22015
rect 20772 21984 22477 22012
rect 20772 21972 20778 21984
rect 22465 21981 22477 21984
rect 22511 21981 22523 22015
rect 22465 21975 22523 21981
rect 12176 21916 12434 21944
rect 7653 21907 7711 21913
rect 3234 21836 3240 21888
rect 3292 21876 3298 21888
rect 3421 21879 3479 21885
rect 3421 21876 3433 21879
rect 3292 21848 3433 21876
rect 3292 21836 3298 21848
rect 3421 21845 3433 21848
rect 3467 21845 3479 21879
rect 3421 21839 3479 21845
rect 5905 21879 5963 21885
rect 5905 21845 5917 21879
rect 5951 21876 5963 21879
rect 6086 21876 6092 21888
rect 5951 21848 6092 21876
rect 5951 21845 5963 21848
rect 5905 21839 5963 21845
rect 6086 21836 6092 21848
rect 6144 21836 6150 21888
rect 7374 21836 7380 21888
rect 7432 21876 7438 21888
rect 7745 21879 7803 21885
rect 7745 21876 7757 21879
rect 7432 21848 7757 21876
rect 7432 21836 7438 21848
rect 7745 21845 7757 21848
rect 7791 21845 7803 21879
rect 12406 21876 12434 21916
rect 13170 21904 13176 21956
rect 13228 21904 13234 21956
rect 17037 21947 17095 21953
rect 17037 21913 17049 21947
rect 17083 21944 17095 21947
rect 17402 21944 17408 21956
rect 17083 21916 17408 21944
rect 17083 21913 17095 21916
rect 17037 21907 17095 21913
rect 17402 21904 17408 21916
rect 17460 21944 17466 21956
rect 17589 21947 17647 21953
rect 17589 21944 17601 21947
rect 17460 21916 17601 21944
rect 17460 21904 17466 21916
rect 17589 21913 17601 21916
rect 17635 21913 17647 21947
rect 17589 21907 17647 21913
rect 22646 21904 22652 21956
rect 22704 21904 22710 21956
rect 13078 21876 13084 21888
rect 12406 21848 13084 21876
rect 7745 21839 7803 21845
rect 13078 21836 13084 21848
rect 13136 21876 13142 21888
rect 14277 21879 14335 21885
rect 14277 21876 14289 21879
rect 13136 21848 14289 21876
rect 13136 21836 13142 21848
rect 14277 21845 14289 21848
rect 14323 21845 14335 21879
rect 14277 21839 14335 21845
rect 14734 21836 14740 21888
rect 14792 21876 14798 21888
rect 15013 21879 15071 21885
rect 15013 21876 15025 21879
rect 14792 21848 15025 21876
rect 14792 21836 14798 21848
rect 15013 21845 15025 21848
rect 15059 21845 15071 21879
rect 15013 21839 15071 21845
rect 15657 21879 15715 21885
rect 15657 21845 15669 21879
rect 15703 21876 15715 21879
rect 15838 21876 15844 21888
rect 15703 21848 15844 21876
rect 15703 21845 15715 21848
rect 15657 21839 15715 21845
rect 15838 21836 15844 21848
rect 15896 21836 15902 21888
rect 17681 21879 17739 21885
rect 17681 21845 17693 21879
rect 17727 21876 17739 21879
rect 18874 21876 18880 21888
rect 17727 21848 18880 21876
rect 17727 21845 17739 21848
rect 17681 21839 17739 21845
rect 18874 21836 18880 21848
rect 18932 21836 18938 21888
rect 19242 21836 19248 21888
rect 19300 21876 19306 21888
rect 20533 21879 20591 21885
rect 20533 21876 20545 21879
rect 19300 21848 20545 21876
rect 19300 21836 19306 21848
rect 20533 21845 20545 21848
rect 20579 21876 20591 21879
rect 22830 21876 22836 21888
rect 20579 21848 22836 21876
rect 20579 21845 20591 21848
rect 20533 21839 20591 21845
rect 22830 21836 22836 21848
rect 22888 21836 22894 21888
rect 1104 21786 23987 21808
rect 1104 21734 6630 21786
rect 6682 21734 6694 21786
rect 6746 21734 6758 21786
rect 6810 21734 6822 21786
rect 6874 21734 6886 21786
rect 6938 21734 12311 21786
rect 12363 21734 12375 21786
rect 12427 21734 12439 21786
rect 12491 21734 12503 21786
rect 12555 21734 12567 21786
rect 12619 21734 17992 21786
rect 18044 21734 18056 21786
rect 18108 21734 18120 21786
rect 18172 21734 18184 21786
rect 18236 21734 18248 21786
rect 18300 21734 23673 21786
rect 23725 21734 23737 21786
rect 23789 21734 23801 21786
rect 23853 21734 23865 21786
rect 23917 21734 23929 21786
rect 23981 21734 23987 21786
rect 1104 21712 23987 21734
rect 18601 21675 18659 21681
rect 18601 21672 18613 21675
rect 8588 21644 18613 21672
rect 3694 21564 3700 21616
rect 3752 21604 3758 21616
rect 3890 21607 3948 21613
rect 3890 21604 3902 21607
rect 3752 21576 3902 21604
rect 3752 21564 3758 21576
rect 3890 21573 3902 21576
rect 3936 21573 3948 21607
rect 4522 21604 4528 21616
rect 3890 21567 3948 21573
rect 4172 21576 4528 21604
rect 4172 21548 4200 21576
rect 4522 21564 4528 21576
rect 4580 21604 4586 21616
rect 6816 21607 6874 21613
rect 4580 21576 6040 21604
rect 4580 21564 4586 21576
rect 4154 21496 4160 21548
rect 4212 21496 4218 21548
rect 5718 21496 5724 21548
rect 5776 21545 5782 21548
rect 6012 21545 6040 21576
rect 6816 21573 6828 21607
rect 6862 21604 6874 21607
rect 8588 21604 8616 21644
rect 18601 21641 18613 21644
rect 18647 21641 18659 21675
rect 18601 21635 18659 21641
rect 19242 21632 19248 21684
rect 19300 21632 19306 21684
rect 21085 21675 21143 21681
rect 21085 21672 21097 21675
rect 19996 21644 21097 21672
rect 6862 21576 8616 21604
rect 8656 21607 8714 21613
rect 6862 21573 6874 21576
rect 6816 21567 6874 21573
rect 8656 21573 8668 21607
rect 8702 21604 8714 21607
rect 15010 21604 15016 21616
rect 8702 21576 15016 21604
rect 8702 21573 8714 21576
rect 8656 21567 8714 21573
rect 15010 21564 15016 21576
rect 15068 21564 15074 21616
rect 15930 21564 15936 21616
rect 15988 21564 15994 21616
rect 19426 21604 19432 21616
rect 17972 21576 19432 21604
rect 5776 21499 5788 21545
rect 5997 21539 6055 21545
rect 5997 21505 6009 21539
rect 6043 21505 6055 21539
rect 5997 21499 6055 21505
rect 5776 21496 5782 21499
rect 6086 21496 6092 21548
rect 6144 21536 6150 21548
rect 9950 21536 9956 21548
rect 6144 21508 9956 21536
rect 6144 21496 6150 21508
rect 9950 21496 9956 21508
rect 10008 21496 10014 21548
rect 12158 21496 12164 21548
rect 12216 21536 12222 21548
rect 12345 21539 12403 21545
rect 12345 21536 12357 21539
rect 12216 21508 12357 21536
rect 12216 21496 12222 21508
rect 12345 21505 12357 21508
rect 12391 21505 12403 21539
rect 12345 21499 12403 21505
rect 12434 21496 12440 21548
rect 12492 21496 12498 21548
rect 12526 21496 12532 21548
rect 12584 21496 12590 21548
rect 12710 21496 12716 21548
rect 12768 21496 12774 21548
rect 13078 21496 13084 21548
rect 13136 21536 13142 21548
rect 13173 21539 13231 21545
rect 13173 21536 13185 21539
rect 13136 21508 13185 21536
rect 13136 21496 13142 21508
rect 13173 21505 13185 21508
rect 13219 21505 13231 21539
rect 13173 21499 13231 21505
rect 14182 21496 14188 21548
rect 14240 21496 14246 21548
rect 14642 21496 14648 21548
rect 14700 21496 14706 21548
rect 14829 21539 14887 21545
rect 14829 21505 14841 21539
rect 14875 21536 14887 21539
rect 15838 21536 15844 21548
rect 14875 21508 15844 21536
rect 14875 21505 14887 21508
rect 14829 21499 14887 21505
rect 15838 21496 15844 21508
rect 15896 21496 15902 21548
rect 17402 21496 17408 21548
rect 17460 21536 17466 21548
rect 17773 21539 17831 21545
rect 17773 21536 17785 21539
rect 17460 21508 17785 21536
rect 17460 21496 17466 21508
rect 17773 21505 17785 21508
rect 17819 21505 17831 21539
rect 17773 21499 17831 21505
rect 17862 21496 17868 21548
rect 17920 21496 17926 21548
rect 17972 21545 18000 21576
rect 19426 21564 19432 21576
rect 19484 21564 19490 21616
rect 17957 21539 18015 21545
rect 17957 21505 17969 21539
rect 18003 21505 18015 21539
rect 17957 21499 18015 21505
rect 18138 21496 18144 21548
rect 18196 21536 18202 21548
rect 19702 21536 19708 21548
rect 18196 21508 19708 21536
rect 18196 21496 18202 21508
rect 19702 21496 19708 21508
rect 19760 21496 19766 21548
rect 6549 21471 6607 21477
rect 6549 21437 6561 21471
rect 6595 21437 6607 21471
rect 6549 21431 6607 21437
rect 2777 21335 2835 21341
rect 2777 21301 2789 21335
rect 2823 21332 2835 21335
rect 4430 21332 4436 21344
rect 2823 21304 4436 21332
rect 2823 21301 2835 21304
rect 2777 21295 2835 21301
rect 4430 21292 4436 21304
rect 4488 21292 4494 21344
rect 4614 21292 4620 21344
rect 4672 21292 4678 21344
rect 6564 21332 6592 21431
rect 8202 21428 8208 21480
rect 8260 21468 8266 21480
rect 8389 21471 8447 21477
rect 8389 21468 8401 21471
rect 8260 21440 8401 21468
rect 8260 21428 8266 21440
rect 8389 21437 8401 21440
rect 8435 21437 8447 21471
rect 8389 21431 8447 21437
rect 13814 21428 13820 21480
rect 13872 21468 13878 21480
rect 13909 21471 13967 21477
rect 13909 21468 13921 21471
rect 13872 21440 13921 21468
rect 13872 21428 13878 21440
rect 13909 21437 13921 21440
rect 13955 21437 13967 21471
rect 13909 21431 13967 21437
rect 14090 21428 14096 21480
rect 14148 21468 14154 21480
rect 17497 21471 17555 21477
rect 17497 21468 17509 21471
rect 14148 21440 17509 21468
rect 14148 21428 14154 21440
rect 17497 21437 17509 21440
rect 17543 21437 17555 21471
rect 17497 21431 17555 21437
rect 18785 21471 18843 21477
rect 18785 21437 18797 21471
rect 18831 21437 18843 21471
rect 18785 21431 18843 21437
rect 11974 21360 11980 21412
rect 12032 21400 12038 21412
rect 12161 21403 12219 21409
rect 12161 21400 12173 21403
rect 12032 21372 12173 21400
rect 12032 21360 12038 21372
rect 12161 21369 12173 21372
rect 12207 21369 12219 21403
rect 12161 21363 12219 21369
rect 14642 21360 14648 21412
rect 14700 21400 14706 21412
rect 14826 21400 14832 21412
rect 14700 21372 14832 21400
rect 14700 21360 14706 21372
rect 14826 21360 14832 21372
rect 14884 21400 14890 21412
rect 16301 21403 16359 21409
rect 14884 21372 16160 21400
rect 14884 21360 14890 21372
rect 7190 21332 7196 21344
rect 6564 21304 7196 21332
rect 7190 21292 7196 21304
rect 7248 21292 7254 21344
rect 7929 21335 7987 21341
rect 7929 21301 7941 21335
rect 7975 21332 7987 21335
rect 8110 21332 8116 21344
rect 7975 21304 8116 21332
rect 7975 21301 7987 21304
rect 7929 21295 7987 21301
rect 8110 21292 8116 21304
rect 8168 21292 8174 21344
rect 9769 21335 9827 21341
rect 9769 21301 9781 21335
rect 9815 21332 9827 21335
rect 9858 21332 9864 21344
rect 9815 21304 9864 21332
rect 9815 21301 9827 21304
rect 9769 21295 9827 21301
rect 9858 21292 9864 21304
rect 9916 21292 9922 21344
rect 13262 21292 13268 21344
rect 13320 21332 13326 21344
rect 14737 21335 14795 21341
rect 14737 21332 14749 21335
rect 13320 21304 14749 21332
rect 13320 21292 13326 21304
rect 14737 21301 14749 21304
rect 14783 21301 14795 21335
rect 14737 21295 14795 21301
rect 15746 21292 15752 21344
rect 15804 21292 15810 21344
rect 15933 21335 15991 21341
rect 15933 21301 15945 21335
rect 15979 21332 15991 21335
rect 16022 21332 16028 21344
rect 15979 21304 16028 21332
rect 15979 21301 15991 21304
rect 15933 21295 15991 21301
rect 16022 21292 16028 21304
rect 16080 21292 16086 21344
rect 16132 21332 16160 21372
rect 16301 21369 16313 21403
rect 16347 21400 16359 21403
rect 17126 21400 17132 21412
rect 16347 21372 17132 21400
rect 16347 21369 16359 21372
rect 16301 21363 16359 21369
rect 17126 21360 17132 21372
rect 17184 21360 17190 21412
rect 18800 21400 18828 21431
rect 18874 21428 18880 21480
rect 18932 21428 18938 21480
rect 19996 21400 20024 21644
rect 21085 21641 21097 21644
rect 21131 21672 21143 21675
rect 22278 21672 22284 21684
rect 21131 21644 22284 21672
rect 21131 21641 21143 21644
rect 21085 21635 21143 21641
rect 22278 21632 22284 21644
rect 22336 21632 22342 21684
rect 22370 21632 22376 21684
rect 22428 21672 22434 21684
rect 22646 21672 22652 21684
rect 22428 21644 22652 21672
rect 22428 21632 22434 21644
rect 22646 21632 22652 21644
rect 22704 21632 22710 21684
rect 20714 21564 20720 21616
rect 20772 21564 20778 21616
rect 20254 21496 20260 21548
rect 20312 21496 20318 21548
rect 20438 21496 20444 21548
rect 20496 21536 20502 21548
rect 20901 21539 20959 21545
rect 20901 21536 20913 21539
rect 20496 21508 20913 21536
rect 20496 21496 20502 21508
rect 20901 21505 20913 21508
rect 20947 21505 20959 21539
rect 20901 21499 20959 21505
rect 20073 21471 20131 21477
rect 20073 21437 20085 21471
rect 20119 21468 20131 21471
rect 20714 21468 20720 21480
rect 20119 21440 20720 21468
rect 20119 21437 20131 21440
rect 20073 21431 20131 21437
rect 18800 21372 20024 21400
rect 16945 21335 17003 21341
rect 16945 21332 16957 21335
rect 16132 21304 16957 21332
rect 16945 21301 16957 21304
rect 16991 21332 17003 21335
rect 20088 21332 20116 21431
rect 20714 21428 20720 21440
rect 20772 21428 20778 21480
rect 16991 21304 20116 21332
rect 16991 21301 17003 21304
rect 16945 21295 17003 21301
rect 1104 21242 23828 21264
rect 1104 21190 3790 21242
rect 3842 21190 3854 21242
rect 3906 21190 3918 21242
rect 3970 21190 3982 21242
rect 4034 21190 4046 21242
rect 4098 21190 9471 21242
rect 9523 21190 9535 21242
rect 9587 21190 9599 21242
rect 9651 21190 9663 21242
rect 9715 21190 9727 21242
rect 9779 21190 15152 21242
rect 15204 21190 15216 21242
rect 15268 21190 15280 21242
rect 15332 21190 15344 21242
rect 15396 21190 15408 21242
rect 15460 21190 20833 21242
rect 20885 21190 20897 21242
rect 20949 21190 20961 21242
rect 21013 21190 21025 21242
rect 21077 21190 21089 21242
rect 21141 21190 23828 21242
rect 1104 21168 23828 21190
rect 12069 21131 12127 21137
rect 12069 21097 12081 21131
rect 12115 21128 12127 21131
rect 14182 21128 14188 21140
rect 12115 21100 14188 21128
rect 12115 21097 12127 21100
rect 12069 21091 12127 21097
rect 14182 21088 14188 21100
rect 14240 21088 14246 21140
rect 14737 21131 14795 21137
rect 14737 21097 14749 21131
rect 14783 21097 14795 21131
rect 14737 21091 14795 21097
rect 8386 21020 8392 21072
rect 8444 21060 8450 21072
rect 9125 21063 9183 21069
rect 9125 21060 9137 21063
rect 8444 21032 9137 21060
rect 8444 21020 8450 21032
rect 9125 21029 9137 21032
rect 9171 21029 9183 21063
rect 9125 21023 9183 21029
rect 13173 21063 13231 21069
rect 13173 21029 13185 21063
rect 13219 21029 13231 21063
rect 13173 21023 13231 21029
rect 11425 20995 11483 21001
rect 11425 20961 11437 20995
rect 11471 20992 11483 20995
rect 12434 20992 12440 21004
rect 11471 20964 12440 20992
rect 11471 20961 11483 20964
rect 11425 20955 11483 20961
rect 12434 20952 12440 20964
rect 12492 20992 12498 21004
rect 13188 20992 13216 21023
rect 14274 21020 14280 21072
rect 14332 21060 14338 21072
rect 14752 21060 14780 21091
rect 15010 21088 15016 21140
rect 15068 21128 15074 21140
rect 15381 21131 15439 21137
rect 15381 21128 15393 21131
rect 15068 21100 15393 21128
rect 15068 21088 15074 21100
rect 15381 21097 15393 21100
rect 15427 21097 15439 21131
rect 15381 21091 15439 21097
rect 17126 21088 17132 21140
rect 17184 21088 17190 21140
rect 18138 21128 18144 21140
rect 17236 21100 18144 21128
rect 17236 21060 17264 21100
rect 18138 21088 18144 21100
rect 18196 21088 18202 21140
rect 19429 21131 19487 21137
rect 19429 21097 19441 21131
rect 19475 21128 19487 21131
rect 19518 21128 19524 21140
rect 19475 21100 19524 21128
rect 19475 21097 19487 21100
rect 19429 21091 19487 21097
rect 19518 21088 19524 21100
rect 19576 21088 19582 21140
rect 14332 21032 17264 21060
rect 14332 21020 14338 21032
rect 17402 21020 17408 21072
rect 17460 21020 17466 21072
rect 17862 21060 17868 21072
rect 17604 21032 17868 21060
rect 12492 20964 12664 20992
rect 13188 20964 15608 20992
rect 12492 20952 12498 20964
rect 1949 20927 2007 20933
rect 1949 20893 1961 20927
rect 1995 20924 2007 20927
rect 2038 20924 2044 20936
rect 1995 20896 2044 20924
rect 1995 20893 2007 20896
rect 1949 20887 2007 20893
rect 2038 20884 2044 20896
rect 2096 20884 2102 20936
rect 2498 20884 2504 20936
rect 2556 20924 2562 20936
rect 5810 20924 5816 20936
rect 2556 20896 5816 20924
rect 2556 20884 2562 20896
rect 5810 20884 5816 20896
rect 5868 20884 5874 20936
rect 7190 20884 7196 20936
rect 7248 20884 7254 20936
rect 9122 20884 9128 20936
rect 9180 20924 9186 20936
rect 12636 20933 12664 20964
rect 10505 20927 10563 20933
rect 10505 20924 10517 20927
rect 9180 20896 10517 20924
rect 9180 20884 9186 20896
rect 10505 20893 10517 20896
rect 10551 20893 10563 20927
rect 10505 20887 10563 20893
rect 11333 20927 11391 20933
rect 11333 20893 11345 20927
rect 11379 20893 11391 20927
rect 11333 20887 11391 20893
rect 12161 20927 12219 20933
rect 12161 20893 12173 20927
rect 12207 20924 12219 20927
rect 12621 20927 12679 20933
rect 12207 20896 12434 20924
rect 12207 20893 12219 20896
rect 12161 20887 12219 20893
rect 2216 20859 2274 20865
rect 2216 20825 2228 20859
rect 2262 20856 2274 20859
rect 2314 20856 2320 20868
rect 2262 20828 2320 20856
rect 2262 20825 2274 20828
rect 2216 20819 2274 20825
rect 2314 20816 2320 20828
rect 2372 20816 2378 20868
rect 6948 20859 7006 20865
rect 6948 20825 6960 20859
rect 6994 20856 7006 20859
rect 7098 20856 7104 20868
rect 6994 20828 7104 20856
rect 6994 20825 7006 20828
rect 6948 20819 7006 20825
rect 7098 20816 7104 20828
rect 7156 20816 7162 20868
rect 10260 20859 10318 20865
rect 8496 20828 10180 20856
rect 8496 20800 8524 20828
rect 2682 20748 2688 20800
rect 2740 20788 2746 20800
rect 3329 20791 3387 20797
rect 3329 20788 3341 20791
rect 2740 20760 3341 20788
rect 2740 20748 2746 20760
rect 3329 20757 3341 20760
rect 3375 20757 3387 20791
rect 3329 20751 3387 20757
rect 5626 20748 5632 20800
rect 5684 20788 5690 20800
rect 5813 20791 5871 20797
rect 5813 20788 5825 20791
rect 5684 20760 5825 20788
rect 5684 20748 5690 20760
rect 5813 20757 5825 20760
rect 5859 20757 5871 20791
rect 5813 20751 5871 20757
rect 8478 20748 8484 20800
rect 8536 20748 8542 20800
rect 10152 20788 10180 20828
rect 10260 20825 10272 20859
rect 10306 20856 10318 20859
rect 10962 20856 10968 20868
rect 10306 20828 10968 20856
rect 10306 20825 10318 20828
rect 10260 20819 10318 20825
rect 10962 20816 10968 20828
rect 11020 20816 11026 20868
rect 11054 20788 11060 20800
rect 10152 20760 11060 20788
rect 11054 20748 11060 20760
rect 11112 20788 11118 20800
rect 11348 20788 11376 20887
rect 11112 20760 11376 20788
rect 12406 20788 12434 20896
rect 12621 20893 12633 20927
rect 12667 20924 12679 20927
rect 12710 20924 12716 20936
rect 12667 20896 12716 20924
rect 12667 20893 12679 20896
rect 12621 20887 12679 20893
rect 12710 20884 12716 20896
rect 12768 20884 12774 20936
rect 12894 20884 12900 20936
rect 12952 20884 12958 20936
rect 13173 20927 13231 20933
rect 13173 20893 13185 20927
rect 13219 20924 13231 20927
rect 13262 20924 13268 20936
rect 13219 20896 13268 20924
rect 13219 20893 13231 20896
rect 13173 20887 13231 20893
rect 13262 20884 13268 20896
rect 13320 20884 13326 20936
rect 14550 20884 14556 20936
rect 14608 20884 14614 20936
rect 14734 20884 14740 20936
rect 14792 20884 14798 20936
rect 15580 20933 15608 20964
rect 16298 20952 16304 21004
rect 16356 20992 16362 21004
rect 17420 20992 17448 21020
rect 16356 20964 17448 20992
rect 16356 20952 16362 20964
rect 15473 20927 15531 20933
rect 15473 20893 15485 20927
rect 15519 20893 15531 20927
rect 15473 20887 15531 20893
rect 15565 20927 15623 20933
rect 15565 20893 15577 20927
rect 15611 20893 15623 20927
rect 15565 20887 15623 20893
rect 13449 20859 13507 20865
rect 13449 20825 13461 20859
rect 13495 20856 13507 20859
rect 14366 20856 14372 20868
rect 13495 20828 14372 20856
rect 13495 20825 13507 20828
rect 13449 20819 13507 20825
rect 14366 20816 14372 20828
rect 14424 20816 14430 20868
rect 14752 20856 14780 20884
rect 15488 20856 15516 20887
rect 15654 20884 15660 20936
rect 15712 20924 15718 20936
rect 15841 20927 15899 20933
rect 15841 20924 15853 20927
rect 15712 20896 15853 20924
rect 15712 20884 15718 20896
rect 15841 20893 15853 20896
rect 15887 20893 15899 20927
rect 15841 20887 15899 20893
rect 16206 20884 16212 20936
rect 16264 20884 16270 20936
rect 17313 20927 17371 20933
rect 17313 20893 17325 20927
rect 17359 20924 17371 20927
rect 17402 20924 17408 20936
rect 17359 20896 17408 20924
rect 17359 20893 17371 20896
rect 17313 20887 17371 20893
rect 17402 20884 17408 20896
rect 17460 20884 17466 20936
rect 17494 20884 17500 20936
rect 17552 20884 17558 20936
rect 17604 20933 17632 21032
rect 17862 21020 17868 21032
rect 17920 21060 17926 21072
rect 19334 21060 19340 21072
rect 17920 21032 19340 21060
rect 17920 21020 17926 21032
rect 19334 21020 19340 21032
rect 19392 21020 19398 21072
rect 18874 20952 18880 21004
rect 18932 20992 18938 21004
rect 18932 20964 22600 20992
rect 18932 20952 18938 20964
rect 17589 20927 17647 20933
rect 17589 20893 17601 20927
rect 17635 20893 17647 20927
rect 17589 20887 17647 20893
rect 17773 20927 17831 20933
rect 17773 20893 17785 20927
rect 17819 20924 17831 20927
rect 18138 20924 18144 20936
rect 17819 20896 18144 20924
rect 17819 20893 17831 20896
rect 17773 20887 17831 20893
rect 18138 20884 18144 20896
rect 18196 20884 18202 20936
rect 18417 20927 18475 20933
rect 18417 20893 18429 20927
rect 18463 20893 18475 20927
rect 18417 20887 18475 20893
rect 18601 20927 18659 20933
rect 18601 20893 18613 20927
rect 18647 20924 18659 20927
rect 19518 20924 19524 20936
rect 18647 20896 19524 20924
rect 18647 20893 18659 20896
rect 18601 20887 18659 20893
rect 18322 20856 18328 20868
rect 14752 20828 15424 20856
rect 15488 20828 18328 20856
rect 14274 20788 14280 20800
rect 12406 20760 14280 20788
rect 11112 20748 11118 20760
rect 14274 20748 14280 20760
rect 14332 20748 14338 20800
rect 14918 20748 14924 20800
rect 14976 20748 14982 20800
rect 15396 20788 15424 20828
rect 18322 20816 18328 20828
rect 18380 20816 18386 20868
rect 18230 20788 18236 20800
rect 15396 20760 18236 20788
rect 18230 20748 18236 20760
rect 18288 20748 18294 20800
rect 18432 20788 18460 20887
rect 19518 20884 19524 20896
rect 19576 20884 19582 20936
rect 19610 20884 19616 20936
rect 19668 20884 19674 20936
rect 19705 20927 19763 20933
rect 19705 20893 19717 20927
rect 19751 20924 19763 20927
rect 19794 20924 19800 20936
rect 19751 20896 19800 20924
rect 19751 20893 19763 20896
rect 19705 20887 19763 20893
rect 19794 20884 19800 20896
rect 19852 20884 19858 20936
rect 19889 20927 19947 20933
rect 19889 20893 19901 20927
rect 19935 20893 19947 20927
rect 19889 20887 19947 20893
rect 19981 20927 20039 20933
rect 19981 20893 19993 20927
rect 20027 20924 20039 20927
rect 20162 20924 20168 20936
rect 20027 20896 20168 20924
rect 20027 20893 20039 20896
rect 19981 20887 20039 20893
rect 18509 20859 18567 20865
rect 18509 20825 18521 20859
rect 18555 20856 18567 20859
rect 19904 20856 19932 20887
rect 20162 20884 20168 20896
rect 20220 20884 20226 20936
rect 20441 20927 20499 20933
rect 20441 20893 20453 20927
rect 20487 20924 20499 20927
rect 20622 20924 20628 20936
rect 20487 20896 20628 20924
rect 20487 20893 20499 20896
rect 20441 20887 20499 20893
rect 20622 20884 20628 20896
rect 20680 20884 20686 20936
rect 22572 20933 22600 20964
rect 22646 20952 22652 21004
rect 22704 20952 22710 21004
rect 22557 20927 22615 20933
rect 22557 20893 22569 20927
rect 22603 20893 22615 20927
rect 22557 20887 22615 20893
rect 18555 20828 19932 20856
rect 18555 20825 18567 20828
rect 18509 20819 18567 20825
rect 20070 20816 20076 20868
rect 20128 20856 20134 20868
rect 20717 20859 20775 20865
rect 20717 20856 20729 20859
rect 20128 20828 20729 20856
rect 20128 20816 20134 20828
rect 20717 20825 20729 20828
rect 20763 20825 20775 20859
rect 20717 20819 20775 20825
rect 21910 20816 21916 20868
rect 21968 20816 21974 20868
rect 20254 20788 20260 20800
rect 18432 20760 20260 20788
rect 20254 20748 20260 20760
rect 20312 20748 20318 20800
rect 1104 20698 23987 20720
rect 1104 20646 6630 20698
rect 6682 20646 6694 20698
rect 6746 20646 6758 20698
rect 6810 20646 6822 20698
rect 6874 20646 6886 20698
rect 6938 20646 12311 20698
rect 12363 20646 12375 20698
rect 12427 20646 12439 20698
rect 12491 20646 12503 20698
rect 12555 20646 12567 20698
rect 12619 20646 17992 20698
rect 18044 20646 18056 20698
rect 18108 20646 18120 20698
rect 18172 20646 18184 20698
rect 18236 20646 18248 20698
rect 18300 20646 23673 20698
rect 23725 20646 23737 20698
rect 23789 20646 23801 20698
rect 23853 20646 23865 20698
rect 23917 20646 23929 20698
rect 23981 20646 23987 20698
rect 1104 20624 23987 20646
rect 2038 20544 2044 20596
rect 2096 20584 2102 20596
rect 3053 20587 3111 20593
rect 3053 20584 3065 20587
rect 2096 20556 3065 20584
rect 2096 20544 2102 20556
rect 3053 20553 3065 20556
rect 3099 20584 3111 20587
rect 4154 20584 4160 20596
rect 3099 20556 4160 20584
rect 3099 20553 3111 20556
rect 3053 20547 3111 20553
rect 4154 20544 4160 20556
rect 4212 20544 4218 20596
rect 11054 20544 11060 20596
rect 11112 20584 11118 20596
rect 13630 20584 13636 20596
rect 11112 20556 12434 20584
rect 11112 20544 11118 20556
rect 12406 20516 12434 20556
rect 13096 20556 13636 20584
rect 13096 20528 13124 20556
rect 13630 20544 13636 20556
rect 13688 20584 13694 20596
rect 13688 20556 15332 20584
rect 13688 20544 13694 20556
rect 13078 20516 13084 20528
rect 12406 20488 13084 20516
rect 13078 20476 13084 20488
rect 13136 20476 13142 20528
rect 13541 20519 13599 20525
rect 13541 20485 13553 20519
rect 13587 20516 13599 20519
rect 14090 20516 14096 20528
rect 13587 20488 14096 20516
rect 13587 20485 13599 20488
rect 13541 20479 13599 20485
rect 14090 20476 14096 20488
rect 14148 20476 14154 20528
rect 15194 20516 15200 20528
rect 14476 20488 15200 20516
rect 4338 20408 4344 20460
rect 4396 20408 4402 20460
rect 8472 20451 8530 20457
rect 8472 20417 8484 20451
rect 8518 20448 8530 20451
rect 10045 20451 10103 20457
rect 10045 20448 10057 20451
rect 8518 20420 10057 20448
rect 8518 20417 8530 20420
rect 8472 20411 8530 20417
rect 10045 20417 10057 20420
rect 10091 20448 10103 20451
rect 11422 20448 11428 20460
rect 10091 20420 11428 20448
rect 10091 20417 10103 20420
rect 10045 20411 10103 20417
rect 11422 20408 11428 20420
rect 11480 20408 11486 20460
rect 12529 20451 12587 20457
rect 12529 20417 12541 20451
rect 12575 20448 12587 20451
rect 12575 20420 13676 20448
rect 12575 20417 12587 20420
rect 12529 20411 12587 20417
rect 8202 20340 8208 20392
rect 8260 20340 8266 20392
rect 12621 20383 12679 20389
rect 12621 20349 12633 20383
rect 12667 20349 12679 20383
rect 12621 20343 12679 20349
rect 12805 20383 12863 20389
rect 12805 20349 12817 20383
rect 12851 20380 12863 20383
rect 13078 20380 13084 20392
rect 12851 20352 13084 20380
rect 12851 20349 12863 20352
rect 12805 20343 12863 20349
rect 8220 20244 8248 20340
rect 9585 20315 9643 20321
rect 9585 20281 9597 20315
rect 9631 20312 9643 20315
rect 11238 20312 11244 20324
rect 9631 20284 11244 20312
rect 9631 20281 9643 20284
rect 9585 20275 9643 20281
rect 11238 20272 11244 20284
rect 11296 20272 11302 20324
rect 12636 20312 12664 20343
rect 13078 20340 13084 20352
rect 13136 20340 13142 20392
rect 13541 20315 13599 20321
rect 13541 20312 13553 20315
rect 12636 20284 13553 20312
rect 13541 20281 13553 20284
rect 13587 20281 13599 20315
rect 13648 20312 13676 20420
rect 13722 20408 13728 20460
rect 13780 20408 13786 20460
rect 13814 20408 13820 20460
rect 13872 20408 13878 20460
rect 14274 20408 14280 20460
rect 14332 20408 14338 20460
rect 14476 20457 14504 20488
rect 15194 20476 15200 20488
rect 15252 20476 15258 20528
rect 14461 20451 14519 20457
rect 14461 20417 14473 20451
rect 14507 20417 14519 20451
rect 14461 20411 14519 20417
rect 14918 20408 14924 20460
rect 14976 20448 14982 20460
rect 15304 20457 15332 20556
rect 18322 20544 18328 20596
rect 18380 20584 18386 20596
rect 20073 20587 20131 20593
rect 20073 20584 20085 20587
rect 18380 20556 20085 20584
rect 18380 20544 18386 20556
rect 20073 20553 20085 20556
rect 20119 20553 20131 20587
rect 20073 20547 20131 20553
rect 20714 20544 20720 20596
rect 20772 20544 20778 20596
rect 22646 20544 22652 20596
rect 22704 20544 22710 20596
rect 15654 20476 15660 20528
rect 15712 20516 15718 20528
rect 16390 20516 16396 20528
rect 15712 20488 16396 20516
rect 15712 20476 15718 20488
rect 16390 20476 16396 20488
rect 16448 20516 16454 20528
rect 16448 20488 20024 20516
rect 16448 20476 16454 20488
rect 15105 20451 15163 20457
rect 15105 20448 15117 20451
rect 14976 20420 15117 20448
rect 14976 20408 14982 20420
rect 15105 20417 15117 20420
rect 15151 20417 15163 20451
rect 15105 20411 15163 20417
rect 15289 20451 15347 20457
rect 15289 20417 15301 20451
rect 15335 20417 15347 20451
rect 15289 20411 15347 20417
rect 15381 20451 15439 20457
rect 15381 20417 15393 20451
rect 15427 20448 15439 20451
rect 15746 20448 15752 20460
rect 15427 20420 15752 20448
rect 15427 20417 15439 20420
rect 15381 20411 15439 20417
rect 14369 20383 14427 20389
rect 14369 20349 14381 20383
rect 14415 20380 14427 20383
rect 15197 20383 15255 20389
rect 15197 20380 15209 20383
rect 14415 20352 15209 20380
rect 14415 20349 14427 20352
rect 14369 20343 14427 20349
rect 15197 20349 15209 20352
rect 15243 20349 15255 20383
rect 15304 20380 15332 20411
rect 15746 20408 15752 20420
rect 15804 20408 15810 20460
rect 19996 20457 20024 20488
rect 20254 20476 20260 20528
rect 20312 20516 20318 20528
rect 22097 20519 22155 20525
rect 22097 20516 22109 20519
rect 20312 20488 22109 20516
rect 20312 20476 20318 20488
rect 22097 20485 22109 20488
rect 22143 20485 22155 20519
rect 22097 20479 22155 20485
rect 19981 20451 20039 20457
rect 19981 20417 19993 20451
rect 20027 20417 20039 20451
rect 19981 20411 20039 20417
rect 20165 20451 20223 20457
rect 20165 20417 20177 20451
rect 20211 20417 20223 20451
rect 20165 20411 20223 20417
rect 15562 20380 15568 20392
rect 15304 20352 15568 20380
rect 15197 20343 15255 20349
rect 15562 20340 15568 20352
rect 15620 20340 15626 20392
rect 20180 20380 20208 20411
rect 22002 20408 22008 20460
rect 22060 20408 22066 20460
rect 22278 20408 22284 20460
rect 22336 20448 22342 20460
rect 22649 20451 22707 20457
rect 22649 20448 22661 20451
rect 22336 20420 22661 20448
rect 22336 20408 22342 20420
rect 22649 20417 22661 20420
rect 22695 20417 22707 20451
rect 22649 20411 22707 20417
rect 22830 20408 22836 20460
rect 22888 20408 22894 20460
rect 22554 20380 22560 20392
rect 20180 20352 22560 20380
rect 22554 20340 22560 20352
rect 22612 20340 22618 20392
rect 15746 20312 15752 20324
rect 13648 20284 15752 20312
rect 13541 20275 13599 20281
rect 15746 20272 15752 20284
rect 15804 20272 15810 20324
rect 16025 20315 16083 20321
rect 16025 20281 16037 20315
rect 16071 20312 16083 20315
rect 16114 20312 16120 20324
rect 16071 20284 16120 20312
rect 16071 20281 16083 20284
rect 16025 20275 16083 20281
rect 16114 20272 16120 20284
rect 16172 20312 16178 20324
rect 19337 20315 19395 20321
rect 19337 20312 19349 20315
rect 16172 20284 19349 20312
rect 16172 20272 16178 20284
rect 19337 20281 19349 20284
rect 19383 20312 19395 20315
rect 20162 20312 20168 20324
rect 19383 20284 20168 20312
rect 19383 20281 19395 20284
rect 19337 20275 19395 20281
rect 20162 20272 20168 20284
rect 20220 20312 20226 20324
rect 20530 20312 20536 20324
rect 20220 20284 20536 20312
rect 20220 20272 20226 20284
rect 20530 20272 20536 20284
rect 20588 20272 20594 20324
rect 9122 20244 9128 20256
rect 8220 20216 9128 20244
rect 9122 20204 9128 20216
rect 9180 20204 9186 20256
rect 11054 20204 11060 20256
rect 11112 20244 11118 20256
rect 12161 20247 12219 20253
rect 12161 20244 12173 20247
rect 11112 20216 12173 20244
rect 11112 20204 11118 20216
rect 12161 20213 12173 20216
rect 12207 20213 12219 20247
rect 12161 20207 12219 20213
rect 14918 20204 14924 20256
rect 14976 20204 14982 20256
rect 1104 20154 23828 20176
rect 1104 20102 3790 20154
rect 3842 20102 3854 20154
rect 3906 20102 3918 20154
rect 3970 20102 3982 20154
rect 4034 20102 4046 20154
rect 4098 20102 9471 20154
rect 9523 20102 9535 20154
rect 9587 20102 9599 20154
rect 9651 20102 9663 20154
rect 9715 20102 9727 20154
rect 9779 20102 15152 20154
rect 15204 20102 15216 20154
rect 15268 20102 15280 20154
rect 15332 20102 15344 20154
rect 15396 20102 15408 20154
rect 15460 20102 20833 20154
rect 20885 20102 20897 20154
rect 20949 20102 20961 20154
rect 21013 20102 21025 20154
rect 21077 20102 21089 20154
rect 21141 20102 23828 20154
rect 1104 20080 23828 20102
rect 11422 20000 11428 20052
rect 11480 20000 11486 20052
rect 11977 20043 12035 20049
rect 11977 20009 11989 20043
rect 12023 20040 12035 20043
rect 12066 20040 12072 20052
rect 12023 20012 12072 20040
rect 12023 20009 12035 20012
rect 11977 20003 12035 20009
rect 12066 20000 12072 20012
rect 12124 20000 12130 20052
rect 13265 20043 13323 20049
rect 13265 20009 13277 20043
rect 13311 20040 13323 20043
rect 14274 20040 14280 20052
rect 13311 20012 14280 20040
rect 13311 20009 13323 20012
rect 13265 20003 13323 20009
rect 14274 20000 14280 20012
rect 14332 20000 14338 20052
rect 15010 20040 15016 20052
rect 14476 20012 15016 20040
rect 3421 19907 3479 19913
rect 3421 19873 3433 19907
rect 3467 19904 3479 19907
rect 4154 19904 4160 19916
rect 3467 19876 4160 19904
rect 3467 19873 3479 19876
rect 3421 19867 3479 19873
rect 4154 19864 4160 19876
rect 4212 19864 4218 19916
rect 6733 19839 6791 19845
rect 6733 19805 6745 19839
rect 6779 19836 6791 19839
rect 7190 19836 7196 19848
rect 6779 19808 7196 19836
rect 6779 19805 6791 19808
rect 6733 19799 6791 19805
rect 7190 19796 7196 19808
rect 7248 19836 7254 19848
rect 8202 19836 8208 19848
rect 7248 19808 8208 19836
rect 7248 19796 7254 19808
rect 8202 19796 8208 19808
rect 8260 19836 8266 19848
rect 9122 19836 9128 19848
rect 8260 19808 9128 19836
rect 8260 19796 8266 19808
rect 9122 19796 9128 19808
rect 9180 19796 9186 19848
rect 9401 19839 9459 19845
rect 9401 19805 9413 19839
rect 9447 19836 9459 19839
rect 11330 19836 11336 19848
rect 9447 19808 11336 19836
rect 9447 19805 9459 19808
rect 9401 19799 9459 19805
rect 11330 19796 11336 19808
rect 11388 19796 11394 19848
rect 11440 19836 11468 20000
rect 12253 19975 12311 19981
rect 12253 19941 12265 19975
rect 12299 19972 12311 19975
rect 14476 19972 14504 20012
rect 15010 20000 15016 20012
rect 15068 20000 15074 20052
rect 15562 20000 15568 20052
rect 15620 20000 15626 20052
rect 19426 20000 19432 20052
rect 19484 20000 19490 20052
rect 12299 19944 14504 19972
rect 12299 19941 12311 19944
rect 12253 19935 12311 19941
rect 14550 19932 14556 19984
rect 14608 19972 14614 19984
rect 22278 19972 22284 19984
rect 14608 19944 22284 19972
rect 14608 19932 14614 19944
rect 22278 19932 22284 19944
rect 22336 19932 22342 19984
rect 11974 19864 11980 19916
rect 12032 19904 12038 19916
rect 12345 19907 12403 19913
rect 12345 19904 12357 19907
rect 12032 19876 12357 19904
rect 12032 19864 12038 19876
rect 12345 19873 12357 19876
rect 12391 19873 12403 19907
rect 12345 19867 12403 19873
rect 12437 19907 12495 19913
rect 12437 19873 12449 19907
rect 12483 19904 12495 19907
rect 14568 19904 14596 19932
rect 12483 19876 14596 19904
rect 12483 19873 12495 19876
rect 12437 19867 12495 19873
rect 15102 19864 15108 19916
rect 15160 19904 15166 19916
rect 15654 19904 15660 19916
rect 15160 19876 15660 19904
rect 15160 19864 15166 19876
rect 15654 19864 15660 19876
rect 15712 19904 15718 19916
rect 16114 19904 16120 19916
rect 15712 19876 16120 19904
rect 15712 19864 15718 19876
rect 16114 19864 16120 19876
rect 16172 19864 16178 19916
rect 22002 19904 22008 19916
rect 19628 19876 22008 19904
rect 12161 19839 12219 19845
rect 12161 19836 12173 19839
rect 11440 19808 12173 19836
rect 12161 19805 12173 19808
rect 12207 19805 12219 19839
rect 12161 19799 12219 19805
rect 12621 19839 12679 19845
rect 12621 19805 12633 19839
rect 12667 19805 12679 19839
rect 12621 19799 12679 19805
rect 2958 19728 2964 19780
rect 3016 19768 3022 19780
rect 3154 19771 3212 19777
rect 3154 19768 3166 19771
rect 3016 19740 3166 19768
rect 3016 19728 3022 19740
rect 3154 19737 3166 19740
rect 3200 19737 3212 19771
rect 3154 19731 3212 19737
rect 6178 19728 6184 19780
rect 6236 19768 6242 19780
rect 6466 19771 6524 19777
rect 6466 19768 6478 19771
rect 6236 19740 6478 19768
rect 6236 19728 6242 19740
rect 6466 19737 6478 19740
rect 6512 19737 6524 19771
rect 6466 19731 6524 19737
rect 7460 19771 7518 19777
rect 7460 19737 7472 19771
rect 7506 19768 7518 19771
rect 8478 19768 8484 19780
rect 7506 19740 8484 19768
rect 7506 19737 7518 19740
rect 7460 19731 7518 19737
rect 8478 19728 8484 19740
rect 8536 19728 8542 19780
rect 2041 19703 2099 19709
rect 2041 19669 2053 19703
rect 2087 19700 2099 19703
rect 2406 19700 2412 19712
rect 2087 19672 2412 19700
rect 2087 19669 2099 19672
rect 2041 19663 2099 19669
rect 2406 19660 2412 19672
rect 2464 19660 2470 19712
rect 5350 19660 5356 19712
rect 5408 19660 5414 19712
rect 8573 19703 8631 19709
rect 8573 19669 8585 19703
rect 8619 19700 8631 19703
rect 9214 19700 9220 19712
rect 8619 19672 9220 19700
rect 8619 19669 8631 19672
rect 8573 19663 8631 19669
rect 9214 19660 9220 19672
rect 9272 19660 9278 19712
rect 10318 19660 10324 19712
rect 10376 19700 10382 19712
rect 10505 19703 10563 19709
rect 10505 19700 10517 19703
rect 10376 19672 10517 19700
rect 10376 19660 10382 19672
rect 10505 19669 10517 19672
rect 10551 19669 10563 19703
rect 12176 19700 12204 19799
rect 12636 19768 12664 19799
rect 13446 19796 13452 19848
rect 13504 19796 13510 19848
rect 14366 19796 14372 19848
rect 14424 19796 14430 19848
rect 14550 19796 14556 19848
rect 14608 19796 14614 19848
rect 17402 19796 17408 19848
rect 17460 19836 17466 19848
rect 18322 19836 18328 19848
rect 17460 19808 18328 19836
rect 17460 19796 17466 19808
rect 18322 19796 18328 19808
rect 18380 19836 18386 19848
rect 19628 19845 19656 19876
rect 22002 19864 22008 19876
rect 22060 19864 22066 19916
rect 19613 19839 19671 19845
rect 19613 19836 19625 19839
rect 18380 19808 19625 19836
rect 18380 19796 18386 19808
rect 19613 19805 19625 19808
rect 19659 19805 19671 19839
rect 19613 19799 19671 19805
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19836 19947 19839
rect 20070 19836 20076 19848
rect 19935 19808 20076 19836
rect 19935 19805 19947 19808
rect 19889 19799 19947 19805
rect 20070 19796 20076 19808
rect 20128 19796 20134 19848
rect 16298 19768 16304 19780
rect 12636 19740 16304 19768
rect 16298 19728 16304 19740
rect 16356 19728 16362 19780
rect 13906 19700 13912 19712
rect 12176 19672 13912 19700
rect 10505 19663 10563 19669
rect 13906 19660 13912 19672
rect 13964 19660 13970 19712
rect 14458 19660 14464 19712
rect 14516 19660 14522 19712
rect 18782 19660 18788 19712
rect 18840 19700 18846 19712
rect 19797 19703 19855 19709
rect 19797 19700 19809 19703
rect 18840 19672 19809 19700
rect 18840 19660 18846 19672
rect 19797 19669 19809 19672
rect 19843 19669 19855 19703
rect 19797 19663 19855 19669
rect 1104 19610 23987 19632
rect 1104 19558 6630 19610
rect 6682 19558 6694 19610
rect 6746 19558 6758 19610
rect 6810 19558 6822 19610
rect 6874 19558 6886 19610
rect 6938 19558 12311 19610
rect 12363 19558 12375 19610
rect 12427 19558 12439 19610
rect 12491 19558 12503 19610
rect 12555 19558 12567 19610
rect 12619 19558 17992 19610
rect 18044 19558 18056 19610
rect 18108 19558 18120 19610
rect 18172 19558 18184 19610
rect 18236 19558 18248 19610
rect 18300 19558 23673 19610
rect 23725 19558 23737 19610
rect 23789 19558 23801 19610
rect 23853 19558 23865 19610
rect 23917 19558 23929 19610
rect 23981 19558 23987 19610
rect 1104 19536 23987 19558
rect 9585 19499 9643 19505
rect 9585 19465 9597 19499
rect 9631 19496 9643 19499
rect 10686 19496 10692 19508
rect 9631 19468 10692 19496
rect 9631 19465 9643 19468
rect 9585 19459 9643 19465
rect 10686 19456 10692 19468
rect 10744 19456 10750 19508
rect 12894 19456 12900 19508
rect 12952 19496 12958 19508
rect 12989 19499 13047 19505
rect 12989 19496 13001 19499
rect 12952 19468 13001 19496
rect 12952 19456 12958 19468
rect 12989 19465 13001 19468
rect 13035 19465 13047 19499
rect 12989 19459 13047 19465
rect 16206 19456 16212 19508
rect 16264 19496 16270 19508
rect 17037 19499 17095 19505
rect 17037 19496 17049 19499
rect 16264 19468 17049 19496
rect 16264 19456 16270 19468
rect 17037 19465 17049 19468
rect 17083 19465 17095 19499
rect 17037 19459 17095 19465
rect 17494 19456 17500 19508
rect 17552 19496 17558 19508
rect 18141 19499 18199 19505
rect 18141 19496 18153 19499
rect 17552 19468 18153 19496
rect 17552 19456 17558 19468
rect 18141 19465 18153 19468
rect 18187 19465 18199 19499
rect 18141 19459 18199 19465
rect 4614 19388 4620 19440
rect 4672 19388 4678 19440
rect 12434 19388 12440 19440
rect 12492 19428 12498 19440
rect 13722 19428 13728 19440
rect 12492 19400 13728 19428
rect 12492 19388 12498 19400
rect 12912 19372 12940 19400
rect 13722 19388 13728 19400
rect 13780 19428 13786 19440
rect 15102 19428 15108 19440
rect 13780 19400 15108 19428
rect 13780 19388 13786 19400
rect 2961 19363 3019 19369
rect 2961 19329 2973 19363
rect 3007 19360 3019 19363
rect 4154 19360 4160 19372
rect 3007 19332 4160 19360
rect 3007 19329 3019 19332
rect 2961 19323 3019 19329
rect 4154 19320 4160 19332
rect 4212 19320 4218 19372
rect 4338 19320 4344 19372
rect 4396 19360 4402 19372
rect 7650 19360 7656 19372
rect 4396 19332 7656 19360
rect 4396 19320 4402 19332
rect 7650 19320 7656 19332
rect 7708 19320 7714 19372
rect 8202 19320 8208 19372
rect 8260 19320 8266 19372
rect 8472 19363 8530 19369
rect 8472 19329 8484 19363
rect 8518 19360 8530 19363
rect 8518 19332 10180 19360
rect 8518 19329 8530 19332
rect 8472 19323 8530 19329
rect 3237 19295 3295 19301
rect 3237 19261 3249 19295
rect 3283 19292 3295 19295
rect 5258 19292 5264 19304
rect 3283 19264 5264 19292
rect 3283 19261 3295 19264
rect 3237 19255 3295 19261
rect 5258 19252 5264 19264
rect 5316 19252 5322 19304
rect 10152 19301 10180 19332
rect 11330 19320 11336 19372
rect 11388 19360 11394 19372
rect 11698 19360 11704 19372
rect 11388 19332 11704 19360
rect 11388 19320 11394 19332
rect 11698 19320 11704 19332
rect 11756 19360 11762 19372
rect 12618 19360 12624 19372
rect 11756 19332 12624 19360
rect 11756 19320 11762 19332
rect 12618 19320 12624 19332
rect 12676 19320 12682 19372
rect 12894 19320 12900 19372
rect 12952 19320 12958 19372
rect 14476 19369 14504 19400
rect 15102 19388 15108 19400
rect 15160 19388 15166 19440
rect 18156 19428 18184 19459
rect 18506 19456 18512 19508
rect 18564 19496 18570 19508
rect 18782 19496 18788 19508
rect 18564 19468 18788 19496
rect 18564 19456 18570 19468
rect 18782 19456 18788 19468
rect 18840 19456 18846 19508
rect 22002 19456 22008 19508
rect 22060 19496 22066 19508
rect 22060 19456 22094 19496
rect 18598 19428 18604 19440
rect 18156 19400 18604 19428
rect 18598 19388 18604 19400
rect 18656 19388 18662 19440
rect 18874 19388 18880 19440
rect 18932 19428 18938 19440
rect 22066 19428 22094 19456
rect 22189 19431 22247 19437
rect 22189 19428 22201 19431
rect 18932 19400 19840 19428
rect 22066 19400 22201 19428
rect 18932 19388 18938 19400
rect 14461 19363 14519 19369
rect 14461 19329 14473 19363
rect 14507 19329 14519 19363
rect 14461 19323 14519 19329
rect 14550 19320 14556 19372
rect 14608 19360 14614 19372
rect 14608 19332 16528 19360
rect 14608 19320 14614 19332
rect 10137 19295 10195 19301
rect 10137 19261 10149 19295
rect 10183 19292 10195 19295
rect 12434 19292 12440 19304
rect 10183 19264 12440 19292
rect 10183 19261 10195 19264
rect 10137 19255 10195 19261
rect 12434 19252 12440 19264
rect 12492 19252 12498 19304
rect 12526 19252 12532 19304
rect 12584 19252 12590 19304
rect 12713 19295 12771 19301
rect 12713 19261 12725 19295
rect 12759 19261 12771 19295
rect 12713 19255 12771 19261
rect 12813 19295 12871 19301
rect 12813 19261 12825 19295
rect 12859 19292 12871 19295
rect 12859 19264 13584 19292
rect 12859 19261 12871 19264
rect 12813 19255 12871 19261
rect 12727 19224 12755 19255
rect 13556 19236 13584 19264
rect 14734 19252 14740 19304
rect 14792 19252 14798 19304
rect 15381 19295 15439 19301
rect 15381 19261 15393 19295
rect 15427 19292 15439 19295
rect 16206 19292 16212 19304
rect 15427 19264 16212 19292
rect 15427 19261 15439 19264
rect 15381 19255 15439 19261
rect 16206 19252 16212 19264
rect 16264 19252 16270 19304
rect 16500 19292 16528 19332
rect 17328 19332 17632 19360
rect 17126 19292 17132 19304
rect 16500 19264 17132 19292
rect 17126 19252 17132 19264
rect 17184 19252 17190 19304
rect 17218 19252 17224 19304
rect 17276 19252 17282 19304
rect 17328 19301 17356 19332
rect 17313 19295 17371 19301
rect 17313 19261 17325 19295
rect 17359 19261 17371 19295
rect 17313 19255 17371 19261
rect 17402 19252 17408 19304
rect 17460 19252 17466 19304
rect 17497 19295 17555 19301
rect 17497 19261 17509 19295
rect 17543 19261 17555 19295
rect 17604 19292 17632 19332
rect 17954 19320 17960 19372
rect 18012 19360 18018 19372
rect 18325 19363 18383 19369
rect 18325 19360 18337 19363
rect 18012 19332 18337 19360
rect 18012 19320 18018 19332
rect 18325 19329 18337 19332
rect 18371 19329 18383 19363
rect 19521 19363 19579 19369
rect 18325 19323 18383 19329
rect 18432 19332 18644 19360
rect 18432 19292 18460 19332
rect 17604 19264 18460 19292
rect 17497 19255 17555 19261
rect 12986 19224 12992 19236
rect 12727 19196 12992 19224
rect 12986 19184 12992 19196
rect 13044 19184 13050 19236
rect 13538 19184 13544 19236
rect 13596 19184 13602 19236
rect 13998 19184 14004 19236
rect 14056 19224 14062 19236
rect 14645 19227 14703 19233
rect 14645 19224 14657 19227
rect 14056 19196 14657 19224
rect 14056 19184 14062 19196
rect 14645 19193 14657 19196
rect 14691 19193 14703 19227
rect 14645 19187 14703 19193
rect 16022 19184 16028 19236
rect 16080 19224 16086 19236
rect 17420 19224 17448 19252
rect 16080 19196 17448 19224
rect 17512 19224 17540 19255
rect 18506 19252 18512 19304
rect 18564 19252 18570 19304
rect 18616 19292 18644 19332
rect 19521 19329 19533 19363
rect 19567 19360 19579 19363
rect 19610 19360 19616 19372
rect 19567 19332 19616 19360
rect 19567 19329 19579 19332
rect 19521 19323 19579 19329
rect 19610 19320 19616 19332
rect 19668 19320 19674 19372
rect 19702 19320 19708 19372
rect 19760 19320 19766 19372
rect 19812 19369 19840 19400
rect 22189 19397 22201 19400
rect 22235 19397 22247 19431
rect 22189 19391 22247 19397
rect 19797 19363 19855 19369
rect 19797 19329 19809 19363
rect 19843 19329 19855 19363
rect 19797 19323 19855 19329
rect 20070 19320 20076 19372
rect 20128 19360 20134 19372
rect 22005 19363 22063 19369
rect 22005 19360 22017 19363
rect 20128 19332 22017 19360
rect 20128 19320 20134 19332
rect 22005 19329 22017 19332
rect 22051 19329 22063 19363
rect 22005 19323 22063 19329
rect 21174 19292 21180 19304
rect 18616 19264 21180 19292
rect 21174 19252 21180 19264
rect 21232 19252 21238 19304
rect 19426 19224 19432 19236
rect 17512 19196 19432 19224
rect 16080 19184 16086 19196
rect 19426 19184 19432 19196
rect 19484 19184 19490 19236
rect 14550 19116 14556 19168
rect 14608 19116 14614 19168
rect 14826 19116 14832 19168
rect 14884 19156 14890 19168
rect 15562 19156 15568 19168
rect 14884 19128 15568 19156
rect 14884 19116 14890 19128
rect 15562 19116 15568 19128
rect 15620 19156 15626 19168
rect 15841 19159 15899 19165
rect 15841 19156 15853 19159
rect 15620 19128 15853 19156
rect 15620 19116 15626 19128
rect 15841 19125 15853 19128
rect 15887 19125 15899 19159
rect 15841 19119 15899 19125
rect 15930 19116 15936 19168
rect 15988 19156 15994 19168
rect 19337 19159 19395 19165
rect 19337 19156 19349 19159
rect 15988 19128 19349 19156
rect 15988 19116 15994 19128
rect 19337 19125 19349 19128
rect 19383 19125 19395 19159
rect 19337 19119 19395 19125
rect 22278 19116 22284 19168
rect 22336 19116 22342 19168
rect 1104 19066 23828 19088
rect 1104 19014 3790 19066
rect 3842 19014 3854 19066
rect 3906 19014 3918 19066
rect 3970 19014 3982 19066
rect 4034 19014 4046 19066
rect 4098 19014 9471 19066
rect 9523 19014 9535 19066
rect 9587 19014 9599 19066
rect 9651 19014 9663 19066
rect 9715 19014 9727 19066
rect 9779 19014 15152 19066
rect 15204 19014 15216 19066
rect 15268 19014 15280 19066
rect 15332 19014 15344 19066
rect 15396 19014 15408 19066
rect 15460 19014 20833 19066
rect 20885 19014 20897 19066
rect 20949 19014 20961 19066
rect 21013 19014 21025 19066
rect 21077 19014 21089 19066
rect 21141 19014 23828 19066
rect 1104 18992 23828 19014
rect 5810 18912 5816 18964
rect 5868 18912 5874 18964
rect 7650 18912 7656 18964
rect 7708 18912 7714 18964
rect 13814 18912 13820 18964
rect 13872 18952 13878 18964
rect 14277 18955 14335 18961
rect 14277 18952 14289 18955
rect 13872 18924 14289 18952
rect 13872 18912 13878 18924
rect 14277 18921 14289 18924
rect 14323 18921 14335 18955
rect 14277 18915 14335 18921
rect 14550 18912 14556 18964
rect 14608 18952 14614 18964
rect 16577 18955 16635 18961
rect 16577 18952 16589 18955
rect 14608 18924 16589 18952
rect 14608 18912 14614 18924
rect 16577 18921 16589 18924
rect 16623 18921 16635 18955
rect 16577 18915 16635 18921
rect 18874 18912 18880 18964
rect 18932 18912 18938 18964
rect 19426 18912 19432 18964
rect 19484 18912 19490 18964
rect 12710 18844 12716 18896
rect 12768 18884 12774 18896
rect 16022 18884 16028 18896
rect 12768 18856 16028 18884
rect 12768 18844 12774 18856
rect 16022 18844 16028 18856
rect 16080 18844 16086 18896
rect 18690 18884 18696 18896
rect 16132 18856 18696 18884
rect 2038 18776 2044 18828
rect 2096 18776 2102 18828
rect 12618 18776 12624 18828
rect 12676 18816 12682 18828
rect 12897 18819 12955 18825
rect 12897 18816 12909 18819
rect 12676 18788 12909 18816
rect 12676 18776 12682 18788
rect 12897 18785 12909 18788
rect 12943 18785 12955 18819
rect 12897 18779 12955 18785
rect 12986 18776 12992 18828
rect 13044 18816 13050 18828
rect 16132 18816 16160 18856
rect 13044 18788 16160 18816
rect 16393 18819 16451 18825
rect 13044 18776 13050 18788
rect 16393 18785 16405 18819
rect 16439 18816 16451 18819
rect 17218 18816 17224 18828
rect 16439 18788 17224 18816
rect 16439 18785 16451 18788
rect 16393 18779 16451 18785
rect 17218 18776 17224 18788
rect 17276 18776 17282 18828
rect 18506 18816 18512 18828
rect 18156 18788 18512 18816
rect 5810 18708 5816 18760
rect 5868 18748 5874 18760
rect 6365 18751 6423 18757
rect 6365 18748 6377 18751
rect 5868 18720 6377 18748
rect 5868 18708 5874 18720
rect 6365 18717 6377 18720
rect 6411 18717 6423 18751
rect 6365 18711 6423 18717
rect 9122 18708 9128 18760
rect 9180 18708 9186 18760
rect 12802 18708 12808 18760
rect 12860 18708 12866 18760
rect 13078 18708 13084 18760
rect 13136 18708 13142 18760
rect 14458 18708 14464 18760
rect 14516 18708 14522 18760
rect 14921 18751 14979 18757
rect 14921 18717 14933 18751
rect 14967 18748 14979 18751
rect 16758 18748 16764 18760
rect 14967 18720 16764 18748
rect 14967 18717 14979 18720
rect 14921 18711 14979 18717
rect 16758 18708 16764 18720
rect 16816 18708 16822 18760
rect 16853 18751 16911 18757
rect 16853 18717 16865 18751
rect 16899 18748 16911 18751
rect 18156 18748 18184 18788
rect 18506 18776 18512 18788
rect 18564 18776 18570 18828
rect 16899 18720 18184 18748
rect 16899 18717 16911 18720
rect 16853 18711 16911 18717
rect 18230 18708 18236 18760
rect 18288 18708 18294 18760
rect 18414 18757 18420 18760
rect 18381 18751 18420 18757
rect 18381 18717 18393 18751
rect 18381 18711 18420 18717
rect 18414 18708 18420 18711
rect 18472 18708 18478 18760
rect 18616 18757 18644 18856
rect 18690 18844 18696 18856
rect 18748 18844 18754 18896
rect 19518 18776 19524 18828
rect 19576 18816 19582 18828
rect 19576 18788 19840 18816
rect 19576 18776 19582 18788
rect 18601 18751 18659 18757
rect 18601 18717 18613 18751
rect 18647 18717 18659 18751
rect 18601 18711 18659 18717
rect 18739 18751 18797 18757
rect 18739 18717 18751 18751
rect 18785 18748 18797 18751
rect 18874 18748 18880 18760
rect 18785 18720 18880 18748
rect 18785 18717 18797 18720
rect 18739 18711 18797 18717
rect 18874 18708 18880 18720
rect 18932 18708 18938 18760
rect 19812 18757 19840 18788
rect 19705 18751 19763 18757
rect 19705 18717 19717 18751
rect 19751 18717 19763 18751
rect 19705 18711 19763 18717
rect 19797 18751 19855 18757
rect 19797 18717 19809 18751
rect 19843 18717 19855 18751
rect 19797 18711 19855 18717
rect 19889 18751 19947 18757
rect 19889 18717 19901 18751
rect 19935 18748 19947 18751
rect 19978 18748 19984 18760
rect 19935 18720 19984 18748
rect 19935 18717 19947 18720
rect 19889 18711 19947 18717
rect 2308 18683 2366 18689
rect 2308 18649 2320 18683
rect 2354 18680 2366 18683
rect 3326 18680 3332 18692
rect 2354 18652 3332 18680
rect 2354 18649 2366 18652
rect 2308 18643 2366 18649
rect 3326 18640 3332 18652
rect 3384 18640 3390 18692
rect 9392 18683 9450 18689
rect 9392 18649 9404 18683
rect 9438 18680 9450 18683
rect 12066 18680 12072 18692
rect 9438 18652 12072 18680
rect 9438 18649 9450 18652
rect 9392 18643 9450 18649
rect 12066 18640 12072 18652
rect 12124 18640 12130 18692
rect 14550 18640 14556 18692
rect 14608 18640 14614 18692
rect 14642 18640 14648 18692
rect 14700 18640 14706 18692
rect 14763 18683 14821 18689
rect 14763 18649 14775 18683
rect 14809 18680 14821 18683
rect 15102 18680 15108 18692
rect 14809 18652 15108 18680
rect 14809 18649 14821 18652
rect 14763 18643 14821 18649
rect 15102 18640 15108 18652
rect 15160 18640 15166 18692
rect 17310 18640 17316 18692
rect 17368 18680 17374 18692
rect 18509 18683 18567 18689
rect 18509 18680 18521 18683
rect 17368 18652 18521 18680
rect 17368 18640 17374 18652
rect 18509 18649 18521 18652
rect 18555 18649 18567 18683
rect 19720 18680 19748 18711
rect 19978 18708 19984 18720
rect 20036 18708 20042 18760
rect 20073 18751 20131 18757
rect 20073 18717 20085 18751
rect 20119 18748 20131 18751
rect 20438 18748 20444 18760
rect 20119 18720 20444 18748
rect 20119 18717 20131 18720
rect 20073 18711 20131 18717
rect 20438 18708 20444 18720
rect 20496 18748 20502 18760
rect 20533 18751 20591 18757
rect 20533 18748 20545 18751
rect 20496 18720 20545 18748
rect 20496 18708 20502 18720
rect 20533 18717 20545 18720
rect 20579 18717 20591 18751
rect 20533 18711 20591 18717
rect 19720 18652 19840 18680
rect 18509 18643 18567 18649
rect 19812 18624 19840 18652
rect 3421 18615 3479 18621
rect 3421 18581 3433 18615
rect 3467 18612 3479 18615
rect 5442 18612 5448 18624
rect 3467 18584 5448 18612
rect 3467 18581 3479 18584
rect 3421 18575 3479 18581
rect 5442 18572 5448 18584
rect 5500 18572 5506 18624
rect 10505 18615 10563 18621
rect 10505 18581 10517 18615
rect 10551 18612 10563 18615
rect 10962 18612 10968 18624
rect 10551 18584 10968 18612
rect 10551 18581 10563 18584
rect 10505 18575 10563 18581
rect 10962 18572 10968 18584
rect 11020 18572 11026 18624
rect 12526 18572 12532 18624
rect 12584 18612 12590 18624
rect 13170 18612 13176 18624
rect 12584 18584 13176 18612
rect 12584 18572 12590 18584
rect 13170 18572 13176 18584
rect 13228 18572 13234 18624
rect 13262 18572 13268 18624
rect 13320 18572 13326 18624
rect 13906 18572 13912 18624
rect 13964 18612 13970 18624
rect 15381 18615 15439 18621
rect 15381 18612 15393 18615
rect 13964 18584 15393 18612
rect 13964 18572 13970 18584
rect 15381 18581 15393 18584
rect 15427 18581 15439 18615
rect 15381 18575 15439 18581
rect 16761 18615 16819 18621
rect 16761 18581 16773 18615
rect 16807 18612 16819 18615
rect 17586 18612 17592 18624
rect 16807 18584 17592 18612
rect 16807 18581 16819 18584
rect 16761 18575 16819 18581
rect 17586 18572 17592 18584
rect 17644 18612 17650 18624
rect 19794 18612 19800 18624
rect 17644 18584 19800 18612
rect 17644 18572 17650 18584
rect 19794 18572 19800 18584
rect 19852 18612 19858 18624
rect 20162 18612 20168 18624
rect 19852 18584 20168 18612
rect 19852 18572 19858 18584
rect 20162 18572 20168 18584
rect 20220 18572 20226 18624
rect 1104 18522 23987 18544
rect 1104 18470 6630 18522
rect 6682 18470 6694 18522
rect 6746 18470 6758 18522
rect 6810 18470 6822 18522
rect 6874 18470 6886 18522
rect 6938 18470 12311 18522
rect 12363 18470 12375 18522
rect 12427 18470 12439 18522
rect 12491 18470 12503 18522
rect 12555 18470 12567 18522
rect 12619 18470 17992 18522
rect 18044 18470 18056 18522
rect 18108 18470 18120 18522
rect 18172 18470 18184 18522
rect 18236 18470 18248 18522
rect 18300 18470 23673 18522
rect 23725 18470 23737 18522
rect 23789 18470 23801 18522
rect 23853 18470 23865 18522
rect 23917 18470 23929 18522
rect 23981 18470 23987 18522
rect 1104 18448 23987 18470
rect 9122 18368 9128 18420
rect 9180 18368 9186 18420
rect 12066 18368 12072 18420
rect 12124 18368 12130 18420
rect 13725 18411 13783 18417
rect 13725 18377 13737 18411
rect 13771 18408 13783 18411
rect 13906 18408 13912 18420
rect 13771 18380 13912 18408
rect 13771 18377 13783 18380
rect 13725 18371 13783 18377
rect 13906 18368 13912 18380
rect 13964 18368 13970 18420
rect 14093 18411 14151 18417
rect 14093 18377 14105 18411
rect 14139 18408 14151 18411
rect 15102 18408 15108 18420
rect 14139 18380 15108 18408
rect 14139 18377 14151 18380
rect 14093 18371 14151 18377
rect 15102 18368 15108 18380
rect 15160 18368 15166 18420
rect 15197 18411 15255 18417
rect 15197 18377 15209 18411
rect 15243 18408 15255 18411
rect 15470 18408 15476 18420
rect 15243 18380 15476 18408
rect 15243 18377 15255 18380
rect 15197 18371 15255 18377
rect 15470 18368 15476 18380
rect 15528 18368 15534 18420
rect 16758 18368 16764 18420
rect 16816 18408 16822 18420
rect 16945 18411 17003 18417
rect 16945 18408 16957 18411
rect 16816 18380 16957 18408
rect 16816 18368 16822 18380
rect 16945 18377 16957 18380
rect 16991 18377 17003 18411
rect 17494 18408 17500 18420
rect 16945 18371 17003 18377
rect 17052 18380 17500 18408
rect 3320 18343 3378 18349
rect 3320 18309 3332 18343
rect 3366 18340 3378 18343
rect 3510 18340 3516 18352
rect 3366 18312 3516 18340
rect 3366 18309 3378 18312
rect 3320 18303 3378 18309
rect 3510 18300 3516 18312
rect 3568 18300 3574 18352
rect 12986 18340 12992 18352
rect 12268 18312 12992 18340
rect 7650 18232 7656 18284
rect 7708 18272 7714 18284
rect 12268 18281 12296 18312
rect 12986 18300 12992 18312
rect 13044 18300 13050 18352
rect 13262 18300 13268 18352
rect 13320 18340 13326 18352
rect 14553 18343 14611 18349
rect 14553 18340 14565 18343
rect 13320 18312 14565 18340
rect 13320 18300 13326 18312
rect 14553 18309 14565 18312
rect 14599 18309 14611 18343
rect 14553 18303 14611 18309
rect 14645 18343 14703 18349
rect 14645 18309 14657 18343
rect 14691 18340 14703 18343
rect 14691 18312 15516 18340
rect 14691 18309 14703 18312
rect 14645 18303 14703 18309
rect 7837 18275 7895 18281
rect 7837 18272 7849 18275
rect 7708 18244 7849 18272
rect 7708 18232 7714 18244
rect 7837 18241 7849 18244
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 12253 18275 12311 18281
rect 12253 18241 12265 18275
rect 12299 18241 12311 18275
rect 12253 18235 12311 18241
rect 12345 18275 12403 18281
rect 12345 18241 12357 18275
rect 12391 18241 12403 18275
rect 12345 18235 12403 18241
rect 12621 18275 12679 18281
rect 12621 18241 12633 18275
rect 12667 18272 12679 18275
rect 12710 18272 12716 18284
rect 12667 18244 12716 18272
rect 12667 18241 12679 18244
rect 12621 18235 12679 18241
rect 3050 18164 3056 18216
rect 3108 18164 3114 18216
rect 12066 18164 12072 18216
rect 12124 18204 12130 18216
rect 12360 18204 12388 18235
rect 12710 18232 12716 18244
rect 12768 18232 12774 18284
rect 13173 18275 13231 18281
rect 13173 18241 13185 18275
rect 13219 18272 13231 18275
rect 13538 18272 13544 18284
rect 13219 18244 13544 18272
rect 13219 18241 13231 18244
rect 13173 18235 13231 18241
rect 13538 18232 13544 18244
rect 13596 18232 13602 18284
rect 13633 18278 13691 18281
rect 13633 18275 13860 18278
rect 13633 18241 13645 18275
rect 13679 18250 13860 18275
rect 13679 18241 13691 18250
rect 13633 18235 13691 18241
rect 12124 18176 12388 18204
rect 12529 18207 12587 18213
rect 12124 18164 12130 18176
rect 12529 18173 12541 18207
rect 12575 18204 12587 18207
rect 13832 18204 13860 18250
rect 13909 18275 13967 18281
rect 13909 18241 13921 18275
rect 13955 18272 13967 18275
rect 13955 18244 14228 18272
rect 13955 18241 13967 18244
rect 13909 18235 13967 18241
rect 14090 18204 14096 18216
rect 12575 18176 13584 18204
rect 13832 18176 14096 18204
rect 12575 18173 12587 18176
rect 12529 18167 12587 18173
rect 4433 18071 4491 18077
rect 4433 18037 4445 18071
rect 4479 18068 4491 18071
rect 5074 18068 5080 18080
rect 4479 18040 5080 18068
rect 4479 18037 4491 18040
rect 4433 18031 4491 18037
rect 5074 18028 5080 18040
rect 5132 18028 5138 18080
rect 13556 18068 13584 18176
rect 14090 18164 14096 18176
rect 14148 18164 14154 18216
rect 14200 18148 14228 18244
rect 14274 18232 14280 18284
rect 14332 18272 14338 18284
rect 14660 18272 14688 18303
rect 15488 18284 15516 18312
rect 14332 18244 14688 18272
rect 14332 18232 14338 18244
rect 14826 18232 14832 18284
rect 14884 18272 14890 18284
rect 14921 18275 14979 18281
rect 14921 18272 14933 18275
rect 14884 18244 14933 18272
rect 14884 18232 14890 18244
rect 14921 18241 14933 18244
rect 14967 18241 14979 18275
rect 14921 18235 14979 18241
rect 15470 18232 15476 18284
rect 15528 18232 15534 18284
rect 16022 18232 16028 18284
rect 16080 18272 16086 18284
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 16080 18244 16865 18272
rect 16080 18232 16086 18244
rect 16853 18241 16865 18244
rect 16899 18272 16911 18275
rect 17052 18272 17080 18380
rect 17494 18368 17500 18380
rect 17552 18408 17558 18420
rect 18322 18408 18328 18420
rect 17552 18380 18328 18408
rect 17552 18368 17558 18380
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 18414 18368 18420 18420
rect 18472 18408 18478 18420
rect 18969 18411 19027 18417
rect 18969 18408 18981 18411
rect 18472 18380 18981 18408
rect 18472 18368 18478 18380
rect 18969 18377 18981 18380
rect 19015 18377 19027 18411
rect 18969 18371 19027 18377
rect 19334 18368 19340 18420
rect 19392 18408 19398 18420
rect 19521 18411 19579 18417
rect 19521 18408 19533 18411
rect 19392 18380 19533 18408
rect 19392 18368 19398 18380
rect 19521 18377 19533 18380
rect 19567 18377 19579 18411
rect 19521 18371 19579 18377
rect 17402 18300 17408 18352
rect 17460 18340 17466 18352
rect 19794 18340 19800 18352
rect 17460 18312 17908 18340
rect 17460 18300 17466 18312
rect 16899 18244 17080 18272
rect 17221 18275 17279 18281
rect 16899 18241 16911 18244
rect 16853 18235 16911 18241
rect 17221 18241 17233 18275
rect 17267 18272 17279 18275
rect 17770 18272 17776 18284
rect 17267 18244 17776 18272
rect 17267 18241 17279 18244
rect 17221 18235 17279 18241
rect 17770 18232 17776 18244
rect 17828 18232 17834 18284
rect 15010 18164 15016 18216
rect 15068 18164 15074 18216
rect 15102 18164 15108 18216
rect 15160 18204 15166 18216
rect 17405 18207 17463 18213
rect 17405 18204 17417 18207
rect 15160 18176 17417 18204
rect 15160 18164 15166 18176
rect 17405 18173 17417 18176
rect 17451 18173 17463 18207
rect 17880 18204 17908 18312
rect 19720 18312 19800 18340
rect 19720 18281 19748 18312
rect 19794 18300 19800 18312
rect 19852 18340 19858 18352
rect 20254 18340 20260 18352
rect 19852 18312 20260 18340
rect 19852 18300 19858 18312
rect 20254 18300 20260 18312
rect 20312 18300 20318 18352
rect 18049 18275 18107 18281
rect 18049 18241 18061 18275
rect 18095 18272 18107 18275
rect 19705 18275 19763 18281
rect 18095 18244 19656 18272
rect 18095 18241 18107 18244
rect 18049 18235 18107 18241
rect 18325 18207 18383 18213
rect 18325 18204 18337 18207
rect 17880 18176 18337 18204
rect 17405 18167 17463 18173
rect 18325 18173 18337 18176
rect 18371 18173 18383 18207
rect 19628 18204 19656 18244
rect 19705 18241 19717 18275
rect 19751 18241 19763 18275
rect 19705 18235 19763 18241
rect 19886 18232 19892 18284
rect 19944 18232 19950 18284
rect 19981 18275 20039 18281
rect 19981 18241 19993 18275
rect 20027 18272 20039 18275
rect 20070 18272 20076 18284
rect 20027 18244 20076 18272
rect 20027 18241 20039 18244
rect 19981 18235 20039 18241
rect 20070 18232 20076 18244
rect 20128 18232 20134 18284
rect 20714 18204 20720 18216
rect 19628 18176 20720 18204
rect 18325 18167 18383 18173
rect 14182 18096 14188 18148
rect 14240 18136 14246 18148
rect 17420 18136 17448 18167
rect 20714 18164 20720 18176
rect 20772 18164 20778 18216
rect 17954 18136 17960 18148
rect 14240 18108 16344 18136
rect 17420 18108 17960 18136
rect 14240 18096 14246 18108
rect 13998 18068 14004 18080
rect 13556 18040 14004 18068
rect 13998 18028 14004 18040
rect 14056 18028 14062 18080
rect 14734 18028 14740 18080
rect 14792 18068 14798 18080
rect 15102 18068 15108 18080
rect 14792 18040 15108 18068
rect 14792 18028 14798 18040
rect 15102 18028 15108 18040
rect 15160 18028 15166 18080
rect 15470 18028 15476 18080
rect 15528 18068 15534 18080
rect 16316 18077 16344 18108
rect 17954 18096 17960 18108
rect 18012 18136 18018 18148
rect 19150 18136 19156 18148
rect 18012 18108 19156 18136
rect 18012 18096 18018 18108
rect 19150 18096 19156 18108
rect 19208 18096 19214 18148
rect 15657 18071 15715 18077
rect 15657 18068 15669 18071
rect 15528 18040 15669 18068
rect 15528 18028 15534 18040
rect 15657 18037 15669 18040
rect 15703 18037 15715 18071
rect 15657 18031 15715 18037
rect 16301 18071 16359 18077
rect 16301 18037 16313 18071
rect 16347 18068 16359 18071
rect 17402 18068 17408 18080
rect 16347 18040 17408 18068
rect 16347 18037 16359 18040
rect 16301 18031 16359 18037
rect 17402 18028 17408 18040
rect 17460 18028 17466 18080
rect 17862 18028 17868 18080
rect 17920 18028 17926 18080
rect 18233 18071 18291 18077
rect 18233 18037 18245 18071
rect 18279 18068 18291 18071
rect 18322 18068 18328 18080
rect 18279 18040 18328 18068
rect 18279 18037 18291 18040
rect 18233 18031 18291 18037
rect 18322 18028 18328 18040
rect 18380 18028 18386 18080
rect 1104 17978 23828 18000
rect 1104 17926 3790 17978
rect 3842 17926 3854 17978
rect 3906 17926 3918 17978
rect 3970 17926 3982 17978
rect 4034 17926 4046 17978
rect 4098 17926 9471 17978
rect 9523 17926 9535 17978
rect 9587 17926 9599 17978
rect 9651 17926 9663 17978
rect 9715 17926 9727 17978
rect 9779 17926 15152 17978
rect 15204 17926 15216 17978
rect 15268 17926 15280 17978
rect 15332 17926 15344 17978
rect 15396 17926 15408 17978
rect 15460 17926 20833 17978
rect 20885 17926 20897 17978
rect 20949 17926 20961 17978
rect 21013 17926 21025 17978
rect 21077 17926 21089 17978
rect 21141 17926 23828 17978
rect 1104 17904 23828 17926
rect 11698 17824 11704 17876
rect 11756 17824 11762 17876
rect 13170 17824 13176 17876
rect 13228 17824 13234 17876
rect 13262 17824 13268 17876
rect 13320 17864 13326 17876
rect 17497 17867 17555 17873
rect 17497 17864 17509 17867
rect 13320 17836 17509 17864
rect 13320 17824 13326 17836
rect 17497 17833 17509 17836
rect 17543 17833 17555 17867
rect 17497 17827 17555 17833
rect 20438 17824 20444 17876
rect 20496 17864 20502 17876
rect 21453 17867 21511 17873
rect 21453 17864 21465 17867
rect 20496 17836 21465 17864
rect 20496 17824 20502 17836
rect 21453 17833 21465 17836
rect 21499 17833 21511 17867
rect 21453 17827 21511 17833
rect 11716 17728 11744 17824
rect 12713 17799 12771 17805
rect 12713 17765 12725 17799
rect 12759 17796 12771 17799
rect 14550 17796 14556 17808
rect 12759 17768 14556 17796
rect 12759 17765 12771 17768
rect 12713 17759 12771 17765
rect 14550 17756 14556 17768
rect 14608 17756 14614 17808
rect 15930 17756 15936 17808
rect 15988 17796 15994 17808
rect 16761 17799 16819 17805
rect 16761 17796 16773 17799
rect 15988 17768 16773 17796
rect 15988 17756 15994 17768
rect 16761 17765 16773 17768
rect 16807 17796 16819 17799
rect 17310 17796 17316 17808
rect 16807 17768 17316 17796
rect 16807 17765 16819 17768
rect 16761 17759 16819 17765
rect 17310 17756 17316 17768
rect 17368 17756 17374 17808
rect 13538 17728 13544 17740
rect 11716 17700 12388 17728
rect 6546 17620 6552 17672
rect 6604 17660 6610 17672
rect 7101 17663 7159 17669
rect 7101 17660 7113 17663
rect 6604 17632 7113 17660
rect 6604 17620 6610 17632
rect 7101 17629 7113 17632
rect 7147 17629 7159 17663
rect 7101 17623 7159 17629
rect 9122 17620 9128 17672
rect 9180 17620 9186 17672
rect 11149 17663 11207 17669
rect 11149 17629 11161 17663
rect 11195 17660 11207 17663
rect 11606 17660 11612 17672
rect 11195 17632 11612 17660
rect 11195 17629 11207 17632
rect 11149 17623 11207 17629
rect 11606 17620 11612 17632
rect 11664 17620 11670 17672
rect 11882 17620 11888 17672
rect 11940 17660 11946 17672
rect 12360 17669 12388 17700
rect 12544 17700 13544 17728
rect 12544 17669 12572 17700
rect 13538 17688 13544 17700
rect 13596 17728 13602 17740
rect 14182 17728 14188 17740
rect 13596 17700 14188 17728
rect 13596 17688 13602 17700
rect 14182 17688 14188 17700
rect 14240 17688 14246 17740
rect 14642 17688 14648 17740
rect 14700 17728 14706 17740
rect 14829 17731 14887 17737
rect 14829 17728 14841 17731
rect 14700 17700 14841 17728
rect 14700 17688 14706 17700
rect 14829 17697 14841 17700
rect 14875 17728 14887 17731
rect 15194 17728 15200 17740
rect 14875 17700 15200 17728
rect 14875 17697 14887 17700
rect 14829 17691 14887 17697
rect 15194 17688 15200 17700
rect 15252 17728 15258 17740
rect 16022 17728 16028 17740
rect 15252 17700 16028 17728
rect 15252 17688 15258 17700
rect 16022 17688 16028 17700
rect 16080 17688 16086 17740
rect 17586 17728 17592 17740
rect 16592 17700 17592 17728
rect 16592 17672 16620 17700
rect 17586 17688 17592 17700
rect 17644 17688 17650 17740
rect 12253 17663 12311 17669
rect 12253 17660 12265 17663
rect 11940 17632 12265 17660
rect 11940 17620 11946 17632
rect 12253 17629 12265 17632
rect 12299 17629 12311 17663
rect 12253 17623 12311 17629
rect 12345 17663 12403 17669
rect 12345 17629 12357 17663
rect 12391 17629 12403 17663
rect 12345 17623 12403 17629
rect 12529 17663 12587 17669
rect 12529 17629 12541 17663
rect 12575 17660 12587 17663
rect 12710 17660 12716 17672
rect 12575 17632 12716 17660
rect 12575 17629 12587 17632
rect 12529 17623 12587 17629
rect 12710 17620 12716 17632
rect 12768 17620 12774 17672
rect 13354 17620 13360 17672
rect 13412 17620 13418 17672
rect 13449 17663 13507 17669
rect 13449 17629 13461 17663
rect 13495 17629 13507 17663
rect 13449 17623 13507 17629
rect 13633 17663 13691 17669
rect 13633 17629 13645 17663
rect 13679 17660 13691 17663
rect 13814 17660 13820 17672
rect 13679 17632 13820 17660
rect 13679 17629 13691 17632
rect 13633 17623 13691 17629
rect 6856 17595 6914 17601
rect 6856 17561 6868 17595
rect 6902 17592 6914 17595
rect 7466 17592 7472 17604
rect 6902 17564 7472 17592
rect 6902 17561 6914 17564
rect 6856 17555 6914 17561
rect 7466 17552 7472 17564
rect 7524 17552 7530 17604
rect 9392 17595 9450 17601
rect 9392 17561 9404 17595
rect 9438 17592 9450 17595
rect 13464 17592 13492 17623
rect 13814 17620 13820 17632
rect 13872 17660 13878 17672
rect 14274 17660 14280 17672
rect 13872 17632 14280 17660
rect 13872 17620 13878 17632
rect 14274 17620 14280 17632
rect 14332 17620 14338 17672
rect 15010 17620 15016 17672
rect 15068 17620 15074 17672
rect 15654 17620 15660 17672
rect 15712 17620 15718 17672
rect 15933 17663 15991 17669
rect 15933 17629 15945 17663
rect 15979 17660 15991 17663
rect 16206 17660 16212 17672
rect 15979 17632 16212 17660
rect 15979 17629 15991 17632
rect 15933 17623 15991 17629
rect 16206 17620 16212 17632
rect 16264 17660 16270 17672
rect 16264 17632 16528 17660
rect 16264 17620 16270 17632
rect 13722 17592 13728 17604
rect 9438 17564 11836 17592
rect 13464 17564 13728 17592
rect 9438 17561 9450 17564
rect 9392 17555 9450 17561
rect 5721 17527 5779 17533
rect 5721 17493 5733 17527
rect 5767 17524 5779 17527
rect 6086 17524 6092 17536
rect 5767 17496 6092 17524
rect 5767 17493 5779 17496
rect 5721 17487 5779 17493
rect 6086 17484 6092 17496
rect 6144 17484 6150 17536
rect 8018 17484 8024 17536
rect 8076 17524 8082 17536
rect 8389 17527 8447 17533
rect 8389 17524 8401 17527
rect 8076 17496 8401 17524
rect 8076 17484 8082 17496
rect 8389 17493 8401 17496
rect 8435 17493 8447 17527
rect 8389 17487 8447 17493
rect 10505 17527 10563 17533
rect 10505 17493 10517 17527
rect 10551 17524 10563 17527
rect 11514 17524 11520 17536
rect 10551 17496 11520 17524
rect 10551 17493 10563 17496
rect 10505 17487 10563 17493
rect 11514 17484 11520 17496
rect 11572 17484 11578 17536
rect 11808 17524 11836 17564
rect 13722 17552 13728 17564
rect 13780 17552 13786 17604
rect 15562 17552 15568 17604
rect 15620 17592 15626 17604
rect 16393 17595 16451 17601
rect 16393 17592 16405 17595
rect 15620 17564 16405 17592
rect 15620 17552 15626 17564
rect 16393 17561 16405 17564
rect 16439 17561 16451 17595
rect 16500 17592 16528 17632
rect 16574 17620 16580 17672
rect 16632 17620 16638 17672
rect 16850 17620 16856 17672
rect 16908 17620 16914 17672
rect 17681 17663 17739 17669
rect 17681 17660 17693 17663
rect 16960 17632 17693 17660
rect 16666 17592 16672 17604
rect 16500 17564 16672 17592
rect 16393 17555 16451 17561
rect 16666 17552 16672 17564
rect 16724 17552 16730 17604
rect 14918 17524 14924 17536
rect 11808 17496 14924 17524
rect 14918 17484 14924 17496
rect 14976 17484 14982 17536
rect 15473 17527 15531 17533
rect 15473 17493 15485 17527
rect 15519 17524 15531 17527
rect 15654 17524 15660 17536
rect 15519 17496 15660 17524
rect 15519 17493 15531 17496
rect 15473 17487 15531 17493
rect 15654 17484 15660 17496
rect 15712 17484 15718 17536
rect 15841 17527 15899 17533
rect 15841 17493 15853 17527
rect 15887 17524 15899 17527
rect 16022 17524 16028 17536
rect 15887 17496 16028 17524
rect 15887 17493 15899 17496
rect 15841 17487 15899 17493
rect 16022 17484 16028 17496
rect 16080 17484 16086 17536
rect 16114 17484 16120 17536
rect 16172 17524 16178 17536
rect 16960 17524 16988 17632
rect 17681 17629 17693 17632
rect 17727 17629 17739 17663
rect 21468 17660 21496 17827
rect 22554 17824 22560 17876
rect 22612 17864 22618 17876
rect 22649 17867 22707 17873
rect 22649 17864 22661 17867
rect 22612 17836 22661 17864
rect 22612 17824 22618 17836
rect 22649 17833 22661 17836
rect 22695 17833 22707 17867
rect 22649 17827 22707 17833
rect 22005 17663 22063 17669
rect 22005 17660 22017 17663
rect 21468 17632 22017 17660
rect 17681 17623 17739 17629
rect 22005 17629 22017 17632
rect 22051 17629 22063 17663
rect 22005 17623 22063 17629
rect 22186 17620 22192 17672
rect 22244 17620 22250 17672
rect 22278 17620 22284 17672
rect 22336 17620 22342 17672
rect 22370 17620 22376 17672
rect 22428 17620 22434 17672
rect 17218 17552 17224 17604
rect 17276 17592 17282 17604
rect 17276 17564 17356 17592
rect 17276 17552 17282 17564
rect 17328 17533 17356 17564
rect 16172 17496 16988 17524
rect 17313 17527 17371 17533
rect 16172 17484 16178 17496
rect 17313 17493 17325 17527
rect 17359 17493 17371 17527
rect 17313 17487 17371 17493
rect 1104 17434 23987 17456
rect 1104 17382 6630 17434
rect 6682 17382 6694 17434
rect 6746 17382 6758 17434
rect 6810 17382 6822 17434
rect 6874 17382 6886 17434
rect 6938 17382 12311 17434
rect 12363 17382 12375 17434
rect 12427 17382 12439 17434
rect 12491 17382 12503 17434
rect 12555 17382 12567 17434
rect 12619 17382 17992 17434
rect 18044 17382 18056 17434
rect 18108 17382 18120 17434
rect 18172 17382 18184 17434
rect 18236 17382 18248 17434
rect 18300 17382 23673 17434
rect 23725 17382 23737 17434
rect 23789 17382 23801 17434
rect 23853 17382 23865 17434
rect 23917 17382 23929 17434
rect 23981 17382 23987 17434
rect 1104 17360 23987 17382
rect 11330 17280 11336 17332
rect 11388 17320 11394 17332
rect 12345 17323 12403 17329
rect 12345 17320 12357 17323
rect 11388 17292 12357 17320
rect 11388 17280 11394 17292
rect 12345 17289 12357 17292
rect 12391 17320 12403 17323
rect 12710 17320 12716 17332
rect 12391 17292 12716 17320
rect 12391 17289 12403 17292
rect 12345 17283 12403 17289
rect 12710 17280 12716 17292
rect 12768 17280 12774 17332
rect 13078 17280 13084 17332
rect 13136 17280 13142 17332
rect 13354 17280 13360 17332
rect 13412 17320 13418 17332
rect 13814 17320 13820 17332
rect 13412 17292 13820 17320
rect 13412 17280 13418 17292
rect 13814 17280 13820 17292
rect 13872 17280 13878 17332
rect 14918 17320 14924 17332
rect 14844 17292 14924 17320
rect 11882 17212 11888 17264
rect 11940 17252 11946 17264
rect 13096 17252 13124 17280
rect 14844 17261 14872 17292
rect 14918 17280 14924 17292
rect 14976 17280 14982 17332
rect 16209 17323 16267 17329
rect 16209 17289 16221 17323
rect 16255 17320 16267 17323
rect 16298 17320 16304 17332
rect 16255 17292 16304 17320
rect 16255 17289 16267 17292
rect 16209 17283 16267 17289
rect 16298 17280 16304 17292
rect 16356 17280 16362 17332
rect 16666 17280 16672 17332
rect 16724 17320 16730 17332
rect 17954 17320 17960 17332
rect 16724 17292 17960 17320
rect 16724 17280 16730 17292
rect 17954 17280 17960 17292
rect 18012 17280 18018 17332
rect 18874 17280 18880 17332
rect 18932 17280 18938 17332
rect 19337 17323 19395 17329
rect 19337 17289 19349 17323
rect 19383 17320 19395 17323
rect 19610 17320 19616 17332
rect 19383 17292 19616 17320
rect 19383 17289 19395 17292
rect 19337 17283 19395 17289
rect 19610 17280 19616 17292
rect 19668 17280 19674 17332
rect 19702 17280 19708 17332
rect 19760 17320 19766 17332
rect 19981 17323 20039 17329
rect 19981 17320 19993 17323
rect 19760 17292 19993 17320
rect 19760 17280 19766 17292
rect 19981 17289 19993 17292
rect 20027 17289 20039 17323
rect 19981 17283 20039 17289
rect 20088 17292 22232 17320
rect 13909 17255 13967 17261
rect 13909 17252 13921 17255
rect 11940 17224 13921 17252
rect 11940 17212 11946 17224
rect 2961 17187 3019 17193
rect 2961 17153 2973 17187
rect 3007 17184 3019 17187
rect 3050 17184 3056 17196
rect 3007 17156 3056 17184
rect 3007 17153 3019 17156
rect 2961 17147 3019 17153
rect 3050 17144 3056 17156
rect 3108 17144 3114 17196
rect 6816 17187 6874 17193
rect 6816 17153 6828 17187
rect 6862 17184 6874 17187
rect 7926 17184 7932 17196
rect 6862 17156 7932 17184
rect 6862 17153 6874 17156
rect 6816 17147 6874 17153
rect 7926 17144 7932 17156
rect 7984 17144 7990 17196
rect 8748 17187 8806 17193
rect 8748 17153 8760 17187
rect 8794 17184 8806 17187
rect 10594 17184 10600 17196
rect 8794 17156 10600 17184
rect 8794 17153 8806 17156
rect 8748 17147 8806 17153
rect 10594 17144 10600 17156
rect 10652 17144 10658 17196
rect 12928 17184 12956 17224
rect 13909 17221 13921 17224
rect 13955 17221 13967 17255
rect 13909 17215 13967 17221
rect 14829 17255 14887 17261
rect 14829 17221 14841 17255
rect 14875 17221 14887 17255
rect 16850 17252 16856 17264
rect 14829 17215 14887 17221
rect 15028 17224 16856 17252
rect 12992 17187 13050 17193
rect 12992 17184 13004 17187
rect 12928 17156 13004 17184
rect 12992 17153 13004 17156
rect 13038 17153 13050 17187
rect 12992 17147 13050 17153
rect 13081 17187 13139 17193
rect 13081 17153 13093 17187
rect 13127 17184 13139 17187
rect 13170 17184 13176 17196
rect 13127 17156 13176 17184
rect 13127 17153 13139 17156
rect 13081 17147 13139 17153
rect 13170 17144 13176 17156
rect 13228 17144 13234 17196
rect 13265 17187 13323 17193
rect 13265 17153 13277 17187
rect 13311 17153 13323 17187
rect 13265 17147 13323 17153
rect 2222 17076 2228 17128
rect 2280 17116 2286 17128
rect 3237 17119 3295 17125
rect 3237 17116 3249 17119
rect 2280 17088 3249 17116
rect 2280 17076 2286 17088
rect 3237 17085 3249 17088
rect 3283 17085 3295 17119
rect 3237 17079 3295 17085
rect 6546 17076 6552 17128
rect 6604 17076 6610 17128
rect 8478 17076 8484 17128
rect 8536 17076 8542 17128
rect 12802 17076 12808 17128
rect 12860 17116 12866 17128
rect 13280 17116 13308 17147
rect 13354 17144 13360 17196
rect 13412 17144 13418 17196
rect 13814 17144 13820 17196
rect 13872 17144 13878 17196
rect 13998 17144 14004 17196
rect 14056 17144 14062 17196
rect 14366 17144 14372 17196
rect 14424 17184 14430 17196
rect 14693 17187 14751 17193
rect 14693 17184 14705 17187
rect 14424 17156 14705 17184
rect 14424 17144 14430 17156
rect 14693 17153 14705 17156
rect 14739 17153 14751 17187
rect 14693 17147 14751 17153
rect 14921 17187 14979 17193
rect 14921 17153 14933 17187
rect 14967 17184 14979 17187
rect 15028 17184 15056 17224
rect 16850 17212 16856 17224
rect 16908 17252 16914 17264
rect 17129 17255 17187 17261
rect 17129 17252 17141 17255
rect 16908 17224 17141 17252
rect 16908 17212 16914 17224
rect 17129 17221 17141 17224
rect 17175 17221 17187 17255
rect 17129 17215 17187 17221
rect 17310 17212 17316 17264
rect 17368 17252 17374 17264
rect 18892 17252 18920 17280
rect 17368 17224 18920 17252
rect 17368 17212 17374 17224
rect 19150 17212 19156 17264
rect 19208 17252 19214 17264
rect 19208 17224 19564 17252
rect 19208 17212 19214 17224
rect 15194 17193 15200 17196
rect 14967 17156 15056 17184
rect 15104 17187 15162 17193
rect 14967 17153 14979 17156
rect 14921 17147 14979 17153
rect 15104 17153 15116 17187
rect 15150 17153 15162 17187
rect 15104 17147 15162 17153
rect 15190 17147 15200 17193
rect 15252 17184 15258 17196
rect 15252 17156 15290 17184
rect 14458 17116 14464 17128
rect 12860 17088 14464 17116
rect 12860 17076 12866 17088
rect 14458 17076 14464 17088
rect 14516 17076 14522 17128
rect 15119 17060 15147 17147
rect 15194 17144 15200 17147
rect 15252 17144 15258 17156
rect 16114 17144 16120 17196
rect 16172 17144 16178 17196
rect 16301 17187 16359 17193
rect 16301 17153 16313 17187
rect 16347 17184 16359 17187
rect 17037 17187 17095 17193
rect 17037 17184 17049 17187
rect 16347 17156 17049 17184
rect 16347 17153 16359 17156
rect 16301 17147 16359 17153
rect 17037 17153 17049 17156
rect 17083 17153 17095 17187
rect 17037 17147 17095 17153
rect 17221 17187 17279 17193
rect 17221 17153 17233 17187
rect 17267 17184 17279 17187
rect 18874 17184 18880 17196
rect 17267 17156 18880 17184
rect 17267 17153 17279 17156
rect 17221 17147 17279 17153
rect 17052 17116 17080 17147
rect 18874 17144 18880 17156
rect 18932 17144 18938 17196
rect 19242 17144 19248 17196
rect 19300 17144 19306 17196
rect 19536 17193 19564 17224
rect 19521 17187 19579 17193
rect 19521 17153 19533 17187
rect 19567 17153 19579 17187
rect 19521 17147 19579 17153
rect 19705 17187 19763 17193
rect 19705 17153 19717 17187
rect 19751 17184 19763 17187
rect 19794 17184 19800 17196
rect 19751 17156 19800 17184
rect 19751 17153 19763 17156
rect 19705 17147 19763 17153
rect 19794 17144 19800 17156
rect 19852 17144 19858 17196
rect 17494 17116 17500 17128
rect 17052 17088 17500 17116
rect 17494 17076 17500 17088
rect 17552 17076 17558 17128
rect 17678 17076 17684 17128
rect 17736 17116 17742 17128
rect 19613 17119 19671 17125
rect 19613 17116 19625 17119
rect 17736 17088 19625 17116
rect 17736 17076 17742 17088
rect 19613 17085 19625 17088
rect 19659 17085 19671 17119
rect 19613 17079 19671 17085
rect 12986 17008 12992 17060
rect 13044 17048 13050 17060
rect 13170 17048 13176 17060
rect 13044 17020 13176 17048
rect 13044 17008 13050 17020
rect 13170 17008 13176 17020
rect 13228 17008 13234 17060
rect 13538 17008 13544 17060
rect 13596 17048 13602 17060
rect 13596 17020 15056 17048
rect 13596 17008 13602 17020
rect 15028 16992 15056 17020
rect 15102 17008 15108 17060
rect 15160 17008 15166 17060
rect 4522 16940 4528 16992
rect 4580 16940 4586 16992
rect 7929 16983 7987 16989
rect 7929 16949 7941 16983
rect 7975 16980 7987 16983
rect 8846 16980 8852 16992
rect 7975 16952 8852 16980
rect 7975 16949 7987 16952
rect 7929 16943 7987 16949
rect 8846 16940 8852 16952
rect 8904 16940 8910 16992
rect 9861 16983 9919 16989
rect 9861 16949 9873 16983
rect 9907 16980 9919 16983
rect 10226 16980 10232 16992
rect 9907 16952 10232 16980
rect 9907 16949 9919 16952
rect 9861 16943 9919 16949
rect 10226 16940 10232 16952
rect 10284 16940 10290 16992
rect 12526 16940 12532 16992
rect 12584 16980 12590 16992
rect 12805 16983 12863 16989
rect 12805 16980 12817 16983
rect 12584 16952 12817 16980
rect 12584 16940 12590 16952
rect 12805 16949 12817 16952
rect 12851 16949 12863 16983
rect 12805 16943 12863 16949
rect 14550 16940 14556 16992
rect 14608 16940 14614 16992
rect 15010 16940 15016 16992
rect 15068 16980 15074 16992
rect 20088 16980 20116 17292
rect 22204 17193 22232 17292
rect 20901 17187 20959 17193
rect 20901 17153 20913 17187
rect 20947 17184 20959 17187
rect 22189 17187 22247 17193
rect 20947 17156 21956 17184
rect 20947 17153 20959 17156
rect 20901 17147 20959 17153
rect 20625 17119 20683 17125
rect 20625 17085 20637 17119
rect 20671 17116 20683 17119
rect 21818 17116 21824 17128
rect 20671 17088 21824 17116
rect 20671 17085 20683 17088
rect 20625 17079 20683 17085
rect 21818 17076 21824 17088
rect 21876 17076 21882 17128
rect 21928 17116 21956 17156
rect 22189 17153 22201 17187
rect 22235 17153 22247 17187
rect 22189 17147 22247 17153
rect 22370 17144 22376 17196
rect 22428 17144 22434 17196
rect 22465 17187 22523 17193
rect 22465 17153 22477 17187
rect 22511 17153 22523 17187
rect 22465 17147 22523 17153
rect 22278 17116 22284 17128
rect 21928 17088 22284 17116
rect 22278 17076 22284 17088
rect 22336 17076 22342 17128
rect 20717 17051 20775 17057
rect 20717 17017 20729 17051
rect 20763 17048 20775 17051
rect 21174 17048 21180 17060
rect 20763 17020 21180 17048
rect 20763 17017 20775 17020
rect 20717 17011 20775 17017
rect 21174 17008 21180 17020
rect 21232 17008 21238 17060
rect 21266 17008 21272 17060
rect 21324 17048 21330 17060
rect 22480 17048 22508 17147
rect 21324 17020 22508 17048
rect 21324 17008 21330 17020
rect 15068 16952 20116 16980
rect 20809 16983 20867 16989
rect 15068 16940 15074 16952
rect 20809 16949 20821 16983
rect 20855 16980 20867 16983
rect 22005 16983 22063 16989
rect 22005 16980 22017 16983
rect 20855 16952 22017 16980
rect 20855 16949 20867 16952
rect 20809 16943 20867 16949
rect 22005 16949 22017 16952
rect 22051 16949 22063 16983
rect 22005 16943 22063 16949
rect 1104 16890 23828 16912
rect 1104 16838 3790 16890
rect 3842 16838 3854 16890
rect 3906 16838 3918 16890
rect 3970 16838 3982 16890
rect 4034 16838 4046 16890
rect 4098 16838 9471 16890
rect 9523 16838 9535 16890
rect 9587 16838 9599 16890
rect 9651 16838 9663 16890
rect 9715 16838 9727 16890
rect 9779 16838 15152 16890
rect 15204 16838 15216 16890
rect 15268 16838 15280 16890
rect 15332 16838 15344 16890
rect 15396 16838 15408 16890
rect 15460 16838 20833 16890
rect 20885 16838 20897 16890
rect 20949 16838 20961 16890
rect 21013 16838 21025 16890
rect 21077 16838 21089 16890
rect 21141 16838 23828 16890
rect 1104 16816 23828 16838
rect 3436 16748 5396 16776
rect 3436 16581 3464 16748
rect 5368 16649 5396 16748
rect 8018 16736 8024 16788
rect 8076 16776 8082 16788
rect 13078 16776 13084 16788
rect 8076 16748 13084 16776
rect 8076 16736 8082 16748
rect 13078 16736 13084 16748
rect 13136 16736 13142 16788
rect 22097 16779 22155 16785
rect 22097 16776 22109 16779
rect 17420 16748 22109 16776
rect 11330 16668 11336 16720
rect 11388 16668 11394 16720
rect 14366 16708 14372 16720
rect 12636 16680 14372 16708
rect 5353 16643 5411 16649
rect 5353 16609 5365 16643
rect 5399 16609 5411 16643
rect 5353 16603 5411 16609
rect 6546 16600 6552 16652
rect 6604 16640 6610 16652
rect 8297 16643 8355 16649
rect 8297 16640 8309 16643
rect 6604 16612 8309 16640
rect 6604 16600 6610 16612
rect 8297 16609 8309 16612
rect 8343 16640 8355 16643
rect 8478 16640 8484 16652
rect 8343 16612 8484 16640
rect 8343 16609 8355 16612
rect 8297 16603 8355 16609
rect 8478 16600 8484 16612
rect 8536 16640 8542 16652
rect 9122 16640 9128 16652
rect 8536 16612 9128 16640
rect 8536 16600 8542 16612
rect 9122 16600 9128 16612
rect 9180 16600 9186 16652
rect 9401 16643 9459 16649
rect 9401 16609 9413 16643
rect 9447 16640 9459 16643
rect 11348 16640 11376 16668
rect 9447 16612 11376 16640
rect 9447 16609 9459 16612
rect 9401 16603 9459 16609
rect 12526 16600 12532 16652
rect 12584 16600 12590 16652
rect 12636 16649 12664 16680
rect 14366 16668 14372 16680
rect 14424 16668 14430 16720
rect 15933 16711 15991 16717
rect 15933 16708 15945 16711
rect 15396 16680 15945 16708
rect 12621 16643 12679 16649
rect 12621 16609 12633 16643
rect 12667 16609 12679 16643
rect 12621 16603 12679 16609
rect 12713 16643 12771 16649
rect 12713 16609 12725 16643
rect 12759 16609 12771 16643
rect 12713 16603 12771 16609
rect 3421 16575 3479 16581
rect 3421 16572 3433 16575
rect 3068 16544 3433 16572
rect 3068 16516 3096 16544
rect 3421 16541 3433 16544
rect 3467 16541 3479 16575
rect 3421 16535 3479 16541
rect 5097 16575 5155 16581
rect 5097 16541 5109 16575
rect 5143 16572 5155 16575
rect 7742 16572 7748 16584
rect 5143 16544 7748 16572
rect 5143 16541 5155 16544
rect 5097 16535 5155 16541
rect 7742 16532 7748 16544
rect 7800 16532 7806 16584
rect 8018 16532 8024 16584
rect 8076 16532 8082 16584
rect 12728 16572 12756 16603
rect 12802 16600 12808 16652
rect 12860 16600 12866 16652
rect 12894 16600 12900 16652
rect 12952 16640 12958 16652
rect 13262 16640 13268 16652
rect 12952 16612 13268 16640
rect 12952 16600 12958 16612
rect 13262 16600 13268 16612
rect 13320 16640 13326 16652
rect 13357 16643 13415 16649
rect 13357 16640 13369 16643
rect 13320 16612 13369 16640
rect 13320 16600 13326 16612
rect 13357 16609 13369 16612
rect 13403 16640 13415 16643
rect 15396 16640 15424 16680
rect 15933 16677 15945 16680
rect 15979 16677 15991 16711
rect 15933 16671 15991 16677
rect 13403 16612 13768 16640
rect 13403 16609 13415 16612
rect 13357 16603 13415 16609
rect 12912 16572 12940 16600
rect 12728 16544 12940 16572
rect 13740 16572 13768 16612
rect 14936 16612 15424 16640
rect 14936 16572 14964 16612
rect 16758 16600 16764 16652
rect 16816 16640 16822 16652
rect 17129 16643 17187 16649
rect 17129 16640 17141 16643
rect 16816 16612 17141 16640
rect 16816 16600 16822 16612
rect 17129 16609 17141 16612
rect 17175 16609 17187 16643
rect 17129 16603 17187 16609
rect 17221 16643 17279 16649
rect 17221 16609 17233 16643
rect 17267 16640 17279 16643
rect 17310 16640 17316 16652
rect 17267 16612 17316 16640
rect 17267 16609 17279 16612
rect 17221 16603 17279 16609
rect 17310 16600 17316 16612
rect 17368 16600 17374 16652
rect 13740 16544 14964 16572
rect 16482 16532 16488 16584
rect 16540 16572 16546 16584
rect 16850 16572 16856 16584
rect 16540 16544 16856 16572
rect 16540 16532 16546 16544
rect 16850 16532 16856 16544
rect 16908 16572 16914 16584
rect 17420 16581 17448 16748
rect 22097 16745 22109 16748
rect 22143 16745 22155 16779
rect 22097 16739 22155 16745
rect 22278 16736 22284 16788
rect 22336 16736 22342 16788
rect 17954 16668 17960 16720
rect 18012 16708 18018 16720
rect 18877 16711 18935 16717
rect 18877 16708 18889 16711
rect 18012 16680 18889 16708
rect 18012 16668 18018 16680
rect 18877 16677 18889 16680
rect 18923 16708 18935 16711
rect 19705 16711 19763 16717
rect 18923 16680 19656 16708
rect 18923 16677 18935 16680
rect 18877 16671 18935 16677
rect 17770 16600 17776 16652
rect 17828 16640 17834 16652
rect 18782 16640 18788 16652
rect 17828 16612 18788 16640
rect 17828 16600 17834 16612
rect 18782 16600 18788 16612
rect 18840 16640 18846 16652
rect 19628 16640 19656 16680
rect 19705 16677 19717 16711
rect 19751 16708 19763 16711
rect 20346 16708 20352 16720
rect 19751 16680 20352 16708
rect 19751 16677 19763 16680
rect 19705 16671 19763 16677
rect 20346 16668 20352 16680
rect 20404 16708 20410 16720
rect 20625 16711 20683 16717
rect 20625 16708 20637 16711
rect 20404 16680 20637 16708
rect 20404 16668 20410 16680
rect 20625 16677 20637 16680
rect 20671 16677 20683 16711
rect 20625 16671 20683 16677
rect 19889 16643 19947 16649
rect 19889 16640 19901 16643
rect 18840 16612 19564 16640
rect 19628 16612 19901 16640
rect 18840 16600 18846 16612
rect 17405 16575 17463 16581
rect 17405 16572 17417 16575
rect 16908 16544 17417 16572
rect 16908 16532 16914 16544
rect 17405 16541 17417 16544
rect 17451 16541 17463 16575
rect 17405 16535 17463 16541
rect 17494 16532 17500 16584
rect 17552 16532 17558 16584
rect 18141 16575 18199 16581
rect 18141 16541 18153 16575
rect 18187 16572 18199 16575
rect 18598 16572 18604 16584
rect 18187 16544 18604 16572
rect 18187 16541 18199 16544
rect 18141 16535 18199 16541
rect 18598 16532 18604 16544
rect 18656 16532 18662 16584
rect 19536 16572 19564 16612
rect 19889 16609 19901 16612
rect 19935 16640 19947 16643
rect 21174 16640 21180 16652
rect 19935 16612 21180 16640
rect 19935 16609 19947 16612
rect 19889 16603 19947 16609
rect 21174 16600 21180 16612
rect 21232 16600 21238 16652
rect 19613 16575 19671 16581
rect 19613 16572 19625 16575
rect 19536 16544 19625 16572
rect 19613 16541 19625 16544
rect 19659 16541 19671 16575
rect 19613 16535 19671 16541
rect 19797 16575 19855 16581
rect 19797 16541 19809 16575
rect 19843 16541 19855 16575
rect 19797 16535 19855 16541
rect 20073 16541 20131 16547
rect 3050 16464 3056 16516
rect 3108 16464 3114 16516
rect 3176 16507 3234 16513
rect 3176 16473 3188 16507
rect 3222 16504 3234 16507
rect 3602 16504 3608 16516
rect 3222 16476 3608 16504
rect 3222 16473 3234 16476
rect 3176 16467 3234 16473
rect 3602 16464 3608 16476
rect 3660 16464 3666 16516
rect 6270 16464 6276 16516
rect 6328 16504 6334 16516
rect 6641 16507 6699 16513
rect 6641 16504 6653 16507
rect 6328 16476 6653 16504
rect 6328 16464 6334 16476
rect 6641 16473 6653 16476
rect 6687 16473 6699 16507
rect 6641 16467 6699 16473
rect 10781 16507 10839 16513
rect 10781 16473 10793 16507
rect 10827 16504 10839 16507
rect 11698 16504 11704 16516
rect 10827 16476 11704 16504
rect 10827 16473 10839 16476
rect 10781 16467 10839 16473
rect 11698 16464 11704 16476
rect 11756 16464 11762 16516
rect 13998 16504 14004 16516
rect 12084 16476 14004 16504
rect 1486 16396 1492 16448
rect 1544 16436 1550 16448
rect 2041 16439 2099 16445
rect 2041 16436 2053 16439
rect 1544 16408 2053 16436
rect 1544 16396 1550 16408
rect 2041 16405 2053 16408
rect 2087 16405 2099 16439
rect 2041 16399 2099 16405
rect 3418 16396 3424 16448
rect 3476 16436 3482 16448
rect 3973 16439 4031 16445
rect 3973 16436 3985 16439
rect 3476 16408 3985 16436
rect 3476 16396 3482 16408
rect 3973 16405 3985 16408
rect 4019 16405 4031 16439
rect 3973 16399 4031 16405
rect 11422 16396 11428 16448
rect 11480 16436 11486 16448
rect 12084 16436 12112 16476
rect 13998 16464 14004 16476
rect 14056 16504 14062 16516
rect 14829 16507 14887 16513
rect 14829 16504 14841 16507
rect 14056 16476 14841 16504
rect 14056 16464 14062 16476
rect 14829 16473 14841 16476
rect 14875 16473 14887 16507
rect 14829 16467 14887 16473
rect 14918 16464 14924 16516
rect 14976 16504 14982 16516
rect 15473 16507 15531 16513
rect 15473 16504 15485 16507
rect 14976 16476 15485 16504
rect 14976 16464 14982 16476
rect 15473 16473 15485 16476
rect 15519 16504 15531 16507
rect 15838 16504 15844 16516
rect 15519 16476 15844 16504
rect 15519 16473 15531 16476
rect 15473 16467 15531 16473
rect 15838 16464 15844 16476
rect 15896 16504 15902 16516
rect 16942 16504 16948 16516
rect 15896 16476 16948 16504
rect 15896 16464 15902 16476
rect 16942 16464 16948 16476
rect 17000 16464 17006 16516
rect 17034 16464 17040 16516
rect 17092 16464 17098 16516
rect 18690 16464 18696 16516
rect 18748 16504 18754 16516
rect 19812 16504 19840 16535
rect 18748 16476 19840 16504
rect 18748 16464 18754 16476
rect 11480 16408 12112 16436
rect 11480 16396 11486 16408
rect 12158 16396 12164 16448
rect 12216 16436 12222 16448
rect 12345 16439 12403 16445
rect 12345 16436 12357 16439
rect 12216 16408 12357 16436
rect 12216 16396 12222 16408
rect 12345 16405 12357 16408
rect 12391 16405 12403 16439
rect 12345 16399 12403 16405
rect 14369 16439 14427 16445
rect 14369 16405 14381 16439
rect 14415 16436 14427 16439
rect 15378 16436 15384 16448
rect 14415 16408 15384 16436
rect 14415 16405 14427 16408
rect 14369 16399 14427 16405
rect 15378 16396 15384 16408
rect 15436 16396 15442 16448
rect 17770 16396 17776 16448
rect 17828 16436 17834 16448
rect 18049 16439 18107 16445
rect 18049 16436 18061 16439
rect 17828 16408 18061 16436
rect 17828 16396 17834 16408
rect 18049 16405 18061 16408
rect 18095 16405 18107 16439
rect 18049 16399 18107 16405
rect 19429 16439 19487 16445
rect 19429 16405 19441 16439
rect 19475 16436 19487 16439
rect 19518 16436 19524 16448
rect 19475 16408 19524 16436
rect 19475 16405 19487 16408
rect 19429 16399 19487 16405
rect 19518 16396 19524 16408
rect 19576 16396 19582 16448
rect 19812 16436 19840 16476
rect 19886 16464 19892 16516
rect 19944 16504 19950 16516
rect 20073 16507 20085 16541
rect 20119 16507 20131 16541
rect 20073 16504 20131 16507
rect 21913 16507 21971 16513
rect 21913 16504 21925 16507
rect 19944 16501 20131 16504
rect 19944 16476 20116 16501
rect 20180 16476 21925 16504
rect 19944 16464 19950 16476
rect 20180 16436 20208 16476
rect 21913 16473 21925 16476
rect 21959 16473 21971 16507
rect 21913 16467 21971 16473
rect 19812 16408 20208 16436
rect 21450 16396 21456 16448
rect 21508 16436 21514 16448
rect 22113 16439 22171 16445
rect 22113 16436 22125 16439
rect 21508 16408 22125 16436
rect 21508 16396 21514 16408
rect 22113 16405 22125 16408
rect 22159 16405 22171 16439
rect 22113 16399 22171 16405
rect 1104 16346 23987 16368
rect 1104 16294 6630 16346
rect 6682 16294 6694 16346
rect 6746 16294 6758 16346
rect 6810 16294 6822 16346
rect 6874 16294 6886 16346
rect 6938 16294 12311 16346
rect 12363 16294 12375 16346
rect 12427 16294 12439 16346
rect 12491 16294 12503 16346
rect 12555 16294 12567 16346
rect 12619 16294 17992 16346
rect 18044 16294 18056 16346
rect 18108 16294 18120 16346
rect 18172 16294 18184 16346
rect 18236 16294 18248 16346
rect 18300 16294 23673 16346
rect 23725 16294 23737 16346
rect 23789 16294 23801 16346
rect 23853 16294 23865 16346
rect 23917 16294 23929 16346
rect 23981 16294 23987 16346
rect 1104 16272 23987 16294
rect 9122 16192 9128 16244
rect 9180 16192 9186 16244
rect 15381 16235 15439 16241
rect 15381 16201 15393 16235
rect 15427 16232 15439 16235
rect 15746 16232 15752 16244
rect 15427 16204 15752 16232
rect 15427 16201 15439 16204
rect 15381 16195 15439 16201
rect 15746 16192 15752 16204
rect 15804 16192 15810 16244
rect 18325 16235 18383 16241
rect 18325 16201 18337 16235
rect 18371 16232 18383 16235
rect 18690 16232 18696 16244
rect 18371 16204 18696 16232
rect 18371 16201 18383 16204
rect 18325 16195 18383 16201
rect 4338 16124 4344 16176
rect 4396 16124 4402 16176
rect 7650 16124 7656 16176
rect 7708 16164 7714 16176
rect 7837 16167 7895 16173
rect 7837 16164 7849 16167
rect 7708 16136 7849 16164
rect 7708 16124 7714 16136
rect 7837 16133 7849 16136
rect 7883 16133 7895 16167
rect 7837 16127 7895 16133
rect 11698 16124 11704 16176
rect 11756 16164 11762 16176
rect 18340 16164 18368 16195
rect 18690 16192 18696 16204
rect 18748 16192 18754 16244
rect 20438 16232 20444 16244
rect 20180 16204 20444 16232
rect 20180 16164 20208 16204
rect 20438 16192 20444 16204
rect 20496 16192 20502 16244
rect 20714 16192 20720 16244
rect 20772 16192 20778 16244
rect 22370 16192 22376 16244
rect 22428 16192 22434 16244
rect 11756 16136 12434 16164
rect 11756 16124 11762 16136
rect 12158 16056 12164 16108
rect 12216 16096 12222 16108
rect 12253 16099 12311 16105
rect 12253 16096 12265 16099
rect 12216 16068 12265 16096
rect 12216 16056 12222 16068
rect 12253 16065 12265 16068
rect 12299 16065 12311 16099
rect 12406 16096 12434 16136
rect 17328 16136 18368 16164
rect 19306 16136 20208 16164
rect 12621 16099 12679 16105
rect 12621 16096 12633 16099
rect 12406 16068 12633 16096
rect 12253 16059 12311 16065
rect 12621 16065 12633 16068
rect 12667 16065 12679 16099
rect 12621 16059 12679 16065
rect 15562 16056 15568 16108
rect 15620 16056 15626 16108
rect 15654 16056 15660 16108
rect 15712 16056 15718 16108
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16096 15991 16099
rect 16390 16096 16396 16108
rect 15979 16068 16396 16096
rect 15979 16065 15991 16068
rect 15933 16059 15991 16065
rect 16390 16056 16396 16068
rect 16448 16056 16454 16108
rect 17034 16056 17040 16108
rect 17092 16096 17098 16108
rect 17218 16096 17224 16108
rect 17092 16068 17224 16096
rect 17092 16056 17098 16068
rect 17218 16056 17224 16068
rect 17276 16056 17282 16108
rect 17328 16105 17356 16136
rect 17313 16099 17371 16105
rect 17313 16065 17325 16099
rect 17359 16065 17371 16099
rect 17313 16059 17371 16065
rect 17586 16056 17592 16108
rect 17644 16056 17650 16108
rect 18509 16099 18567 16105
rect 18509 16065 18521 16099
rect 18555 16096 18567 16099
rect 18966 16096 18972 16108
rect 18555 16068 18972 16096
rect 18555 16065 18567 16068
rect 18509 16059 18567 16065
rect 18966 16056 18972 16068
rect 19024 16056 19030 16108
rect 13630 15988 13636 16040
rect 13688 16028 13694 16040
rect 14553 16031 14611 16037
rect 14553 16028 14565 16031
rect 13688 16000 14565 16028
rect 13688 15988 13694 16000
rect 14553 15997 14565 16000
rect 14599 16028 14611 16031
rect 15010 16028 15016 16040
rect 14599 16000 15016 16028
rect 14599 15997 14611 16000
rect 14553 15991 14611 15997
rect 15010 15988 15016 16000
rect 15068 15988 15074 16040
rect 19058 15988 19064 16040
rect 19116 16028 19122 16040
rect 19306 16028 19334 16136
rect 20180 16105 20208 16136
rect 20165 16099 20223 16105
rect 20165 16065 20177 16099
rect 20211 16065 20223 16099
rect 20165 16059 20223 16065
rect 20254 16056 20260 16108
rect 20312 16056 20318 16108
rect 20441 16099 20499 16105
rect 20441 16065 20453 16099
rect 20487 16065 20499 16099
rect 20441 16059 20499 16065
rect 20533 16099 20591 16105
rect 20533 16065 20545 16099
rect 20579 16096 20591 16099
rect 20622 16096 20628 16108
rect 20579 16068 20628 16096
rect 20579 16065 20591 16068
rect 20533 16059 20591 16065
rect 19116 16000 19334 16028
rect 20456 16028 20484 16059
rect 20622 16056 20628 16068
rect 20680 16056 20686 16108
rect 22097 16099 22155 16105
rect 22097 16065 22109 16099
rect 22143 16096 22155 16099
rect 22922 16096 22928 16108
rect 22143 16068 22928 16096
rect 22143 16065 22155 16068
rect 22097 16059 22155 16065
rect 22922 16056 22928 16068
rect 22980 16056 22986 16108
rect 20456 16000 20576 16028
rect 19116 15988 19122 16000
rect 12618 15920 12624 15972
rect 12676 15960 12682 15972
rect 13648 15960 13676 15988
rect 12676 15932 13676 15960
rect 12676 15920 12682 15932
rect 19150 15920 19156 15972
rect 19208 15960 19214 15972
rect 19886 15960 19892 15972
rect 19208 15932 19892 15960
rect 19208 15920 19214 15932
rect 19886 15920 19892 15932
rect 19944 15920 19950 15972
rect 20548 15904 20576 16000
rect 3050 15852 3056 15904
rect 3108 15852 3114 15904
rect 11238 15852 11244 15904
rect 11296 15892 11302 15904
rect 12342 15892 12348 15904
rect 11296 15864 12348 15892
rect 11296 15852 11302 15864
rect 12342 15852 12348 15864
rect 12400 15852 12406 15904
rect 13906 15852 13912 15904
rect 13964 15852 13970 15904
rect 15841 15895 15899 15901
rect 15841 15861 15853 15895
rect 15887 15892 15899 15895
rect 17034 15892 17040 15904
rect 15887 15864 17040 15892
rect 15887 15861 15899 15864
rect 15841 15855 15899 15861
rect 17034 15852 17040 15864
rect 17092 15852 17098 15904
rect 17310 15852 17316 15904
rect 17368 15892 17374 15904
rect 17405 15895 17463 15901
rect 17405 15892 17417 15895
rect 17368 15864 17417 15892
rect 17368 15852 17374 15864
rect 17405 15861 17417 15864
rect 17451 15861 17463 15895
rect 17405 15855 17463 15861
rect 17678 15852 17684 15904
rect 17736 15892 17742 15904
rect 17773 15895 17831 15901
rect 17773 15892 17785 15895
rect 17736 15864 17785 15892
rect 17736 15852 17742 15864
rect 17773 15861 17785 15864
rect 17819 15861 17831 15895
rect 17773 15855 17831 15861
rect 19705 15895 19763 15901
rect 19705 15861 19717 15895
rect 19751 15892 19763 15895
rect 20530 15892 20536 15904
rect 19751 15864 20536 15892
rect 19751 15861 19763 15864
rect 19705 15855 19763 15861
rect 20530 15852 20536 15864
rect 20588 15852 20594 15904
rect 20714 15852 20720 15904
rect 20772 15892 20778 15904
rect 22370 15892 22376 15904
rect 20772 15864 22376 15892
rect 20772 15852 20778 15864
rect 22370 15852 22376 15864
rect 22428 15852 22434 15904
rect 1104 15802 23828 15824
rect 1104 15750 3790 15802
rect 3842 15750 3854 15802
rect 3906 15750 3918 15802
rect 3970 15750 3982 15802
rect 4034 15750 4046 15802
rect 4098 15750 9471 15802
rect 9523 15750 9535 15802
rect 9587 15750 9599 15802
rect 9651 15750 9663 15802
rect 9715 15750 9727 15802
rect 9779 15750 15152 15802
rect 15204 15750 15216 15802
rect 15268 15750 15280 15802
rect 15332 15750 15344 15802
rect 15396 15750 15408 15802
rect 15460 15750 20833 15802
rect 20885 15750 20897 15802
rect 20949 15750 20961 15802
rect 21013 15750 21025 15802
rect 21077 15750 21089 15802
rect 21141 15750 23828 15802
rect 1104 15728 23828 15750
rect 12066 15648 12072 15700
rect 12124 15688 12130 15700
rect 13173 15691 13231 15697
rect 13173 15688 13185 15691
rect 12124 15660 13185 15688
rect 12124 15648 12130 15660
rect 13173 15657 13185 15660
rect 13219 15657 13231 15691
rect 13173 15651 13231 15657
rect 13446 15648 13452 15700
rect 13504 15688 13510 15700
rect 13504 15660 15700 15688
rect 13504 15648 13510 15660
rect 10594 15580 10600 15632
rect 10652 15620 10658 15632
rect 14461 15623 14519 15629
rect 14461 15620 14473 15623
rect 10652 15592 14473 15620
rect 10652 15580 10658 15592
rect 14461 15589 14473 15592
rect 14507 15589 14519 15623
rect 14461 15583 14519 15589
rect 6546 15512 6552 15564
rect 6604 15552 6610 15564
rect 6733 15555 6791 15561
rect 6733 15552 6745 15555
rect 6604 15524 6745 15552
rect 6604 15512 6610 15524
rect 6733 15521 6745 15524
rect 6779 15521 6791 15555
rect 6733 15515 6791 15521
rect 9122 15512 9128 15564
rect 9180 15512 9186 15564
rect 12158 15512 12164 15564
rect 12216 15552 12222 15564
rect 12345 15555 12403 15561
rect 12345 15552 12357 15555
rect 12216 15524 12357 15552
rect 12216 15512 12222 15524
rect 12345 15521 12357 15524
rect 12391 15521 12403 15555
rect 12345 15515 12403 15521
rect 12434 15512 12440 15564
rect 12492 15552 12498 15564
rect 13541 15555 13599 15561
rect 12492 15524 12572 15552
rect 12492 15512 12498 15524
rect 2406 15444 2412 15496
rect 2464 15444 2470 15496
rect 4522 15444 4528 15496
rect 4580 15484 4586 15496
rect 4982 15484 4988 15496
rect 4580 15456 4988 15484
rect 4580 15444 4586 15456
rect 4982 15444 4988 15456
rect 5040 15484 5046 15496
rect 5629 15487 5687 15493
rect 5629 15484 5641 15487
rect 5040 15456 5641 15484
rect 5040 15444 5046 15456
rect 5629 15453 5641 15456
rect 5675 15484 5687 15487
rect 8294 15484 8300 15496
rect 5675 15456 8300 15484
rect 5675 15453 5687 15456
rect 5629 15447 5687 15453
rect 8294 15444 8300 15456
rect 8352 15444 8358 15496
rect 9392 15487 9450 15493
rect 9392 15453 9404 15487
rect 9438 15484 9450 15487
rect 9438 15456 11192 15484
rect 9438 15453 9450 15456
rect 9392 15447 9450 15453
rect 5166 15376 5172 15428
rect 5224 15416 5230 15428
rect 5261 15419 5319 15425
rect 5261 15416 5273 15419
rect 5224 15388 5273 15416
rect 5224 15376 5230 15388
rect 5261 15385 5273 15388
rect 5307 15385 5319 15419
rect 5261 15379 5319 15385
rect 7000 15419 7058 15425
rect 7000 15385 7012 15419
rect 7046 15416 7058 15419
rect 11054 15416 11060 15428
rect 7046 15388 11060 15416
rect 7046 15385 7058 15388
rect 7000 15379 7058 15385
rect 11054 15376 11060 15388
rect 11112 15376 11118 15428
rect 2225 15351 2283 15357
rect 2225 15317 2237 15351
rect 2271 15348 2283 15351
rect 2498 15348 2504 15360
rect 2271 15320 2504 15348
rect 2271 15317 2283 15320
rect 2225 15311 2283 15317
rect 2498 15308 2504 15320
rect 2556 15308 2562 15360
rect 8113 15351 8171 15357
rect 8113 15317 8125 15351
rect 8159 15348 8171 15351
rect 10134 15348 10140 15360
rect 8159 15320 10140 15348
rect 8159 15317 8171 15320
rect 8113 15311 8171 15317
rect 10134 15308 10140 15320
rect 10192 15308 10198 15360
rect 10410 15308 10416 15360
rect 10468 15348 10474 15360
rect 11164 15357 11192 15456
rect 11330 15444 11336 15496
rect 11388 15484 11394 15496
rect 11698 15484 11704 15496
rect 11388 15456 11704 15484
rect 11388 15444 11394 15456
rect 11698 15444 11704 15456
rect 11756 15484 11762 15496
rect 12544 15493 12572 15524
rect 13541 15521 13553 15555
rect 13587 15552 13599 15555
rect 13587 15524 13768 15552
rect 13587 15521 13599 15524
rect 13541 15515 13599 15521
rect 12253 15487 12311 15493
rect 12253 15484 12265 15487
rect 11756 15456 12265 15484
rect 11756 15444 11762 15456
rect 12253 15453 12265 15456
rect 12299 15453 12311 15487
rect 12253 15447 12311 15453
rect 12529 15487 12587 15493
rect 12529 15453 12541 15487
rect 12575 15453 12587 15487
rect 12529 15447 12587 15453
rect 13354 15444 13360 15496
rect 13412 15444 13418 15496
rect 13449 15487 13507 15493
rect 13449 15453 13461 15487
rect 13495 15453 13507 15487
rect 13449 15447 13507 15453
rect 11793 15419 11851 15425
rect 11793 15385 11805 15419
rect 11839 15416 11851 15419
rect 12618 15416 12624 15428
rect 11839 15388 12624 15416
rect 11839 15385 11851 15388
rect 11793 15379 11851 15385
rect 12618 15376 12624 15388
rect 12676 15376 12682 15428
rect 13464 15416 13492 15447
rect 13630 15444 13636 15496
rect 13688 15444 13694 15496
rect 13740 15484 13768 15524
rect 15010 15512 15016 15564
rect 15068 15512 15074 15564
rect 14274 15484 14280 15496
rect 13740 15456 14280 15484
rect 14274 15444 14280 15456
rect 14332 15444 14338 15496
rect 15470 15484 15476 15496
rect 14384 15456 15476 15484
rect 14384 15416 14412 15456
rect 15470 15444 15476 15456
rect 15528 15444 15534 15496
rect 15672 15493 15700 15660
rect 17034 15648 17040 15700
rect 17092 15648 17098 15700
rect 18877 15691 18935 15697
rect 18877 15657 18889 15691
rect 18923 15688 18935 15691
rect 18923 15660 19932 15688
rect 18923 15657 18935 15660
rect 18877 15651 18935 15657
rect 17494 15580 17500 15632
rect 17552 15620 17558 15632
rect 17552 15592 19380 15620
rect 17552 15580 17558 15592
rect 15933 15555 15991 15561
rect 15933 15521 15945 15555
rect 15979 15552 15991 15555
rect 16390 15552 16396 15564
rect 15979 15524 16396 15552
rect 15979 15521 15991 15524
rect 15933 15515 15991 15521
rect 15657 15487 15715 15493
rect 15657 15453 15669 15487
rect 15703 15453 15715 15487
rect 15657 15447 15715 15453
rect 13464 15388 14412 15416
rect 14829 15419 14887 15425
rect 14829 15385 14841 15419
rect 14875 15416 14887 15419
rect 15838 15416 15844 15428
rect 14875 15388 15844 15416
rect 14875 15385 14887 15388
rect 14829 15379 14887 15385
rect 15838 15376 15844 15388
rect 15896 15376 15902 15428
rect 10505 15351 10563 15357
rect 10505 15348 10517 15351
rect 10468 15320 10517 15348
rect 10468 15308 10474 15320
rect 10505 15317 10517 15320
rect 10551 15317 10563 15351
rect 10505 15311 10563 15317
rect 11149 15351 11207 15357
rect 11149 15317 11161 15351
rect 11195 15348 11207 15351
rect 11422 15348 11428 15360
rect 11195 15320 11428 15348
rect 11195 15317 11207 15320
rect 11149 15311 11207 15317
rect 11422 15308 11428 15320
rect 11480 15308 11486 15360
rect 12710 15308 12716 15360
rect 12768 15308 12774 15360
rect 14918 15308 14924 15360
rect 14976 15308 14982 15360
rect 15194 15308 15200 15360
rect 15252 15348 15258 15360
rect 15948 15348 15976 15515
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 17678 15512 17684 15564
rect 17736 15512 17742 15564
rect 18785 15555 18843 15561
rect 18785 15521 18797 15555
rect 18831 15552 18843 15555
rect 19242 15552 19248 15564
rect 18831 15524 19248 15552
rect 18831 15521 18843 15524
rect 18785 15515 18843 15521
rect 19242 15512 19248 15524
rect 19300 15512 19306 15564
rect 19352 15552 19380 15592
rect 19426 15580 19432 15632
rect 19484 15580 19490 15632
rect 19904 15552 19932 15660
rect 21818 15648 21824 15700
rect 21876 15648 21882 15700
rect 22646 15552 22652 15564
rect 19352 15524 19748 15552
rect 17221 15487 17279 15493
rect 17221 15453 17233 15487
rect 17267 15484 17279 15487
rect 17770 15484 17776 15496
rect 17267 15456 17776 15484
rect 17267 15453 17279 15456
rect 17221 15447 17279 15453
rect 17770 15444 17776 15456
rect 17828 15444 17834 15496
rect 19720 15493 19748 15524
rect 19904 15524 22652 15552
rect 19904 15493 19932 15524
rect 22646 15512 22652 15524
rect 22704 15512 22710 15564
rect 18877 15487 18935 15493
rect 18877 15453 18889 15487
rect 18923 15484 18935 15487
rect 19613 15487 19671 15493
rect 19613 15484 19625 15487
rect 18923 15456 19625 15484
rect 18923 15453 18935 15456
rect 18877 15447 18935 15453
rect 19613 15453 19625 15456
rect 19659 15453 19671 15487
rect 19613 15447 19671 15453
rect 19705 15487 19763 15493
rect 19705 15453 19717 15487
rect 19751 15453 19763 15487
rect 19705 15447 19763 15453
rect 19889 15487 19947 15493
rect 19889 15453 19901 15487
rect 19935 15453 19947 15487
rect 19889 15447 19947 15453
rect 19981 15487 20039 15493
rect 19981 15453 19993 15487
rect 20027 15484 20039 15487
rect 20162 15484 20168 15496
rect 20027 15456 20168 15484
rect 20027 15453 20039 15456
rect 19981 15447 20039 15453
rect 16850 15376 16856 15428
rect 16908 15416 16914 15428
rect 17313 15419 17371 15425
rect 17313 15416 17325 15419
rect 16908 15388 17325 15416
rect 16908 15376 16914 15388
rect 17313 15385 17325 15388
rect 17359 15385 17371 15419
rect 17313 15379 17371 15385
rect 17405 15419 17463 15425
rect 17405 15385 17417 15419
rect 17451 15385 17463 15419
rect 17405 15379 17463 15385
rect 17543 15419 17601 15425
rect 17543 15385 17555 15419
rect 17589 15416 17601 15419
rect 17589 15388 18552 15416
rect 17589 15385 17601 15388
rect 17543 15379 17601 15385
rect 15252 15320 15976 15348
rect 15252 15308 15258 15320
rect 16666 15308 16672 15360
rect 16724 15348 16730 15360
rect 17420 15348 17448 15379
rect 18524 15357 18552 15388
rect 16724 15320 17448 15348
rect 18509 15351 18567 15357
rect 16724 15308 16730 15320
rect 18509 15317 18521 15351
rect 18555 15317 18567 15351
rect 19628 15348 19656 15447
rect 19720 15416 19748 15447
rect 20162 15444 20168 15456
rect 20220 15484 20226 15496
rect 21361 15487 21419 15493
rect 21361 15484 21373 15487
rect 20220 15456 21373 15484
rect 20220 15444 20226 15456
rect 21361 15453 21373 15456
rect 21407 15484 21419 15487
rect 22005 15487 22063 15493
rect 22005 15484 22017 15487
rect 21407 15456 22017 15484
rect 21407 15453 21419 15456
rect 21361 15447 21419 15453
rect 22005 15453 22017 15456
rect 22051 15484 22063 15487
rect 22094 15484 22100 15496
rect 22051 15456 22100 15484
rect 22051 15453 22063 15456
rect 22005 15447 22063 15453
rect 22094 15444 22100 15456
rect 22152 15444 22158 15496
rect 22278 15444 22284 15496
rect 22336 15444 22342 15496
rect 20714 15416 20720 15428
rect 19720 15388 20720 15416
rect 20714 15376 20720 15388
rect 20772 15376 20778 15428
rect 21085 15419 21143 15425
rect 21085 15385 21097 15419
rect 21131 15416 21143 15419
rect 21634 15416 21640 15428
rect 21131 15388 21640 15416
rect 21131 15385 21143 15388
rect 21085 15379 21143 15385
rect 21634 15376 21640 15388
rect 21692 15376 21698 15428
rect 21266 15348 21272 15360
rect 19628 15320 21272 15348
rect 18509 15311 18567 15317
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 22189 15351 22247 15357
rect 22189 15317 22201 15351
rect 22235 15348 22247 15351
rect 22462 15348 22468 15360
rect 22235 15320 22468 15348
rect 22235 15317 22247 15320
rect 22189 15311 22247 15317
rect 22462 15308 22468 15320
rect 22520 15308 22526 15360
rect 1104 15258 23987 15280
rect 1104 15206 6630 15258
rect 6682 15206 6694 15258
rect 6746 15206 6758 15258
rect 6810 15206 6822 15258
rect 6874 15206 6886 15258
rect 6938 15206 12311 15258
rect 12363 15206 12375 15258
rect 12427 15206 12439 15258
rect 12491 15206 12503 15258
rect 12555 15206 12567 15258
rect 12619 15206 17992 15258
rect 18044 15206 18056 15258
rect 18108 15206 18120 15258
rect 18172 15206 18184 15258
rect 18236 15206 18248 15258
rect 18300 15206 23673 15258
rect 23725 15206 23737 15258
rect 23789 15206 23801 15258
rect 23853 15206 23865 15258
rect 23917 15206 23929 15258
rect 23981 15206 23987 15258
rect 1104 15184 23987 15206
rect 2409 15147 2467 15153
rect 2409 15113 2421 15147
rect 2455 15144 2467 15147
rect 2958 15144 2964 15156
rect 2455 15116 2964 15144
rect 2455 15113 2467 15116
rect 2409 15107 2467 15113
rect 2958 15104 2964 15116
rect 3016 15104 3022 15156
rect 14829 15147 14887 15153
rect 12406 15116 14688 15144
rect 2133 15079 2191 15085
rect 2133 15045 2145 15079
rect 2179 15076 2191 15079
rect 2498 15076 2504 15088
rect 2179 15048 2504 15076
rect 2179 15045 2191 15048
rect 2133 15039 2191 15045
rect 2498 15036 2504 15048
rect 2556 15036 2562 15088
rect 5442 15036 5448 15088
rect 5500 15076 5506 15088
rect 5629 15079 5687 15085
rect 5629 15076 5641 15079
rect 5500 15048 5641 15076
rect 5500 15036 5506 15048
rect 5629 15045 5641 15048
rect 5675 15045 5687 15079
rect 5629 15039 5687 15045
rect 6733 15079 6791 15085
rect 6733 15045 6745 15079
rect 6779 15076 6791 15079
rect 7006 15076 7012 15088
rect 6779 15048 7012 15076
rect 6779 15045 6791 15048
rect 6733 15039 6791 15045
rect 7006 15036 7012 15048
rect 7064 15076 7070 15088
rect 7285 15079 7343 15085
rect 7285 15076 7297 15079
rect 7064 15048 7297 15076
rect 7064 15036 7070 15048
rect 7285 15045 7297 15048
rect 7331 15045 7343 15079
rect 7285 15039 7343 15045
rect 9392 15079 9450 15085
rect 9392 15045 9404 15079
rect 9438 15076 9450 15079
rect 12406 15076 12434 15116
rect 9438 15048 12434 15076
rect 9438 15045 9450 15048
rect 9392 15039 9450 15045
rect 13538 15036 13544 15088
rect 13596 15036 13602 15088
rect 14550 15036 14556 15088
rect 14608 15036 14614 15088
rect 14660 15076 14688 15116
rect 14829 15113 14841 15147
rect 14875 15144 14887 15147
rect 14918 15144 14924 15156
rect 14875 15116 14924 15144
rect 14875 15113 14887 15116
rect 14829 15107 14887 15113
rect 14918 15104 14924 15116
rect 14976 15104 14982 15156
rect 15838 15104 15844 15156
rect 15896 15144 15902 15156
rect 16853 15147 16911 15153
rect 16853 15144 16865 15147
rect 15896 15116 16865 15144
rect 15896 15104 15902 15116
rect 16853 15113 16865 15116
rect 16899 15113 16911 15147
rect 16853 15107 16911 15113
rect 17310 15104 17316 15156
rect 17368 15144 17374 15156
rect 17494 15144 17500 15156
rect 17368 15116 17500 15144
rect 17368 15104 17374 15116
rect 17494 15104 17500 15116
rect 17552 15104 17558 15156
rect 17678 15104 17684 15156
rect 17736 15144 17742 15156
rect 18782 15144 18788 15156
rect 17736 15116 18788 15144
rect 17736 15104 17742 15116
rect 18782 15104 18788 15116
rect 18840 15104 18846 15156
rect 19702 15144 19708 15156
rect 19168 15116 19708 15144
rect 17862 15076 17868 15088
rect 14660 15048 17868 15076
rect 17862 15036 17868 15048
rect 17920 15036 17926 15088
rect 19168 15076 19196 15116
rect 19702 15104 19708 15116
rect 19760 15104 19766 15156
rect 21174 15104 21180 15156
rect 21232 15144 21238 15156
rect 21232 15116 22094 15144
rect 21232 15104 21238 15116
rect 20438 15076 20444 15088
rect 18156 15048 19196 15076
rect 19260 15048 20444 15076
rect 1854 14968 1860 15020
rect 1912 14968 1918 15020
rect 2038 14968 2044 15020
rect 2096 14968 2102 15020
rect 2222 14968 2228 15020
rect 2280 14968 2286 15020
rect 5994 14968 6000 15020
rect 6052 15008 6058 15020
rect 6549 15011 6607 15017
rect 6549 15008 6561 15011
rect 6052 14980 6561 15008
rect 6052 14968 6058 14980
rect 6549 14977 6561 14980
rect 6595 14977 6607 15011
rect 6549 14971 6607 14977
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 15008 6883 15011
rect 7374 15008 7380 15020
rect 6871 14980 7380 15008
rect 6871 14977 6883 14980
rect 6825 14971 6883 14977
rect 7374 14968 7380 14980
rect 7432 14968 7438 15020
rect 9122 14968 9128 15020
rect 9180 14968 9186 15020
rect 11054 14968 11060 15020
rect 11112 15008 11118 15020
rect 11793 15011 11851 15017
rect 11793 15008 11805 15011
rect 11112 14980 11805 15008
rect 11112 14968 11118 14980
rect 11793 14977 11805 14980
rect 11839 14977 11851 15011
rect 11793 14971 11851 14977
rect 12894 14968 12900 15020
rect 12952 14968 12958 15020
rect 13265 15011 13323 15017
rect 13265 14977 13277 15011
rect 13311 15008 13323 15011
rect 14090 15008 14096 15020
rect 13311 14980 14096 15008
rect 13311 14977 13323 14980
rect 13265 14971 13323 14977
rect 14090 14968 14096 14980
rect 14148 14968 14154 15020
rect 14274 14968 14280 15020
rect 14332 14968 14338 15020
rect 14458 14968 14464 15020
rect 14516 14968 14522 15020
rect 14642 14968 14648 15020
rect 14700 14968 14706 15020
rect 15654 14968 15660 15020
rect 15712 15008 15718 15020
rect 15930 15008 15936 15020
rect 15712 14980 15936 15008
rect 15712 14968 15718 14980
rect 15930 14968 15936 14980
rect 15988 14968 15994 15020
rect 16022 14968 16028 15020
rect 16080 14968 16086 15020
rect 16209 15011 16267 15017
rect 16209 14977 16221 15011
rect 16255 14977 16267 15011
rect 16209 14971 16267 14977
rect 3050 14900 3056 14952
rect 3108 14900 3114 14952
rect 3329 14943 3387 14949
rect 3329 14909 3341 14943
rect 3375 14940 3387 14943
rect 6086 14940 6092 14952
rect 3375 14912 6092 14940
rect 3375 14909 3387 14912
rect 3329 14903 3387 14909
rect 6086 14900 6092 14912
rect 6144 14900 6150 14952
rect 12066 14900 12072 14952
rect 12124 14900 12130 14952
rect 12710 14900 12716 14952
rect 12768 14940 12774 14952
rect 13357 14943 13415 14949
rect 13357 14940 13369 14943
rect 12768 14912 13369 14940
rect 12768 14900 12774 14912
rect 13357 14909 13369 14912
rect 13403 14909 13415 14943
rect 14292 14940 14320 14968
rect 15194 14940 15200 14952
rect 14292 14912 15200 14940
rect 13357 14903 13415 14909
rect 15194 14900 15200 14912
rect 15252 14900 15258 14952
rect 16224 14940 16252 14971
rect 16298 14968 16304 15020
rect 16356 14968 16362 15020
rect 16666 14968 16672 15020
rect 16724 15008 16730 15020
rect 16724 14980 17172 15008
rect 16724 14968 16730 14980
rect 15948 14912 16252 14940
rect 15948 14884 15976 14912
rect 17034 14900 17040 14952
rect 17092 14900 17098 14952
rect 17144 14949 17172 14980
rect 17218 14968 17224 15020
rect 17276 14968 17282 15020
rect 17313 15011 17371 15017
rect 17313 14977 17325 15011
rect 17359 15008 17371 15011
rect 18156 15008 18184 15048
rect 17359 14980 18184 15008
rect 18233 15011 18291 15017
rect 17359 14977 17371 14980
rect 17313 14971 17371 14977
rect 18233 14977 18245 15011
rect 18279 14977 18291 15011
rect 18233 14971 18291 14977
rect 18417 15011 18475 15017
rect 18417 14977 18429 15011
rect 18463 15008 18475 15011
rect 18782 15008 18788 15020
rect 18463 14980 18788 15008
rect 18463 14977 18475 14980
rect 18417 14971 18475 14977
rect 17129 14943 17187 14949
rect 17129 14909 17141 14943
rect 17175 14940 17187 14943
rect 17770 14940 17776 14952
rect 17175 14912 17776 14940
rect 17175 14909 17187 14912
rect 17129 14903 17187 14909
rect 17770 14900 17776 14912
rect 17828 14900 17834 14952
rect 18248 14940 18276 14971
rect 18782 14968 18788 14980
rect 18840 14968 18846 15020
rect 19260 15017 19288 15048
rect 20438 15036 20444 15048
rect 20496 15036 20502 15088
rect 22066 15076 22094 15116
rect 22554 15104 22560 15156
rect 22612 15104 22618 15156
rect 22066 15048 22876 15076
rect 19245 15011 19303 15017
rect 19245 15008 19257 15011
rect 18892 14980 19257 15008
rect 18690 14940 18696 14952
rect 18248 14912 18696 14940
rect 18690 14900 18696 14912
rect 18748 14900 18754 14952
rect 4617 14875 4675 14881
rect 4617 14841 4629 14875
rect 4663 14872 4675 14875
rect 5902 14872 5908 14884
rect 4663 14844 5908 14872
rect 4663 14841 4675 14844
rect 4617 14835 4675 14841
rect 5902 14832 5908 14844
rect 5960 14872 5966 14884
rect 6638 14872 6644 14884
rect 5960 14844 6644 14872
rect 5960 14832 5966 14844
rect 6638 14832 6644 14844
rect 6696 14832 6702 14884
rect 14550 14832 14556 14884
rect 14608 14872 14614 14884
rect 14608 14844 15884 14872
rect 14608 14832 14614 14844
rect 5350 14764 5356 14816
rect 5408 14804 5414 14816
rect 5721 14807 5779 14813
rect 5721 14804 5733 14807
rect 5408 14776 5733 14804
rect 5408 14764 5414 14776
rect 5721 14773 5733 14776
rect 5767 14773 5779 14807
rect 5721 14767 5779 14773
rect 6546 14764 6552 14816
rect 6604 14764 6610 14816
rect 10505 14807 10563 14813
rect 10505 14773 10517 14807
rect 10551 14804 10563 14807
rect 10870 14804 10876 14816
rect 10551 14776 10876 14804
rect 10551 14773 10563 14776
rect 10505 14767 10563 14773
rect 10870 14764 10876 14776
rect 10928 14764 10934 14816
rect 14734 14764 14740 14816
rect 14792 14804 14798 14816
rect 15749 14807 15807 14813
rect 15749 14804 15761 14807
rect 14792 14776 15761 14804
rect 14792 14764 14798 14776
rect 15749 14773 15761 14776
rect 15795 14773 15807 14807
rect 15856 14804 15884 14844
rect 15930 14832 15936 14884
rect 15988 14832 15994 14884
rect 16850 14832 16856 14884
rect 16908 14872 16914 14884
rect 18325 14875 18383 14881
rect 18325 14872 18337 14875
rect 16908 14844 18337 14872
rect 16908 14832 16914 14844
rect 18325 14841 18337 14844
rect 18371 14841 18383 14875
rect 18325 14835 18383 14841
rect 18892 14804 18920 14980
rect 19245 14977 19257 14980
rect 19291 14977 19303 15011
rect 19245 14971 19303 14977
rect 19426 14968 19432 15020
rect 19484 14968 19490 15020
rect 21453 15011 21511 15017
rect 21453 14977 21465 15011
rect 21499 15008 21511 15011
rect 21726 15008 21732 15020
rect 21499 14980 21732 15008
rect 21499 14977 21511 14980
rect 21453 14971 21511 14977
rect 21726 14968 21732 14980
rect 21784 15008 21790 15020
rect 22848 15017 22876 15048
rect 22281 15011 22339 15017
rect 22281 15008 22293 15011
rect 21784 14980 22293 15008
rect 21784 14968 21790 14980
rect 22281 14977 22293 14980
rect 22327 14977 22339 15011
rect 22281 14971 22339 14977
rect 22833 15011 22891 15017
rect 22833 14977 22845 15011
rect 22879 14977 22891 15011
rect 22833 14971 22891 14977
rect 19613 14943 19671 14949
rect 19613 14909 19625 14943
rect 19659 14940 19671 14943
rect 20070 14940 20076 14952
rect 19659 14912 20076 14940
rect 19659 14909 19671 14912
rect 19613 14903 19671 14909
rect 20070 14900 20076 14912
rect 20128 14940 20134 14952
rect 20530 14940 20536 14952
rect 20128 14912 20536 14940
rect 20128 14900 20134 14912
rect 20530 14900 20536 14912
rect 20588 14900 20594 14952
rect 22002 14900 22008 14952
rect 22060 14900 22066 14952
rect 22649 14943 22707 14949
rect 22649 14909 22661 14943
rect 22695 14909 22707 14943
rect 22649 14903 22707 14909
rect 21542 14832 21548 14884
rect 21600 14872 21606 14884
rect 22664 14872 22692 14903
rect 21600 14844 22692 14872
rect 21600 14832 21606 14844
rect 15856 14776 18920 14804
rect 20901 14807 20959 14813
rect 15749 14767 15807 14773
rect 20901 14773 20913 14807
rect 20947 14804 20959 14807
rect 21174 14804 21180 14816
rect 20947 14776 21180 14804
rect 20947 14773 20959 14776
rect 20901 14767 20959 14773
rect 21174 14764 21180 14776
rect 21232 14764 21238 14816
rect 1104 14714 23828 14736
rect 1104 14662 3790 14714
rect 3842 14662 3854 14714
rect 3906 14662 3918 14714
rect 3970 14662 3982 14714
rect 4034 14662 4046 14714
rect 4098 14662 9471 14714
rect 9523 14662 9535 14714
rect 9587 14662 9599 14714
rect 9651 14662 9663 14714
rect 9715 14662 9727 14714
rect 9779 14662 15152 14714
rect 15204 14662 15216 14714
rect 15268 14662 15280 14714
rect 15332 14662 15344 14714
rect 15396 14662 15408 14714
rect 15460 14662 20833 14714
rect 20885 14662 20897 14714
rect 20949 14662 20961 14714
rect 21013 14662 21025 14714
rect 21077 14662 21089 14714
rect 21141 14662 23828 14714
rect 1104 14640 23828 14662
rect 2314 14560 2320 14612
rect 2372 14560 2378 14612
rect 3326 14560 3332 14612
rect 3384 14600 3390 14612
rect 5077 14603 5135 14609
rect 5077 14600 5089 14603
rect 3384 14572 5089 14600
rect 3384 14560 3390 14572
rect 5077 14569 5089 14572
rect 5123 14569 5135 14603
rect 5077 14563 5135 14569
rect 6086 14560 6092 14612
rect 6144 14560 6150 14612
rect 7742 14560 7748 14612
rect 7800 14600 7806 14612
rect 9125 14603 9183 14609
rect 9125 14600 9137 14603
rect 7800 14572 9137 14600
rect 7800 14560 7806 14572
rect 9125 14569 9137 14572
rect 9171 14569 9183 14603
rect 9125 14563 9183 14569
rect 9214 14560 9220 14612
rect 9272 14600 9278 14612
rect 9272 14572 10916 14600
rect 9272 14560 9278 14572
rect 8202 14492 8208 14544
rect 8260 14532 8266 14544
rect 8260 14504 8340 14532
rect 8260 14492 8266 14504
rect 5166 14464 5172 14476
rect 2240 14436 4200 14464
rect 2240 14408 2268 14436
rect 1765 14399 1823 14405
rect 1765 14365 1777 14399
rect 1811 14396 1823 14399
rect 1854 14396 1860 14408
rect 1811 14368 1860 14396
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 1854 14356 1860 14368
rect 1912 14356 1918 14408
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14396 2191 14399
rect 2222 14396 2228 14408
rect 2179 14368 2228 14396
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 2222 14356 2228 14368
rect 2280 14356 2286 14408
rect 2866 14356 2872 14408
rect 2924 14396 2930 14408
rect 4172 14405 4200 14436
rect 4540 14436 5172 14464
rect 4540 14405 4568 14436
rect 5166 14424 5172 14436
rect 5224 14464 5230 14476
rect 8312 14464 8340 14504
rect 8662 14492 8668 14544
rect 8720 14532 8726 14544
rect 10413 14535 10471 14541
rect 8720 14504 9628 14532
rect 8720 14492 8726 14504
rect 5224 14436 7328 14464
rect 5224 14424 5230 14436
rect 3421 14399 3479 14405
rect 3421 14396 3433 14399
rect 2924 14368 3433 14396
rect 2924 14356 2930 14368
rect 3421 14365 3433 14368
rect 3467 14365 3479 14399
rect 3421 14359 3479 14365
rect 4157 14399 4215 14405
rect 4157 14365 4169 14399
rect 4203 14396 4215 14399
rect 4525 14399 4583 14405
rect 4203 14368 4476 14396
rect 4203 14365 4215 14368
rect 4157 14359 4215 14365
rect 1946 14288 1952 14340
rect 2004 14288 2010 14340
rect 2041 14331 2099 14337
rect 2041 14297 2053 14331
rect 2087 14328 2099 14331
rect 2682 14328 2688 14340
rect 2087 14300 2688 14328
rect 2087 14297 2099 14300
rect 2041 14291 2099 14297
rect 1670 14220 1676 14272
rect 1728 14260 1734 14272
rect 2056 14260 2084 14291
rect 2682 14288 2688 14300
rect 2740 14288 2746 14340
rect 3145 14331 3203 14337
rect 3145 14297 3157 14331
rect 3191 14328 3203 14331
rect 4249 14331 4307 14337
rect 4249 14328 4261 14331
rect 3191 14300 4261 14328
rect 3191 14297 3203 14300
rect 3145 14291 3203 14297
rect 4249 14297 4261 14300
rect 4295 14297 4307 14331
rect 4249 14291 4307 14297
rect 1728 14232 2084 14260
rect 1728 14220 1734 14232
rect 2222 14220 2228 14272
rect 2280 14260 2286 14272
rect 3160 14260 3188 14291
rect 2280 14232 3188 14260
rect 2280 14220 2286 14232
rect 3970 14220 3976 14272
rect 4028 14220 4034 14272
rect 4264 14260 4292 14291
rect 4338 14288 4344 14340
rect 4396 14288 4402 14340
rect 4448 14328 4476 14368
rect 4525 14365 4537 14399
rect 4571 14365 4583 14399
rect 4525 14359 4583 14365
rect 5261 14399 5319 14405
rect 5261 14365 5273 14399
rect 5307 14365 5319 14399
rect 5261 14359 5319 14365
rect 5276 14328 5304 14359
rect 5350 14356 5356 14408
rect 5408 14356 5414 14408
rect 5644 14405 5672 14436
rect 7300 14408 7328 14436
rect 8312 14436 9352 14464
rect 8215 14409 8273 14415
rect 5629 14399 5687 14405
rect 5629 14365 5641 14399
rect 5675 14365 5687 14399
rect 5629 14359 5687 14365
rect 5810 14356 5816 14408
rect 5868 14396 5874 14408
rect 6273 14399 6331 14405
rect 6273 14396 6285 14399
rect 5868 14368 6285 14396
rect 5868 14356 5874 14368
rect 6273 14365 6285 14368
rect 6319 14365 6331 14399
rect 6273 14359 6331 14365
rect 6638 14356 6644 14408
rect 6696 14356 6702 14408
rect 7282 14356 7288 14408
rect 7340 14396 7346 14408
rect 7340 14368 7696 14396
rect 7340 14356 7346 14368
rect 4448 14300 5304 14328
rect 4522 14260 4528 14272
rect 4264 14232 4528 14260
rect 4522 14220 4528 14232
rect 4580 14220 4586 14272
rect 5276 14260 5304 14300
rect 5442 14288 5448 14340
rect 5500 14288 5506 14340
rect 6362 14288 6368 14340
rect 6420 14288 6426 14340
rect 6454 14288 6460 14340
rect 6512 14288 6518 14340
rect 7558 14328 7564 14340
rect 7024 14300 7564 14328
rect 7024 14260 7052 14300
rect 7558 14288 7564 14300
rect 7616 14288 7622 14340
rect 7668 14328 7696 14368
rect 7834 14356 7840 14408
rect 7892 14356 7898 14408
rect 7929 14399 7987 14405
rect 7929 14365 7941 14399
rect 7975 14365 7987 14399
rect 7929 14359 7987 14365
rect 7944 14328 7972 14359
rect 8018 14356 8024 14408
rect 8076 14396 8082 14408
rect 8113 14399 8171 14405
rect 8113 14396 8125 14399
rect 8076 14368 8125 14396
rect 8076 14356 8082 14368
rect 8113 14365 8125 14368
rect 8159 14365 8171 14399
rect 8215 14375 8227 14409
rect 8261 14406 8273 14409
rect 8312 14406 8340 14436
rect 8261 14378 8340 14406
rect 9324 14405 9352 14436
rect 9309 14399 9367 14405
rect 8261 14375 8273 14378
rect 8215 14369 8273 14375
rect 8113 14359 8171 14365
rect 9309 14365 9321 14399
rect 9355 14365 9367 14399
rect 9600 14396 9628 14504
rect 10413 14501 10425 14535
rect 10459 14532 10471 14535
rect 10778 14532 10784 14544
rect 10459 14504 10784 14532
rect 10459 14501 10471 14504
rect 10413 14495 10471 14501
rect 10778 14492 10784 14504
rect 10836 14492 10842 14544
rect 9677 14399 9735 14405
rect 9677 14396 9689 14399
rect 9600 14368 9689 14396
rect 9309 14359 9367 14365
rect 9677 14365 9689 14368
rect 9723 14365 9735 14399
rect 9677 14359 9735 14365
rect 10134 14356 10140 14408
rect 10192 14396 10198 14408
rect 10689 14399 10747 14405
rect 10689 14396 10701 14399
rect 10192 14368 10701 14396
rect 10192 14356 10198 14368
rect 10689 14365 10701 14368
rect 10735 14365 10747 14399
rect 10888 14396 10916 14572
rect 11606 14560 11612 14612
rect 11664 14600 11670 14612
rect 11664 14572 12434 14600
rect 11664 14560 11670 14572
rect 12406 14532 12434 14572
rect 13262 14560 13268 14612
rect 13320 14600 13326 14612
rect 13633 14603 13691 14609
rect 13633 14600 13645 14603
rect 13320 14572 13645 14600
rect 13320 14560 13326 14572
rect 13633 14569 13645 14572
rect 13679 14600 13691 14603
rect 14553 14603 14611 14609
rect 13679 14572 14504 14600
rect 13679 14569 13691 14572
rect 13633 14563 13691 14569
rect 14274 14532 14280 14544
rect 12406 14504 14280 14532
rect 14274 14492 14280 14504
rect 14332 14492 14338 14544
rect 11609 14467 11667 14473
rect 11609 14433 11621 14467
rect 11655 14464 11667 14467
rect 11882 14464 11888 14476
rect 11655 14436 11888 14464
rect 11655 14433 11667 14436
rect 11609 14427 11667 14433
rect 11882 14424 11888 14436
rect 11940 14424 11946 14476
rect 12713 14467 12771 14473
rect 12713 14433 12725 14467
rect 12759 14464 12771 14467
rect 13630 14464 13636 14476
rect 12759 14436 13636 14464
rect 12759 14433 12771 14436
rect 12713 14427 12771 14433
rect 13630 14424 13636 14436
rect 13688 14424 13694 14476
rect 14476 14464 14504 14572
rect 14553 14569 14565 14603
rect 14599 14600 14611 14603
rect 14642 14600 14648 14612
rect 14599 14572 14648 14600
rect 14599 14569 14611 14572
rect 14553 14563 14611 14569
rect 14642 14560 14648 14572
rect 14700 14560 14706 14612
rect 15470 14560 15476 14612
rect 15528 14600 15534 14612
rect 15657 14603 15715 14609
rect 15657 14600 15669 14603
rect 15528 14572 15669 14600
rect 15528 14560 15534 14572
rect 15657 14569 15669 14572
rect 15703 14569 15715 14603
rect 15657 14563 15715 14569
rect 15838 14560 15844 14612
rect 15896 14600 15902 14612
rect 16114 14600 16120 14612
rect 15896 14572 16120 14600
rect 15896 14560 15902 14572
rect 16114 14560 16120 14572
rect 16172 14560 16178 14612
rect 19978 14560 19984 14612
rect 20036 14600 20042 14612
rect 20073 14603 20131 14609
rect 20073 14600 20085 14603
rect 20036 14572 20085 14600
rect 20036 14560 20042 14572
rect 20073 14569 20085 14572
rect 20119 14569 20131 14603
rect 21818 14600 21824 14612
rect 20073 14563 20131 14569
rect 20180 14572 21824 14600
rect 18874 14492 18880 14544
rect 18932 14532 18938 14544
rect 20180 14532 20208 14572
rect 21818 14560 21824 14572
rect 21876 14560 21882 14612
rect 22186 14560 22192 14612
rect 22244 14600 22250 14612
rect 22281 14603 22339 14609
rect 22281 14600 22293 14603
rect 22244 14572 22293 14600
rect 22244 14560 22250 14572
rect 22281 14569 22293 14572
rect 22327 14569 22339 14603
rect 22281 14563 22339 14569
rect 18932 14504 20208 14532
rect 18932 14492 18938 14504
rect 20438 14492 20444 14544
rect 20496 14532 20502 14544
rect 20496 14504 20668 14532
rect 20496 14492 20502 14504
rect 14921 14467 14979 14473
rect 14921 14464 14933 14467
rect 14476 14436 14933 14464
rect 14921 14433 14933 14436
rect 14967 14433 14979 14467
rect 16298 14464 16304 14476
rect 14921 14427 14979 14433
rect 15672 14436 16304 14464
rect 11698 14396 11704 14408
rect 10888 14368 11704 14396
rect 10689 14359 10747 14365
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 11790 14356 11796 14408
rect 11848 14396 11854 14408
rect 11977 14399 12035 14405
rect 11977 14396 11989 14399
rect 11848 14368 11989 14396
rect 11848 14356 11854 14368
rect 11977 14365 11989 14368
rect 12023 14365 12035 14399
rect 11977 14359 12035 14365
rect 12069 14399 12127 14405
rect 12069 14365 12081 14399
rect 12115 14396 12127 14399
rect 14090 14396 14096 14408
rect 12115 14368 14096 14396
rect 12115 14365 12127 14368
rect 12069 14359 12127 14365
rect 14090 14356 14096 14368
rect 14148 14356 14154 14408
rect 14734 14356 14740 14408
rect 14792 14356 14798 14408
rect 15672 14405 15700 14436
rect 16298 14424 16304 14436
rect 16356 14424 16362 14476
rect 17126 14424 17132 14476
rect 17184 14464 17190 14476
rect 17184 14436 17448 14464
rect 17184 14424 17190 14436
rect 15657 14399 15715 14405
rect 15657 14365 15669 14399
rect 15703 14365 15715 14399
rect 15657 14359 15715 14365
rect 15933 14399 15991 14405
rect 15933 14365 15945 14399
rect 15979 14396 15991 14399
rect 16850 14396 16856 14408
rect 15979 14368 16856 14396
rect 15979 14365 15991 14368
rect 15933 14359 15991 14365
rect 16850 14356 16856 14368
rect 16908 14356 16914 14408
rect 17420 14396 17448 14436
rect 19058 14424 19064 14476
rect 19116 14464 19122 14476
rect 20640 14464 20668 14504
rect 20714 14492 20720 14544
rect 20772 14532 20778 14544
rect 20772 14504 21772 14532
rect 20772 14492 20778 14504
rect 20990 14464 20996 14476
rect 19116 14436 20576 14464
rect 20640 14436 20996 14464
rect 19116 14424 19122 14436
rect 19429 14399 19487 14405
rect 19429 14396 19441 14399
rect 17420 14368 19441 14396
rect 19429 14365 19441 14368
rect 19475 14365 19487 14399
rect 19429 14359 19487 14365
rect 19521 14399 19579 14405
rect 19521 14365 19533 14399
rect 19567 14365 19579 14399
rect 19521 14359 19579 14365
rect 7668 14300 7972 14328
rect 5276 14232 7052 14260
rect 7098 14220 7104 14272
rect 7156 14260 7162 14272
rect 7653 14263 7711 14269
rect 7653 14260 7665 14263
rect 7156 14232 7665 14260
rect 7156 14220 7162 14232
rect 7653 14229 7665 14232
rect 7699 14229 7711 14263
rect 7944 14260 7972 14300
rect 8478 14288 8484 14340
rect 8536 14328 8542 14340
rect 9401 14331 9459 14337
rect 9401 14328 9413 14331
rect 8536 14300 9413 14328
rect 8536 14288 8542 14300
rect 9401 14297 9413 14300
rect 9447 14297 9459 14331
rect 9401 14291 9459 14297
rect 9493 14331 9551 14337
rect 9493 14297 9505 14331
rect 9539 14297 9551 14331
rect 9493 14291 9551 14297
rect 8662 14260 8668 14272
rect 7944 14232 8668 14260
rect 7653 14223 7711 14229
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 9214 14220 9220 14272
rect 9272 14260 9278 14272
rect 9508 14260 9536 14291
rect 10870 14288 10876 14340
rect 10928 14288 10934 14340
rect 10965 14331 11023 14337
rect 10965 14297 10977 14331
rect 11011 14328 11023 14331
rect 11146 14328 11152 14340
rect 11011 14300 11152 14328
rect 11011 14297 11023 14300
rect 10965 14291 11023 14297
rect 11146 14288 11152 14300
rect 11204 14288 11210 14340
rect 13906 14288 13912 14340
rect 13964 14328 13970 14340
rect 15102 14328 15108 14340
rect 13964 14300 15108 14328
rect 13964 14288 13970 14300
rect 15102 14288 15108 14300
rect 15160 14288 15166 14340
rect 15562 14288 15568 14340
rect 15620 14328 15626 14340
rect 15749 14331 15807 14337
rect 15749 14328 15761 14331
rect 15620 14300 15761 14328
rect 15620 14288 15626 14300
rect 15749 14297 15761 14300
rect 15795 14297 15807 14331
rect 19536 14328 19564 14359
rect 19886 14356 19892 14408
rect 19944 14356 19950 14408
rect 15749 14291 15807 14297
rect 15948 14300 19564 14328
rect 19705 14331 19763 14337
rect 15948 14272 15976 14300
rect 19705 14297 19717 14331
rect 19751 14297 19763 14331
rect 19705 14291 19763 14297
rect 19797 14331 19855 14337
rect 19797 14297 19809 14331
rect 19843 14328 19855 14331
rect 20438 14328 20444 14340
rect 19843 14300 20444 14328
rect 19843 14297 19855 14300
rect 19797 14291 19855 14297
rect 9272 14232 9536 14260
rect 9272 14220 9278 14232
rect 13814 14220 13820 14272
rect 13872 14260 13878 14272
rect 14550 14260 14556 14272
rect 13872 14232 14556 14260
rect 13872 14220 13878 14232
rect 14550 14220 14556 14232
rect 14608 14220 14614 14272
rect 15930 14220 15936 14272
rect 15988 14220 15994 14272
rect 18601 14263 18659 14269
rect 18601 14229 18613 14263
rect 18647 14260 18659 14263
rect 18690 14260 18696 14272
rect 18647 14232 18696 14260
rect 18647 14229 18659 14232
rect 18601 14223 18659 14229
rect 18690 14220 18696 14232
rect 18748 14220 18754 14272
rect 19334 14220 19340 14272
rect 19392 14260 19398 14272
rect 19610 14260 19616 14272
rect 19392 14232 19616 14260
rect 19392 14220 19398 14232
rect 19610 14220 19616 14232
rect 19668 14260 19674 14272
rect 19720 14260 19748 14291
rect 20438 14288 20444 14300
rect 20496 14288 20502 14340
rect 20548 14328 20576 14436
rect 20990 14424 20996 14436
rect 21048 14424 21054 14476
rect 21634 14356 21640 14408
rect 21692 14356 21698 14408
rect 21744 14405 21772 14504
rect 21730 14399 21788 14405
rect 21730 14365 21742 14399
rect 21776 14365 21788 14399
rect 21730 14359 21788 14365
rect 22002 14356 22008 14408
rect 22060 14356 22066 14408
rect 22143 14399 22201 14405
rect 22143 14365 22155 14399
rect 22189 14396 22201 14399
rect 22278 14396 22284 14408
rect 22189 14368 22284 14396
rect 22189 14365 22201 14368
rect 22143 14359 22201 14365
rect 22278 14356 22284 14368
rect 22336 14356 22342 14408
rect 22925 14399 22983 14405
rect 22925 14365 22937 14399
rect 22971 14396 22983 14399
rect 23198 14396 23204 14408
rect 22971 14368 23204 14396
rect 22971 14365 22983 14368
rect 22925 14359 22983 14365
rect 23198 14356 23204 14368
rect 23256 14356 23262 14408
rect 20548 14300 21036 14328
rect 19668 14232 19748 14260
rect 19668 14220 19674 14232
rect 20898 14220 20904 14272
rect 20956 14220 20962 14272
rect 21008 14260 21036 14300
rect 21450 14288 21456 14340
rect 21508 14328 21514 14340
rect 21913 14331 21971 14337
rect 21913 14328 21925 14331
rect 21508 14300 21925 14328
rect 21508 14288 21514 14300
rect 21913 14297 21925 14300
rect 21959 14297 21971 14331
rect 21913 14291 21971 14297
rect 22020 14260 22048 14356
rect 21008 14232 22048 14260
rect 22830 14220 22836 14272
rect 22888 14220 22894 14272
rect 1104 14170 23987 14192
rect 1104 14118 6630 14170
rect 6682 14118 6694 14170
rect 6746 14118 6758 14170
rect 6810 14118 6822 14170
rect 6874 14118 6886 14170
rect 6938 14118 12311 14170
rect 12363 14118 12375 14170
rect 12427 14118 12439 14170
rect 12491 14118 12503 14170
rect 12555 14118 12567 14170
rect 12619 14118 17992 14170
rect 18044 14118 18056 14170
rect 18108 14118 18120 14170
rect 18172 14118 18184 14170
rect 18236 14118 18248 14170
rect 18300 14118 23673 14170
rect 23725 14118 23737 14170
rect 23789 14118 23801 14170
rect 23853 14118 23865 14170
rect 23917 14118 23929 14170
rect 23981 14118 23987 14170
rect 1104 14096 23987 14118
rect 2038 14016 2044 14068
rect 2096 14056 2102 14068
rect 2133 14059 2191 14065
rect 2133 14056 2145 14059
rect 2096 14028 2145 14056
rect 2096 14016 2102 14028
rect 2133 14025 2145 14028
rect 2179 14025 2191 14059
rect 2133 14019 2191 14025
rect 2866 14016 2872 14068
rect 2924 14016 2930 14068
rect 4430 14016 4436 14068
rect 4488 14056 4494 14068
rect 4709 14059 4767 14065
rect 4709 14056 4721 14059
rect 4488 14028 4721 14056
rect 4488 14016 4494 14028
rect 4709 14025 4721 14028
rect 4755 14056 4767 14059
rect 4798 14056 4804 14068
rect 4755 14028 4804 14056
rect 4755 14025 4767 14028
rect 4709 14019 4767 14025
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 5258 14016 5264 14068
rect 5316 14016 5322 14068
rect 5721 14059 5779 14065
rect 5721 14025 5733 14059
rect 5767 14056 5779 14059
rect 6454 14056 6460 14068
rect 5767 14028 6460 14056
rect 5767 14025 5779 14028
rect 5721 14019 5779 14025
rect 6454 14016 6460 14028
rect 6512 14056 6518 14068
rect 7193 14059 7251 14065
rect 7193 14056 7205 14059
rect 6512 14028 7205 14056
rect 6512 14016 6518 14028
rect 7193 14025 7205 14028
rect 7239 14025 7251 14059
rect 7193 14019 7251 14025
rect 7558 14016 7564 14068
rect 7616 14056 7622 14068
rect 8202 14056 8208 14068
rect 7616 14028 8208 14056
rect 7616 14016 7622 14028
rect 8202 14016 8208 14028
rect 8260 14016 8266 14068
rect 11790 14016 11796 14068
rect 11848 14016 11854 14068
rect 12526 14016 12532 14068
rect 12584 14056 12590 14068
rect 12897 14059 12955 14065
rect 12897 14056 12909 14059
rect 12584 14028 12909 14056
rect 12584 14016 12590 14028
rect 12897 14025 12909 14028
rect 12943 14056 12955 14059
rect 13262 14056 13268 14068
rect 12943 14028 13268 14056
rect 12943 14025 12955 14028
rect 12897 14019 12955 14025
rect 13262 14016 13268 14028
rect 13320 14016 13326 14068
rect 13633 14059 13691 14065
rect 13633 14025 13645 14059
rect 13679 14056 13691 14059
rect 14182 14056 14188 14068
rect 13679 14028 14188 14056
rect 13679 14025 13691 14028
rect 13633 14019 13691 14025
rect 14182 14016 14188 14028
rect 14240 14056 14246 14068
rect 16390 14056 16396 14068
rect 14240 14028 16396 14056
rect 14240 14016 14246 14028
rect 16390 14016 16396 14028
rect 16448 14016 16454 14068
rect 16482 14016 16488 14068
rect 16540 14056 16546 14068
rect 16540 14028 17448 14056
rect 16540 14016 16546 14028
rect 3050 13948 3056 14000
rect 3108 13988 3114 14000
rect 5629 13991 5687 13997
rect 3108 13960 4292 13988
rect 3108 13948 3114 13960
rect 2406 13880 2412 13932
rect 2464 13880 2470 13932
rect 3970 13880 3976 13932
rect 4028 13929 4034 13932
rect 4264 13929 4292 13960
rect 5629 13957 5641 13991
rect 5675 13988 5687 13991
rect 5810 13988 5816 14000
rect 5675 13960 5816 13988
rect 5675 13957 5687 13960
rect 5629 13951 5687 13957
rect 5810 13948 5816 13960
rect 5868 13988 5874 14000
rect 6733 13991 6791 13997
rect 6733 13988 6745 13991
rect 5868 13960 6745 13988
rect 5868 13948 5874 13960
rect 6733 13957 6745 13960
rect 6779 13957 6791 13991
rect 6733 13951 6791 13957
rect 7374 13948 7380 14000
rect 7432 13988 7438 14000
rect 7742 13988 7748 14000
rect 7432 13960 7748 13988
rect 7432 13948 7438 13960
rect 7742 13948 7748 13960
rect 7800 13988 7806 14000
rect 7800 13960 8892 13988
rect 7800 13948 7806 13960
rect 4028 13920 4040 13929
rect 4249 13923 4307 13929
rect 4028 13892 4073 13920
rect 4028 13883 4040 13892
rect 4249 13889 4261 13923
rect 4295 13889 4307 13923
rect 4249 13883 4307 13889
rect 4028 13880 4034 13883
rect 8294 13880 8300 13932
rect 8352 13880 8358 13932
rect 8864 13929 8892 13960
rect 13078 13948 13084 14000
rect 13136 13988 13142 14000
rect 13136 13960 14412 13988
rect 13136 13948 13142 13960
rect 8849 13923 8907 13929
rect 8849 13889 8861 13923
rect 8895 13889 8907 13923
rect 8849 13883 8907 13889
rect 11698 13880 11704 13932
rect 11756 13880 11762 13932
rect 11882 13880 11888 13932
rect 11940 13880 11946 13932
rect 14001 13923 14059 13929
rect 14001 13889 14013 13923
rect 14047 13920 14059 13923
rect 14090 13920 14096 13932
rect 14047 13892 14096 13920
rect 14047 13889 14059 13892
rect 14001 13883 14059 13889
rect 14090 13880 14096 13892
rect 14148 13880 14154 13932
rect 14384 13929 14412 13960
rect 14826 13948 14832 14000
rect 14884 13988 14890 14000
rect 14884 13960 17356 13988
rect 14884 13948 14890 13960
rect 14369 13923 14427 13929
rect 14369 13889 14381 13923
rect 14415 13920 14427 13923
rect 14918 13920 14924 13932
rect 14415 13892 14924 13920
rect 14415 13889 14427 13892
rect 14369 13883 14427 13889
rect 14918 13880 14924 13892
rect 14976 13880 14982 13932
rect 15102 13880 15108 13932
rect 15160 13920 15166 13932
rect 15657 13923 15715 13929
rect 15657 13920 15669 13923
rect 15160 13892 15669 13920
rect 15160 13880 15166 13892
rect 15657 13889 15669 13892
rect 15703 13920 15715 13923
rect 16206 13920 16212 13932
rect 15703 13892 16212 13920
rect 15703 13889 15715 13892
rect 15657 13883 15715 13889
rect 16206 13880 16212 13892
rect 16264 13880 16270 13932
rect 17037 13923 17095 13929
rect 17037 13889 17049 13923
rect 17083 13889 17095 13923
rect 17037 13883 17095 13889
rect 2130 13812 2136 13864
rect 2188 13812 2194 13864
rect 5813 13855 5871 13861
rect 5813 13821 5825 13855
rect 5859 13821 5871 13855
rect 5813 13815 5871 13821
rect 4614 13744 4620 13796
rect 4672 13784 4678 13796
rect 5534 13784 5540 13796
rect 4672 13756 5540 13784
rect 4672 13744 4678 13756
rect 5534 13744 5540 13756
rect 5592 13784 5598 13796
rect 5828 13784 5856 13815
rect 11146 13812 11152 13864
rect 11204 13852 11210 13864
rect 12066 13852 12072 13864
rect 11204 13824 12072 13852
rect 11204 13812 11210 13824
rect 12066 13812 12072 13824
rect 12124 13812 12130 13864
rect 13906 13812 13912 13864
rect 13964 13812 13970 13864
rect 14274 13812 14280 13864
rect 14332 13852 14338 13864
rect 15010 13852 15016 13864
rect 14332 13824 15016 13852
rect 14332 13812 14338 13824
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 15470 13812 15476 13864
rect 15528 13852 15534 13864
rect 17052 13852 17080 13883
rect 17126 13880 17132 13932
rect 17184 13880 17190 13932
rect 17328 13929 17356 13960
rect 17420 13929 17448 14028
rect 20254 14016 20260 14068
rect 20312 14056 20318 14068
rect 20441 14059 20499 14065
rect 20441 14056 20453 14059
rect 20312 14028 20453 14056
rect 20312 14016 20318 14028
rect 20441 14025 20453 14028
rect 20487 14025 20499 14059
rect 20441 14019 20499 14025
rect 20530 14016 20536 14068
rect 20588 14056 20594 14068
rect 20588 14028 21680 14056
rect 20588 14016 20594 14028
rect 21652 13988 21680 14028
rect 21818 14016 21824 14068
rect 21876 14056 21882 14068
rect 22097 14059 22155 14065
rect 22097 14056 22109 14059
rect 21876 14028 22109 14056
rect 21876 14016 21882 14028
rect 22097 14025 22109 14028
rect 22143 14025 22155 14059
rect 22097 14019 22155 14025
rect 20180 13960 21588 13988
rect 21652 13960 22048 13988
rect 17313 13923 17371 13929
rect 17313 13889 17325 13923
rect 17359 13889 17371 13923
rect 17313 13883 17371 13889
rect 17405 13923 17463 13929
rect 17405 13889 17417 13923
rect 17451 13920 17463 13923
rect 19794 13920 19800 13932
rect 17451 13892 19800 13920
rect 17451 13889 17463 13892
rect 17405 13883 17463 13889
rect 19794 13880 19800 13892
rect 19852 13880 19858 13932
rect 19978 13880 19984 13932
rect 20036 13880 20042 13932
rect 20070 13880 20076 13932
rect 20128 13880 20134 13932
rect 20180 13929 20208 13960
rect 20165 13923 20223 13929
rect 20165 13889 20177 13923
rect 20211 13889 20223 13923
rect 20165 13883 20223 13889
rect 21085 13923 21143 13929
rect 21085 13889 21097 13923
rect 21131 13920 21143 13923
rect 21174 13920 21180 13932
rect 21131 13892 21180 13920
rect 21131 13889 21143 13892
rect 21085 13883 21143 13889
rect 21174 13880 21180 13892
rect 21232 13880 21238 13932
rect 21269 13923 21327 13929
rect 21269 13889 21281 13923
rect 21315 13889 21327 13923
rect 21269 13883 21327 13889
rect 19242 13852 19248 13864
rect 15528 13824 16252 13852
rect 15528 13812 15534 13824
rect 5592 13756 5856 13784
rect 5592 13744 5598 13756
rect 7098 13744 7104 13796
rect 7156 13744 7162 13796
rect 11514 13744 11520 13796
rect 11572 13784 11578 13796
rect 11698 13784 11704 13796
rect 11572 13756 11704 13784
rect 11572 13744 11578 13756
rect 11698 13744 11704 13756
rect 11756 13744 11762 13796
rect 16224 13793 16252 13824
rect 16776 13824 16988 13852
rect 17052 13824 19248 13852
rect 16209 13787 16267 13793
rect 16209 13753 16221 13787
rect 16255 13784 16267 13787
rect 16776 13784 16804 13824
rect 16255 13756 16804 13784
rect 16255 13753 16267 13756
rect 16209 13747 16267 13753
rect 16850 13744 16856 13796
rect 16908 13744 16914 13796
rect 16960 13784 16988 13824
rect 19242 13812 19248 13824
rect 19300 13812 19306 13864
rect 21284 13796 21312 13883
rect 21453 13855 21511 13861
rect 21453 13821 21465 13855
rect 21499 13821 21511 13855
rect 21560 13852 21588 13960
rect 22020 13929 22048 13960
rect 22005 13923 22063 13929
rect 22005 13889 22017 13923
rect 22051 13889 22063 13923
rect 22005 13883 22063 13889
rect 21560 13824 22048 13852
rect 21453 13815 21511 13821
rect 18414 13784 18420 13796
rect 16960 13756 18420 13784
rect 18414 13744 18420 13756
rect 18472 13784 18478 13796
rect 18598 13784 18604 13796
rect 18472 13756 18604 13784
rect 18472 13744 18478 13756
rect 18598 13744 18604 13756
rect 18656 13784 18662 13796
rect 20898 13784 20904 13796
rect 18656 13756 20904 13784
rect 18656 13744 18662 13756
rect 20898 13744 20904 13756
rect 20956 13744 20962 13796
rect 20990 13744 20996 13796
rect 21048 13784 21054 13796
rect 21266 13784 21272 13796
rect 21048 13756 21272 13784
rect 21048 13744 21054 13756
rect 21266 13744 21272 13756
rect 21324 13744 21330 13796
rect 2317 13719 2375 13725
rect 2317 13685 2329 13719
rect 2363 13716 2375 13719
rect 2774 13716 2780 13728
rect 2363 13688 2780 13716
rect 2363 13685 2375 13688
rect 2317 13679 2375 13685
rect 2774 13676 2780 13688
rect 2832 13676 2838 13728
rect 5902 13676 5908 13728
rect 5960 13716 5966 13728
rect 6454 13716 6460 13728
rect 5960 13688 6460 13716
rect 5960 13676 5966 13688
rect 6454 13676 6460 13688
rect 6512 13676 6518 13728
rect 20916 13716 20944 13744
rect 21468 13716 21496 13815
rect 21910 13716 21916 13728
rect 20916 13688 21916 13716
rect 21910 13676 21916 13688
rect 21968 13676 21974 13728
rect 22020 13716 22048 13824
rect 22094 13744 22100 13796
rect 22152 13784 22158 13796
rect 22465 13787 22523 13793
rect 22465 13784 22477 13787
rect 22152 13756 22477 13784
rect 22152 13744 22158 13756
rect 22465 13753 22477 13756
rect 22511 13753 22523 13787
rect 22465 13747 22523 13753
rect 22186 13716 22192 13728
rect 22020 13688 22192 13716
rect 22186 13676 22192 13688
rect 22244 13716 22250 13728
rect 22281 13719 22339 13725
rect 22281 13716 22293 13719
rect 22244 13688 22293 13716
rect 22244 13676 22250 13688
rect 22281 13685 22293 13688
rect 22327 13685 22339 13719
rect 22281 13679 22339 13685
rect 22370 13676 22376 13728
rect 22428 13676 22434 13728
rect 22738 13676 22744 13728
rect 22796 13676 22802 13728
rect 1104 13626 23828 13648
rect 1104 13574 3790 13626
rect 3842 13574 3854 13626
rect 3906 13574 3918 13626
rect 3970 13574 3982 13626
rect 4034 13574 4046 13626
rect 4098 13574 9471 13626
rect 9523 13574 9535 13626
rect 9587 13574 9599 13626
rect 9651 13574 9663 13626
rect 9715 13574 9727 13626
rect 9779 13574 15152 13626
rect 15204 13574 15216 13626
rect 15268 13574 15280 13626
rect 15332 13574 15344 13626
rect 15396 13574 15408 13626
rect 15460 13574 20833 13626
rect 20885 13574 20897 13626
rect 20949 13574 20961 13626
rect 21013 13574 21025 13626
rect 21077 13574 21089 13626
rect 21141 13574 23828 13626
rect 1104 13552 23828 13574
rect 4157 13515 4215 13521
rect 4157 13481 4169 13515
rect 4203 13512 4215 13515
rect 5442 13512 5448 13524
rect 4203 13484 5448 13512
rect 4203 13481 4215 13484
rect 4157 13475 4215 13481
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 5902 13472 5908 13524
rect 5960 13512 5966 13524
rect 6089 13515 6147 13521
rect 6089 13512 6101 13515
rect 5960 13484 6101 13512
rect 5960 13472 5966 13484
rect 6089 13481 6101 13484
rect 6135 13481 6147 13515
rect 6089 13475 6147 13481
rect 6825 13515 6883 13521
rect 6825 13481 6837 13515
rect 6871 13512 6883 13515
rect 7006 13512 7012 13524
rect 6871 13484 7012 13512
rect 6871 13481 6883 13484
rect 6825 13475 6883 13481
rect 7006 13472 7012 13484
rect 7064 13472 7070 13524
rect 7469 13515 7527 13521
rect 7469 13481 7481 13515
rect 7515 13512 7527 13515
rect 9214 13512 9220 13524
rect 7515 13484 9220 13512
rect 7515 13481 7527 13484
rect 7469 13475 7527 13481
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 12802 13472 12808 13524
rect 12860 13472 12866 13524
rect 13170 13472 13176 13524
rect 13228 13512 13234 13524
rect 13630 13512 13636 13524
rect 13228 13484 13636 13512
rect 13228 13472 13234 13484
rect 13630 13472 13636 13484
rect 13688 13472 13694 13524
rect 14182 13472 14188 13524
rect 14240 13512 14246 13524
rect 14642 13512 14648 13524
rect 14240 13484 14648 13512
rect 14240 13472 14246 13484
rect 14642 13472 14648 13484
rect 14700 13472 14706 13524
rect 14826 13472 14832 13524
rect 14884 13472 14890 13524
rect 14918 13472 14924 13524
rect 14976 13512 14982 13524
rect 15289 13515 15347 13521
rect 15289 13512 15301 13515
rect 14976 13484 15301 13512
rect 14976 13472 14982 13484
rect 15289 13481 15301 13484
rect 15335 13481 15347 13515
rect 15289 13475 15347 13481
rect 15378 13472 15384 13524
rect 15436 13512 15442 13524
rect 16022 13512 16028 13524
rect 15436 13484 16028 13512
rect 15436 13472 15442 13484
rect 16022 13472 16028 13484
rect 16080 13472 16086 13524
rect 16853 13515 16911 13521
rect 16853 13481 16865 13515
rect 16899 13512 16911 13515
rect 17034 13512 17040 13524
rect 16899 13484 17040 13512
rect 16899 13481 16911 13484
rect 16853 13475 16911 13481
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 19242 13472 19248 13524
rect 19300 13512 19306 13524
rect 19981 13515 20039 13521
rect 19981 13512 19993 13515
rect 19300 13484 19993 13512
rect 19300 13472 19306 13484
rect 19981 13481 19993 13484
rect 20027 13481 20039 13515
rect 22922 13512 22928 13524
rect 19981 13475 20039 13481
rect 22066 13484 22928 13512
rect 2222 13444 2228 13456
rect 1872 13416 2228 13444
rect 1872 13385 1900 13416
rect 2222 13404 2228 13416
rect 2280 13404 2286 13456
rect 3694 13404 3700 13456
rect 3752 13444 3758 13456
rect 4709 13447 4767 13453
rect 4709 13444 4721 13447
rect 3752 13416 4721 13444
rect 3752 13404 3758 13416
rect 4709 13413 4721 13416
rect 4755 13413 4767 13447
rect 4709 13407 4767 13413
rect 4798 13404 4804 13456
rect 4856 13444 4862 13456
rect 4856 13416 5212 13444
rect 4856 13404 4862 13416
rect 1857 13379 1915 13385
rect 1857 13345 1869 13379
rect 1903 13345 1915 13379
rect 1857 13339 1915 13345
rect 2130 13336 2136 13388
rect 2188 13376 2194 13388
rect 5184 13376 5212 13416
rect 7926 13404 7932 13456
rect 7984 13444 7990 13456
rect 8021 13447 8079 13453
rect 8021 13444 8033 13447
rect 7984 13416 8033 13444
rect 7984 13404 7990 13416
rect 8021 13413 8033 13416
rect 8067 13413 8079 13447
rect 8021 13407 8079 13413
rect 12713 13447 12771 13453
rect 12713 13413 12725 13447
rect 12759 13444 12771 13447
rect 14734 13444 14740 13456
rect 12759 13416 14740 13444
rect 12759 13413 12771 13416
rect 12713 13407 12771 13413
rect 14734 13404 14740 13416
rect 14792 13404 14798 13456
rect 16040 13444 16068 13472
rect 16040 13416 17816 13444
rect 5261 13379 5319 13385
rect 5261 13376 5273 13379
rect 2188 13348 4108 13376
rect 5184 13348 5273 13376
rect 2188 13336 2194 13348
rect 1670 13268 1676 13320
rect 1728 13268 1734 13320
rect 2041 13311 2099 13317
rect 2041 13277 2053 13311
rect 2087 13308 2099 13311
rect 2314 13308 2320 13320
rect 2087 13280 2320 13308
rect 2087 13277 2099 13280
rect 2041 13271 2099 13277
rect 2314 13268 2320 13280
rect 2372 13268 2378 13320
rect 2406 13268 2412 13320
rect 2464 13308 2470 13320
rect 2961 13311 3019 13317
rect 2961 13308 2973 13311
rect 2464 13280 2973 13308
rect 2464 13268 2470 13280
rect 2961 13277 2973 13280
rect 3007 13277 3019 13311
rect 2961 13271 3019 13277
rect 3234 13268 3240 13320
rect 3292 13268 3298 13320
rect 4080 13317 4108 13348
rect 5261 13345 5273 13348
rect 5307 13345 5319 13379
rect 5261 13339 5319 13345
rect 7650 13336 7656 13388
rect 7708 13376 7714 13388
rect 11977 13379 12035 13385
rect 11977 13376 11989 13379
rect 7708 13348 8616 13376
rect 7708 13336 7714 13348
rect 4065 13311 4123 13317
rect 4065 13277 4077 13311
rect 4111 13277 4123 13311
rect 4065 13271 4123 13277
rect 1854 13200 1860 13252
rect 1912 13240 1918 13252
rect 3053 13243 3111 13249
rect 3053 13240 3065 13243
rect 1912 13212 3065 13240
rect 1912 13200 1918 13212
rect 3053 13209 3065 13212
rect 3099 13240 3111 13243
rect 4080 13240 4108 13271
rect 4246 13268 4252 13320
rect 4304 13268 4310 13320
rect 4890 13268 4896 13320
rect 4948 13308 4954 13320
rect 5077 13311 5135 13317
rect 5077 13308 5089 13311
rect 4948 13280 5089 13308
rect 4948 13268 4954 13280
rect 5077 13277 5089 13280
rect 5123 13277 5135 13311
rect 5077 13271 5135 13277
rect 5169 13311 5227 13317
rect 5169 13277 5181 13311
rect 5215 13308 5227 13311
rect 5534 13308 5540 13320
rect 5215 13280 5540 13308
rect 5215 13277 5227 13280
rect 5169 13271 5227 13277
rect 5534 13268 5540 13280
rect 5592 13308 5598 13320
rect 6546 13308 6552 13320
rect 5592 13280 6552 13308
rect 5592 13268 5598 13280
rect 6546 13268 6552 13280
rect 6604 13268 6610 13320
rect 7006 13268 7012 13320
rect 7064 13308 7070 13320
rect 7377 13311 7435 13317
rect 7377 13308 7389 13311
rect 7064 13280 7389 13308
rect 7064 13268 7070 13280
rect 7377 13277 7389 13280
rect 7423 13277 7435 13311
rect 7377 13271 7435 13277
rect 7561 13311 7619 13317
rect 7561 13277 7573 13311
rect 7607 13277 7619 13311
rect 7561 13271 7619 13277
rect 6273 13243 6331 13249
rect 3099 13212 4025 13240
rect 4080 13212 6224 13240
rect 3099 13209 3111 13212
rect 3053 13203 3111 13209
rect 1762 13132 1768 13184
rect 1820 13132 1826 13184
rect 1949 13175 2007 13181
rect 1949 13141 1961 13175
rect 1995 13172 2007 13175
rect 2038 13172 2044 13184
rect 1995 13144 2044 13172
rect 1995 13141 2007 13144
rect 1949 13135 2007 13141
rect 2038 13132 2044 13144
rect 2096 13132 2102 13184
rect 3418 13132 3424 13184
rect 3476 13132 3482 13184
rect 3997 13172 4025 13212
rect 5166 13172 5172 13184
rect 3997 13144 5172 13172
rect 5166 13132 5172 13144
rect 5224 13132 5230 13184
rect 5810 13132 5816 13184
rect 5868 13172 5874 13184
rect 6086 13181 6092 13184
rect 5905 13175 5963 13181
rect 5905 13172 5917 13175
rect 5868 13144 5917 13172
rect 5868 13132 5874 13144
rect 5905 13141 5917 13144
rect 5951 13141 5963 13175
rect 5905 13135 5963 13141
rect 6073 13175 6092 13181
rect 6073 13141 6085 13175
rect 6073 13135 6092 13141
rect 6086 13132 6092 13135
rect 6144 13132 6150 13184
rect 6196 13172 6224 13212
rect 6273 13209 6285 13243
rect 6319 13240 6331 13243
rect 7282 13240 7288 13252
rect 6319 13212 7288 13240
rect 6319 13209 6331 13212
rect 6273 13203 6331 13209
rect 7282 13200 7288 13212
rect 7340 13200 7346 13252
rect 7576 13172 7604 13271
rect 8202 13268 8208 13320
rect 8260 13268 8266 13320
rect 8588 13317 8616 13348
rect 10888 13348 11989 13376
rect 8297 13311 8355 13317
rect 8297 13277 8309 13311
rect 8343 13308 8355 13311
rect 8573 13311 8631 13317
rect 8343 13280 8524 13308
rect 8343 13277 8355 13280
rect 8297 13271 8355 13277
rect 7926 13200 7932 13252
rect 7984 13240 7990 13252
rect 8312 13240 8340 13271
rect 7984 13212 8340 13240
rect 8389 13243 8447 13249
rect 7984 13200 7990 13212
rect 8389 13209 8401 13243
rect 8435 13209 8447 13243
rect 8496 13240 8524 13280
rect 8573 13277 8585 13311
rect 8619 13277 8631 13311
rect 8573 13271 8631 13277
rect 8846 13268 8852 13320
rect 8904 13308 8910 13320
rect 9125 13311 9183 13317
rect 9125 13308 9137 13311
rect 8904 13280 9137 13308
rect 8904 13268 8910 13280
rect 9125 13277 9137 13280
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 10686 13268 10692 13320
rect 10744 13317 10750 13320
rect 10888 13317 10916 13348
rect 11977 13345 11989 13348
rect 12023 13376 12035 13379
rect 12894 13376 12900 13388
rect 12023 13348 12900 13376
rect 12023 13345 12035 13348
rect 11977 13339 12035 13345
rect 12894 13336 12900 13348
rect 12952 13336 12958 13388
rect 13541 13379 13599 13385
rect 13541 13345 13553 13379
rect 13587 13376 13599 13379
rect 13814 13376 13820 13388
rect 13587 13348 13820 13376
rect 13587 13345 13599 13348
rect 13541 13339 13599 13345
rect 13814 13336 13820 13348
rect 13872 13376 13878 13388
rect 17126 13376 17132 13388
rect 13872 13348 17132 13376
rect 13872 13336 13878 13348
rect 17126 13336 17132 13348
rect 17184 13336 17190 13388
rect 17402 13336 17408 13388
rect 17460 13376 17466 13388
rect 17788 13376 17816 13416
rect 19518 13404 19524 13456
rect 19576 13404 19582 13456
rect 19610 13404 19616 13456
rect 19668 13444 19674 13456
rect 19668 13416 21220 13444
rect 19668 13404 19674 13416
rect 19334 13376 19340 13388
rect 17460 13348 17540 13376
rect 17788 13348 19340 13376
rect 17460 13336 17466 13348
rect 10744 13311 10777 13317
rect 10765 13277 10777 13311
rect 10744 13271 10777 13277
rect 10873 13311 10931 13317
rect 10873 13277 10885 13311
rect 10919 13277 10931 13311
rect 10873 13271 10931 13277
rect 10744 13268 10750 13271
rect 11330 13268 11336 13320
rect 11388 13268 11394 13320
rect 11609 13311 11667 13317
rect 11609 13277 11621 13311
rect 11655 13277 11667 13311
rect 11609 13271 11667 13277
rect 9953 13243 10011 13249
rect 9953 13240 9965 13243
rect 8496 13212 9965 13240
rect 8389 13203 8447 13209
rect 9953 13209 9965 13212
rect 9999 13240 10011 13243
rect 11054 13240 11060 13252
rect 9999 13212 11060 13240
rect 9999 13209 10011 13212
rect 9953 13203 10011 13209
rect 8404 13172 8432 13203
rect 11054 13200 11060 13212
rect 11112 13200 11118 13252
rect 11146 13200 11152 13252
rect 11204 13240 11210 13252
rect 11624 13240 11652 13271
rect 11698 13268 11704 13320
rect 11756 13308 11762 13320
rect 11793 13311 11851 13317
rect 11793 13308 11805 13311
rect 11756 13280 11805 13308
rect 11756 13268 11762 13280
rect 11793 13277 11805 13280
rect 11839 13308 11851 13311
rect 12158 13308 12164 13320
rect 11839 13280 12164 13308
rect 11839 13277 11851 13280
rect 11793 13271 11851 13277
rect 12158 13268 12164 13280
rect 12216 13268 12222 13320
rect 12526 13268 12532 13320
rect 12584 13268 12590 13320
rect 12805 13311 12863 13317
rect 12805 13277 12817 13311
rect 12851 13308 12863 13311
rect 13170 13308 13176 13320
rect 12851 13280 13176 13308
rect 12851 13277 12863 13280
rect 12805 13271 12863 13277
rect 13170 13268 13176 13280
rect 13228 13268 13234 13320
rect 13265 13311 13323 13317
rect 13265 13277 13277 13311
rect 13311 13277 13323 13311
rect 13265 13271 13323 13277
rect 11204 13212 11652 13240
rect 13280 13240 13308 13271
rect 13998 13268 14004 13320
rect 14056 13308 14062 13320
rect 14553 13311 14611 13317
rect 14553 13308 14565 13311
rect 14056 13280 14565 13308
rect 14056 13268 14062 13280
rect 14553 13277 14565 13280
rect 14599 13308 14611 13311
rect 15286 13308 15292 13320
rect 14599 13280 15292 13308
rect 14599 13277 14611 13280
rect 14553 13271 14611 13277
rect 15286 13268 15292 13280
rect 15344 13308 15350 13320
rect 15562 13308 15568 13320
rect 15344 13280 15568 13308
rect 15344 13268 15350 13280
rect 15562 13268 15568 13280
rect 15620 13268 15626 13320
rect 16390 13268 16396 13320
rect 16448 13268 16454 13320
rect 16485 13311 16543 13317
rect 16485 13277 16497 13311
rect 16531 13308 16543 13311
rect 16574 13308 16580 13320
rect 16531 13280 16580 13308
rect 16531 13277 16543 13280
rect 16485 13271 16543 13277
rect 16574 13268 16580 13280
rect 16632 13268 16638 13320
rect 16666 13268 16672 13320
rect 16724 13268 16730 13320
rect 13538 13240 13544 13252
rect 13280 13212 13544 13240
rect 11204 13200 11210 13212
rect 13538 13200 13544 13212
rect 13596 13200 13602 13252
rect 14277 13243 14335 13249
rect 14277 13209 14289 13243
rect 14323 13209 14335 13243
rect 14277 13203 14335 13209
rect 10042 13172 10048 13184
rect 6196 13144 10048 13172
rect 10042 13132 10048 13144
rect 10100 13132 10106 13184
rect 10502 13132 10508 13184
rect 10560 13132 10566 13184
rect 11330 13132 11336 13184
rect 11388 13172 11394 13184
rect 11974 13172 11980 13184
rect 11388 13144 11980 13172
rect 11388 13132 11394 13144
rect 11974 13132 11980 13144
rect 12032 13132 12038 13184
rect 14292 13172 14320 13203
rect 14458 13200 14464 13252
rect 14516 13200 14522 13252
rect 14568 13212 14872 13240
rect 14568 13172 14596 13212
rect 14844 13184 14872 13212
rect 14918 13200 14924 13252
rect 14976 13240 14982 13252
rect 16408 13240 16436 13268
rect 17402 13240 17408 13252
rect 14976 13212 16344 13240
rect 16408 13212 17408 13240
rect 14976 13200 14982 13212
rect 14292 13144 14596 13172
rect 14642 13132 14648 13184
rect 14700 13132 14706 13184
rect 14826 13132 14832 13184
rect 14884 13172 14890 13184
rect 15746 13172 15752 13184
rect 14884 13144 15752 13172
rect 14884 13132 14890 13144
rect 15746 13132 15752 13144
rect 15804 13172 15810 13184
rect 15933 13175 15991 13181
rect 15933 13172 15945 13175
rect 15804 13144 15945 13172
rect 15804 13132 15810 13144
rect 15933 13141 15945 13144
rect 15979 13172 15991 13175
rect 16206 13172 16212 13184
rect 15979 13144 16212 13172
rect 15979 13141 15991 13144
rect 15933 13135 15991 13141
rect 16206 13132 16212 13144
rect 16264 13132 16270 13184
rect 16316 13172 16344 13212
rect 17402 13200 17408 13212
rect 17460 13200 17466 13252
rect 17512 13240 17540 13348
rect 19334 13336 19340 13348
rect 19392 13376 19398 13388
rect 19536 13376 19564 13404
rect 19705 13379 19763 13385
rect 19392 13348 19656 13376
rect 19392 13336 19398 13348
rect 18782 13268 18788 13320
rect 18840 13308 18846 13320
rect 19628 13317 19656 13348
rect 19705 13345 19717 13379
rect 19751 13376 19763 13379
rect 20806 13376 20812 13388
rect 19751 13348 20812 13376
rect 19751 13345 19763 13348
rect 19705 13339 19763 13345
rect 20806 13336 20812 13348
rect 20864 13336 20870 13388
rect 21192 13385 21220 13416
rect 21177 13379 21235 13385
rect 21177 13345 21189 13379
rect 21223 13376 21235 13379
rect 21818 13376 21824 13388
rect 21223 13348 21824 13376
rect 21223 13345 21235 13348
rect 21177 13339 21235 13345
rect 21818 13336 21824 13348
rect 21876 13336 21882 13388
rect 19521 13311 19579 13317
rect 19521 13308 19533 13311
rect 18840 13280 19533 13308
rect 18840 13268 18846 13280
rect 19521 13277 19533 13280
rect 19567 13277 19579 13311
rect 19521 13271 19579 13277
rect 19613 13311 19671 13317
rect 19613 13277 19625 13311
rect 19659 13277 19671 13311
rect 19613 13271 19671 13277
rect 19797 13311 19855 13317
rect 19797 13277 19809 13311
rect 19843 13308 19855 13311
rect 20714 13308 20720 13320
rect 19843 13280 20720 13308
rect 19843 13277 19855 13280
rect 19797 13271 19855 13277
rect 20714 13268 20720 13280
rect 20772 13268 20778 13320
rect 20993 13311 21051 13317
rect 20993 13277 21005 13311
rect 21039 13308 21051 13311
rect 21913 13311 21971 13317
rect 21913 13308 21925 13311
rect 21039 13280 21925 13308
rect 21039 13277 21051 13280
rect 20993 13271 21051 13277
rect 21913 13277 21925 13280
rect 21959 13308 21971 13311
rect 22066 13308 22094 13484
rect 22922 13472 22928 13484
rect 22980 13472 22986 13524
rect 21959 13280 22094 13308
rect 22281 13311 22339 13317
rect 21959 13277 21971 13280
rect 21913 13271 21971 13277
rect 22281 13277 22293 13311
rect 22327 13308 22339 13311
rect 22830 13308 22836 13320
rect 22327 13280 22836 13308
rect 22327 13277 22339 13280
rect 22281 13271 22339 13277
rect 19242 13240 19248 13252
rect 17512 13212 19248 13240
rect 19242 13200 19248 13212
rect 19300 13240 19306 13252
rect 21008 13240 21036 13271
rect 22830 13268 22836 13280
rect 22888 13268 22894 13320
rect 19300 13212 21036 13240
rect 19300 13200 19306 13212
rect 20346 13172 20352 13184
rect 16316 13144 20352 13172
rect 20346 13132 20352 13144
rect 20404 13132 20410 13184
rect 1104 13082 23987 13104
rect 1104 13030 6630 13082
rect 6682 13030 6694 13082
rect 6746 13030 6758 13082
rect 6810 13030 6822 13082
rect 6874 13030 6886 13082
rect 6938 13030 12311 13082
rect 12363 13030 12375 13082
rect 12427 13030 12439 13082
rect 12491 13030 12503 13082
rect 12555 13030 12567 13082
rect 12619 13030 17992 13082
rect 18044 13030 18056 13082
rect 18108 13030 18120 13082
rect 18172 13030 18184 13082
rect 18236 13030 18248 13082
rect 18300 13030 23673 13082
rect 23725 13030 23737 13082
rect 23789 13030 23801 13082
rect 23853 13030 23865 13082
rect 23917 13030 23929 13082
rect 23981 13030 23987 13082
rect 1104 13008 23987 13030
rect 2590 12928 2596 12980
rect 2648 12968 2654 12980
rect 4341 12971 4399 12977
rect 4341 12968 4353 12971
rect 2648 12940 4353 12968
rect 2648 12928 2654 12940
rect 4341 12937 4353 12940
rect 4387 12937 4399 12971
rect 5369 12971 5427 12977
rect 5369 12968 5381 12971
rect 4341 12931 4399 12937
rect 4724 12940 5381 12968
rect 2406 12860 2412 12912
rect 2464 12900 2470 12912
rect 4724 12900 4752 12940
rect 5369 12937 5381 12940
rect 5415 12968 5427 12971
rect 6086 12968 6092 12980
rect 5415 12940 6092 12968
rect 5415 12937 5427 12940
rect 5369 12931 5427 12937
rect 6086 12928 6092 12940
rect 6144 12928 6150 12980
rect 10502 12928 10508 12980
rect 10560 12968 10566 12980
rect 12913 12971 12971 12977
rect 12913 12968 12925 12971
rect 10560 12940 12925 12968
rect 10560 12928 10566 12940
rect 12913 12937 12925 12940
rect 12959 12937 12971 12971
rect 12913 12931 12971 12937
rect 13170 12928 13176 12980
rect 13228 12968 13234 12980
rect 13541 12971 13599 12977
rect 13541 12968 13553 12971
rect 13228 12940 13553 12968
rect 13228 12928 13234 12940
rect 13541 12937 13553 12940
rect 13587 12937 13599 12971
rect 13541 12931 13599 12937
rect 13906 12928 13912 12980
rect 13964 12928 13970 12980
rect 14366 12928 14372 12980
rect 14424 12968 14430 12980
rect 14737 12971 14795 12977
rect 14737 12968 14749 12971
rect 14424 12940 14749 12968
rect 14424 12928 14430 12940
rect 14737 12937 14749 12940
rect 14783 12937 14795 12971
rect 14737 12931 14795 12937
rect 17126 12928 17132 12980
rect 17184 12968 17190 12980
rect 17586 12968 17592 12980
rect 17184 12940 17592 12968
rect 17184 12928 17190 12940
rect 17586 12928 17592 12940
rect 17644 12928 17650 12980
rect 18325 12971 18383 12977
rect 18325 12937 18337 12971
rect 18371 12968 18383 12971
rect 18506 12968 18512 12980
rect 18371 12940 18512 12968
rect 18371 12937 18383 12940
rect 18325 12931 18383 12937
rect 18506 12928 18512 12940
rect 18564 12928 18570 12980
rect 20070 12928 20076 12980
rect 20128 12968 20134 12980
rect 22005 12971 22063 12977
rect 22005 12968 22017 12971
rect 20128 12940 22017 12968
rect 20128 12928 20134 12940
rect 22005 12937 22017 12940
rect 22051 12937 22063 12971
rect 22005 12931 22063 12937
rect 2464 12872 4752 12900
rect 2464 12860 2470 12872
rect 5166 12860 5172 12912
rect 5224 12860 5230 12912
rect 6914 12860 6920 12912
rect 6972 12900 6978 12912
rect 7009 12903 7067 12909
rect 7009 12900 7021 12903
rect 6972 12872 7021 12900
rect 6972 12860 6978 12872
rect 7009 12869 7021 12872
rect 7055 12900 7067 12903
rect 7098 12900 7104 12912
rect 7055 12872 7104 12900
rect 7055 12869 7067 12872
rect 7009 12863 7067 12869
rect 7098 12860 7104 12872
rect 7156 12860 7162 12912
rect 8846 12860 8852 12912
rect 8904 12900 8910 12912
rect 8904 12872 10456 12900
rect 8904 12860 8910 12872
rect 2225 12835 2283 12841
rect 2225 12801 2237 12835
rect 2271 12801 2283 12835
rect 2225 12795 2283 12801
rect 2240 12764 2268 12795
rect 2682 12792 2688 12844
rect 2740 12832 2746 12844
rect 2777 12835 2835 12841
rect 2777 12832 2789 12835
rect 2740 12804 2789 12832
rect 2740 12792 2746 12804
rect 2777 12801 2789 12804
rect 2823 12801 2835 12835
rect 2777 12795 2835 12801
rect 2958 12792 2964 12844
rect 3016 12792 3022 12844
rect 3053 12835 3111 12841
rect 3053 12801 3065 12835
rect 3099 12832 3111 12835
rect 3234 12832 3240 12844
rect 3099 12804 3240 12832
rect 3099 12801 3111 12804
rect 3053 12795 3111 12801
rect 3234 12792 3240 12804
rect 3292 12792 3298 12844
rect 3418 12792 3424 12844
rect 3476 12832 3482 12844
rect 4525 12835 4583 12841
rect 4525 12832 4537 12835
rect 3476 12804 4537 12832
rect 3476 12792 3482 12804
rect 4525 12801 4537 12804
rect 4571 12801 4583 12835
rect 4525 12795 4583 12801
rect 4709 12835 4767 12841
rect 4709 12801 4721 12835
rect 4755 12832 4767 12835
rect 5534 12832 5540 12844
rect 4755 12804 5540 12832
rect 4755 12801 4767 12804
rect 4709 12795 4767 12801
rect 5534 12792 5540 12804
rect 5592 12792 5598 12844
rect 6086 12792 6092 12844
rect 6144 12832 6150 12844
rect 6454 12832 6460 12844
rect 6144 12804 6460 12832
rect 6144 12792 6150 12804
rect 6454 12792 6460 12804
rect 6512 12832 6518 12844
rect 6733 12835 6791 12841
rect 6733 12832 6745 12835
rect 6512 12804 6745 12832
rect 6512 12792 6518 12804
rect 6733 12801 6745 12804
rect 6779 12801 6791 12835
rect 6733 12795 6791 12801
rect 6825 12835 6883 12841
rect 6825 12801 6837 12835
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 3142 12764 3148 12776
rect 2240 12736 3148 12764
rect 3142 12724 3148 12736
rect 3200 12724 3206 12776
rect 5442 12724 5448 12776
rect 5500 12764 5506 12776
rect 6840 12764 6868 12795
rect 9030 12792 9036 12844
rect 9088 12792 9094 12844
rect 9214 12792 9220 12844
rect 9272 12792 9278 12844
rect 9950 12792 9956 12844
rect 10008 12832 10014 12844
rect 10137 12835 10195 12841
rect 10137 12832 10149 12835
rect 10008 12804 10149 12832
rect 10008 12792 10014 12804
rect 10137 12801 10149 12804
rect 10183 12801 10195 12835
rect 10137 12795 10195 12801
rect 10226 12792 10232 12844
rect 10284 12792 10290 12844
rect 10428 12841 10456 12872
rect 10686 12860 10692 12912
rect 10744 12860 10750 12912
rect 11698 12860 11704 12912
rect 11756 12860 11762 12912
rect 12710 12860 12716 12912
rect 12768 12860 12774 12912
rect 13722 12860 13728 12912
rect 13780 12900 13786 12912
rect 14001 12903 14059 12909
rect 14001 12900 14013 12903
rect 13780 12872 14013 12900
rect 13780 12860 13786 12872
rect 14001 12869 14013 12872
rect 14047 12900 14059 12903
rect 15378 12900 15384 12912
rect 14047 12872 14136 12900
rect 14047 12869 14059 12872
rect 14001 12863 14059 12869
rect 10413 12835 10471 12841
rect 10413 12801 10425 12835
rect 10459 12801 10471 12835
rect 10704 12832 10732 12860
rect 11885 12835 11943 12841
rect 11885 12832 11897 12835
rect 10704 12804 11897 12832
rect 10413 12795 10471 12801
rect 11885 12801 11897 12804
rect 11931 12801 11943 12835
rect 11885 12795 11943 12801
rect 11974 12792 11980 12844
rect 12032 12792 12038 12844
rect 13814 12792 13820 12844
rect 13872 12792 13878 12844
rect 5500 12736 6868 12764
rect 5500 12724 5506 12736
rect 6472 12708 6500 12736
rect 10686 12724 10692 12776
rect 10744 12764 10750 12776
rect 10873 12767 10931 12773
rect 10873 12764 10885 12767
rect 10744 12736 10885 12764
rect 10744 12724 10750 12736
rect 10873 12733 10885 12736
rect 10919 12733 10931 12767
rect 14108 12764 14136 12872
rect 14292 12872 15384 12900
rect 14182 12792 14188 12844
rect 14240 12792 14246 12844
rect 14292 12841 14320 12872
rect 15378 12860 15384 12872
rect 15436 12860 15442 12912
rect 15470 12860 15476 12912
rect 15528 12860 15534 12912
rect 15703 12869 15761 12875
rect 15703 12866 15715 12869
rect 14277 12835 14335 12841
rect 14277 12801 14289 12835
rect 14323 12801 14335 12835
rect 14277 12795 14335 12801
rect 14737 12835 14795 12841
rect 14737 12801 14749 12835
rect 14783 12832 14795 12835
rect 14826 12832 14832 12844
rect 14783 12804 14832 12832
rect 14783 12801 14795 12804
rect 14737 12795 14795 12801
rect 14826 12792 14832 12804
rect 14884 12792 14890 12844
rect 14921 12835 14979 12841
rect 14921 12801 14933 12835
rect 14967 12801 14979 12835
rect 14921 12795 14979 12801
rect 14458 12764 14464 12776
rect 14108 12736 14464 12764
rect 10873 12727 10931 12733
rect 14458 12724 14464 12736
rect 14516 12724 14522 12776
rect 14936 12764 14964 12795
rect 15286 12792 15292 12844
rect 15344 12832 15350 12844
rect 15688 12835 15715 12866
rect 15749 12844 15761 12869
rect 16022 12860 16028 12912
rect 16080 12900 16086 12912
rect 16298 12900 16304 12912
rect 16080 12872 16304 12900
rect 16080 12860 16086 12872
rect 16298 12860 16304 12872
rect 16356 12900 16362 12912
rect 16356 12872 21680 12900
rect 16356 12860 16362 12872
rect 15749 12835 15752 12844
rect 15688 12832 15752 12835
rect 15344 12804 15752 12832
rect 15344 12792 15350 12804
rect 15746 12792 15752 12804
rect 15804 12792 15810 12844
rect 16868 12841 16896 12872
rect 21652 12844 21680 12872
rect 21818 12860 21824 12912
rect 21876 12900 21882 12912
rect 22373 12903 22431 12909
rect 22373 12900 22385 12903
rect 21876 12872 22385 12900
rect 21876 12860 21882 12872
rect 22373 12869 22385 12872
rect 22419 12869 22431 12903
rect 22373 12863 22431 12869
rect 16853 12835 16911 12841
rect 16853 12801 16865 12835
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 16942 12792 16948 12844
rect 17000 12832 17006 12844
rect 17000 12804 17045 12832
rect 17000 12792 17006 12804
rect 17126 12792 17132 12844
rect 17184 12792 17190 12844
rect 17218 12792 17224 12844
rect 17276 12792 17282 12844
rect 17402 12841 17408 12844
rect 17359 12835 17408 12841
rect 17359 12801 17371 12835
rect 17405 12801 17408 12835
rect 17359 12795 17408 12801
rect 17402 12792 17408 12795
rect 17460 12792 17466 12844
rect 18601 12835 18659 12841
rect 18601 12801 18613 12835
rect 18647 12832 18659 12835
rect 19058 12832 19064 12844
rect 18647 12804 19064 12832
rect 18647 12801 18659 12804
rect 18601 12795 18659 12801
rect 19058 12792 19064 12804
rect 19116 12792 19122 12844
rect 21634 12792 21640 12844
rect 21692 12832 21698 12844
rect 22094 12832 22100 12844
rect 21692 12804 22100 12832
rect 21692 12792 21698 12804
rect 22094 12792 22100 12804
rect 22152 12832 22158 12844
rect 22189 12835 22247 12841
rect 22189 12832 22201 12835
rect 22152 12804 22201 12832
rect 22152 12792 22158 12804
rect 22189 12801 22201 12804
rect 22235 12801 22247 12835
rect 22189 12795 22247 12801
rect 22462 12792 22468 12844
rect 22520 12792 22526 12844
rect 18230 12764 18236 12776
rect 14936 12736 18236 12764
rect 18230 12724 18236 12736
rect 18288 12724 18294 12776
rect 18506 12724 18512 12776
rect 18564 12724 18570 12776
rect 18693 12767 18751 12773
rect 18693 12764 18705 12767
rect 18616 12736 18705 12764
rect 18616 12708 18644 12736
rect 18693 12733 18705 12736
rect 18739 12733 18751 12767
rect 18693 12727 18751 12733
rect 18782 12724 18788 12776
rect 18840 12724 18846 12776
rect 2774 12656 2780 12708
rect 2832 12656 2838 12708
rect 3050 12656 3056 12708
rect 3108 12696 3114 12708
rect 3418 12696 3424 12708
rect 3108 12668 3424 12696
rect 3108 12656 3114 12668
rect 3418 12656 3424 12668
rect 3476 12696 3482 12708
rect 5537 12699 5595 12705
rect 3476 12668 5396 12696
rect 3476 12656 3482 12668
rect 2038 12588 2044 12640
rect 2096 12628 2102 12640
rect 2133 12631 2191 12637
rect 2133 12628 2145 12631
rect 2096 12600 2145 12628
rect 2096 12588 2102 12600
rect 2133 12597 2145 12600
rect 2179 12628 2191 12631
rect 2498 12628 2504 12640
rect 2179 12600 2504 12628
rect 2179 12597 2191 12600
rect 2133 12591 2191 12597
rect 2498 12588 2504 12600
rect 2556 12588 2562 12640
rect 2590 12588 2596 12640
rect 2648 12628 2654 12640
rect 2958 12628 2964 12640
rect 2648 12600 2964 12628
rect 2648 12588 2654 12600
rect 2958 12588 2964 12600
rect 3016 12628 3022 12640
rect 5258 12628 5264 12640
rect 3016 12600 5264 12628
rect 3016 12588 3022 12600
rect 5258 12588 5264 12600
rect 5316 12588 5322 12640
rect 5368 12637 5396 12668
rect 5537 12665 5549 12699
rect 5583 12696 5595 12699
rect 5994 12696 6000 12708
rect 5583 12668 6000 12696
rect 5583 12665 5595 12668
rect 5537 12659 5595 12665
rect 5994 12656 6000 12668
rect 6052 12656 6058 12708
rect 6454 12656 6460 12708
rect 6512 12656 6518 12708
rect 7009 12699 7067 12705
rect 7009 12665 7021 12699
rect 7055 12696 7067 12699
rect 8018 12696 8024 12708
rect 7055 12668 8024 12696
rect 7055 12665 7067 12668
rect 7009 12659 7067 12665
rect 8018 12656 8024 12668
rect 8076 12656 8082 12708
rect 11882 12656 11888 12708
rect 11940 12696 11946 12708
rect 12161 12699 12219 12705
rect 12161 12696 12173 12699
rect 11940 12668 12173 12696
rect 11940 12656 11946 12668
rect 12161 12665 12173 12668
rect 12207 12696 12219 12699
rect 13081 12699 13139 12705
rect 12207 12668 12434 12696
rect 12207 12665 12219 12668
rect 12161 12659 12219 12665
rect 5353 12631 5411 12637
rect 5353 12597 5365 12631
rect 5399 12597 5411 12631
rect 5353 12591 5411 12597
rect 9306 12588 9312 12640
rect 9364 12588 9370 12640
rect 11146 12588 11152 12640
rect 11204 12628 11210 12640
rect 11701 12631 11759 12637
rect 11701 12628 11713 12631
rect 11204 12600 11713 12628
rect 11204 12588 11210 12600
rect 11701 12597 11713 12600
rect 11747 12597 11759 12631
rect 12406 12628 12434 12668
rect 13081 12665 13093 12699
rect 13127 12696 13139 12699
rect 13446 12696 13452 12708
rect 13127 12668 13452 12696
rect 13127 12665 13139 12668
rect 13081 12659 13139 12665
rect 13446 12656 13452 12668
rect 13504 12656 13510 12708
rect 17034 12696 17040 12708
rect 15672 12668 17040 12696
rect 12897 12631 12955 12637
rect 12897 12628 12909 12631
rect 12406 12600 12909 12628
rect 11701 12591 11759 12597
rect 12897 12597 12909 12600
rect 12943 12597 12955 12631
rect 12897 12591 12955 12597
rect 13262 12588 13268 12640
rect 13320 12628 13326 12640
rect 15470 12628 15476 12640
rect 13320 12600 15476 12628
rect 13320 12588 13326 12600
rect 15470 12588 15476 12600
rect 15528 12588 15534 12640
rect 15672 12637 15700 12668
rect 17034 12656 17040 12668
rect 17092 12656 17098 12708
rect 18598 12656 18604 12708
rect 18656 12696 18662 12708
rect 19150 12696 19156 12708
rect 18656 12668 19156 12696
rect 18656 12656 18662 12668
rect 19150 12656 19156 12668
rect 19208 12696 19214 12708
rect 19337 12699 19395 12705
rect 19337 12696 19349 12699
rect 19208 12668 19349 12696
rect 19208 12656 19214 12668
rect 19337 12665 19349 12668
rect 19383 12665 19395 12699
rect 19337 12659 19395 12665
rect 15657 12631 15715 12637
rect 15657 12597 15669 12631
rect 15703 12597 15715 12631
rect 15657 12591 15715 12597
rect 15841 12631 15899 12637
rect 15841 12597 15853 12631
rect 15887 12628 15899 12631
rect 16574 12628 16580 12640
rect 15887 12600 16580 12628
rect 15887 12597 15899 12600
rect 15841 12591 15899 12597
rect 16574 12588 16580 12600
rect 16632 12588 16638 12640
rect 17497 12631 17555 12637
rect 17497 12597 17509 12631
rect 17543 12628 17555 12631
rect 17862 12628 17868 12640
rect 17543 12600 17868 12628
rect 17543 12597 17555 12600
rect 17497 12591 17555 12597
rect 17862 12588 17868 12600
rect 17920 12588 17926 12640
rect 20346 12588 20352 12640
rect 20404 12628 20410 12640
rect 22922 12628 22928 12640
rect 20404 12600 22928 12628
rect 20404 12588 20410 12600
rect 22922 12588 22928 12600
rect 22980 12588 22986 12640
rect 1104 12538 23828 12560
rect 1104 12486 3790 12538
rect 3842 12486 3854 12538
rect 3906 12486 3918 12538
rect 3970 12486 3982 12538
rect 4034 12486 4046 12538
rect 4098 12486 9471 12538
rect 9523 12486 9535 12538
rect 9587 12486 9599 12538
rect 9651 12486 9663 12538
rect 9715 12486 9727 12538
rect 9779 12486 15152 12538
rect 15204 12486 15216 12538
rect 15268 12486 15280 12538
rect 15332 12486 15344 12538
rect 15396 12486 15408 12538
rect 15460 12486 20833 12538
rect 20885 12486 20897 12538
rect 20949 12486 20961 12538
rect 21013 12486 21025 12538
rect 21077 12486 21089 12538
rect 21141 12486 23828 12538
rect 1104 12464 23828 12486
rect 1762 12384 1768 12436
rect 1820 12384 1826 12436
rect 1857 12427 1915 12433
rect 1857 12393 1869 12427
rect 1903 12424 1915 12427
rect 1946 12424 1952 12436
rect 1903 12396 1952 12424
rect 1903 12393 1915 12396
rect 1857 12387 1915 12393
rect 1946 12384 1952 12396
rect 2004 12384 2010 12436
rect 2406 12384 2412 12436
rect 2464 12384 2470 12436
rect 2590 12384 2596 12436
rect 2648 12384 2654 12436
rect 4798 12384 4804 12436
rect 4856 12424 4862 12436
rect 5258 12424 5264 12436
rect 4856 12396 5264 12424
rect 4856 12384 4862 12396
rect 5258 12384 5264 12396
rect 5316 12384 5322 12436
rect 5626 12384 5632 12436
rect 5684 12424 5690 12436
rect 7282 12424 7288 12436
rect 5684 12396 7288 12424
rect 5684 12384 5690 12396
rect 7282 12384 7288 12396
rect 7340 12384 7346 12436
rect 7558 12384 7564 12436
rect 7616 12384 7622 12436
rect 8110 12384 8116 12436
rect 8168 12384 8174 12436
rect 13633 12427 13691 12433
rect 13633 12393 13645 12427
rect 13679 12424 13691 12427
rect 14642 12424 14648 12436
rect 13679 12396 14648 12424
rect 13679 12393 13691 12396
rect 13633 12387 13691 12393
rect 14642 12384 14648 12396
rect 14700 12384 14706 12436
rect 16942 12424 16948 12436
rect 14844 12396 16948 12424
rect 4433 12359 4491 12365
rect 4433 12325 4445 12359
rect 4479 12356 4491 12359
rect 7006 12356 7012 12368
rect 4479 12328 7012 12356
rect 4479 12325 4491 12328
rect 4433 12319 4491 12325
rect 7006 12316 7012 12328
rect 7064 12316 7070 12368
rect 8202 12316 8208 12368
rect 8260 12356 8266 12368
rect 9214 12356 9220 12368
rect 8260 12328 9220 12356
rect 8260 12316 8266 12328
rect 1946 12248 1952 12300
rect 2004 12288 2010 12300
rect 2130 12288 2136 12300
rect 2004 12260 2136 12288
rect 2004 12248 2010 12260
rect 2130 12248 2136 12260
rect 2188 12248 2194 12300
rect 4522 12248 4528 12300
rect 4580 12288 4586 12300
rect 4580 12260 8340 12288
rect 4580 12248 4586 12260
rect 1673 12223 1731 12229
rect 1673 12189 1685 12223
rect 1719 12189 1731 12223
rect 1673 12183 1731 12189
rect 1688 12084 1716 12183
rect 3694 12180 3700 12232
rect 3752 12220 3758 12232
rect 4065 12223 4123 12229
rect 4065 12220 4077 12223
rect 3752 12192 4077 12220
rect 3752 12180 3758 12192
rect 4065 12189 4077 12192
rect 4111 12189 4123 12223
rect 4065 12183 4123 12189
rect 4219 12223 4277 12229
rect 4219 12189 4231 12223
rect 4265 12220 4277 12223
rect 4430 12220 4436 12232
rect 4265 12192 4436 12220
rect 4265 12189 4277 12192
rect 4219 12183 4277 12189
rect 4430 12180 4436 12192
rect 4488 12180 4494 12232
rect 6914 12180 6920 12232
rect 6972 12220 6978 12232
rect 7374 12220 7380 12232
rect 6972 12192 7380 12220
rect 6972 12180 6978 12192
rect 7374 12180 7380 12192
rect 7432 12180 7438 12232
rect 7558 12180 7564 12232
rect 7616 12220 7622 12232
rect 7926 12220 7932 12232
rect 7616 12192 7932 12220
rect 7616 12180 7622 12192
rect 7926 12180 7932 12192
rect 7984 12180 7990 12232
rect 8312 12229 8340 12260
rect 8021 12223 8079 12229
rect 8021 12189 8033 12223
rect 8067 12189 8079 12223
rect 8021 12183 8079 12189
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12189 8355 12223
rect 8297 12183 8355 12189
rect 2774 12112 2780 12164
rect 2832 12152 2838 12164
rect 2958 12152 2964 12164
rect 2832 12124 2964 12152
rect 2832 12112 2838 12124
rect 2958 12112 2964 12124
rect 3016 12112 3022 12164
rect 7098 12152 7104 12164
rect 7024 12124 7104 12152
rect 2567 12087 2625 12093
rect 2567 12084 2579 12087
rect 1688 12056 2579 12084
rect 2567 12053 2579 12056
rect 2613 12084 2625 12087
rect 3234 12084 3240 12096
rect 2613 12056 3240 12084
rect 2613 12053 2625 12056
rect 2567 12047 2625 12053
rect 3234 12044 3240 12056
rect 3292 12044 3298 12096
rect 3786 12044 3792 12096
rect 3844 12084 3850 12096
rect 4893 12087 4951 12093
rect 4893 12084 4905 12087
rect 3844 12056 4905 12084
rect 3844 12044 3850 12056
rect 4893 12053 4905 12056
rect 4939 12053 4951 12087
rect 4893 12047 4951 12053
rect 5442 12044 5448 12096
rect 5500 12084 5506 12096
rect 6365 12087 6423 12093
rect 6365 12084 6377 12087
rect 5500 12056 6377 12084
rect 5500 12044 5506 12056
rect 6365 12053 6377 12056
rect 6411 12084 6423 12087
rect 7024 12084 7052 12124
rect 7098 12112 7104 12124
rect 7156 12112 7162 12164
rect 8036 12152 8064 12183
rect 8386 12180 8392 12232
rect 8444 12180 8450 12232
rect 9140 12229 9168 12328
rect 9214 12316 9220 12328
rect 9272 12316 9278 12368
rect 10318 12316 10324 12368
rect 10376 12356 10382 12368
rect 13814 12356 13820 12368
rect 10376 12328 13820 12356
rect 10376 12316 10382 12328
rect 13814 12316 13820 12328
rect 13872 12316 13878 12368
rect 11606 12248 11612 12300
rect 11664 12288 11670 12300
rect 11885 12291 11943 12297
rect 11885 12288 11897 12291
rect 11664 12260 11897 12288
rect 11664 12248 11670 12260
rect 11885 12257 11897 12260
rect 11931 12257 11943 12291
rect 11885 12251 11943 12257
rect 12986 12248 12992 12300
rect 13044 12288 13050 12300
rect 14550 12288 14556 12300
rect 13044 12260 13308 12288
rect 13044 12248 13050 12260
rect 13280 12232 13308 12260
rect 13740 12260 14556 12288
rect 13740 12232 13768 12260
rect 14550 12248 14556 12260
rect 14608 12248 14614 12300
rect 14844 12297 14872 12396
rect 16942 12384 16948 12396
rect 17000 12424 17006 12436
rect 17494 12424 17500 12436
rect 17000 12396 17500 12424
rect 17000 12384 17006 12396
rect 17494 12384 17500 12396
rect 17552 12384 17558 12436
rect 18141 12427 18199 12433
rect 18141 12393 18153 12427
rect 18187 12424 18199 12427
rect 18322 12424 18328 12436
rect 18187 12396 18328 12424
rect 18187 12393 18199 12396
rect 18141 12387 18199 12393
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 19334 12384 19340 12436
rect 19392 12424 19398 12436
rect 19518 12424 19524 12436
rect 19392 12396 19524 12424
rect 19392 12384 19398 12396
rect 19518 12384 19524 12396
rect 19576 12384 19582 12436
rect 19702 12384 19708 12436
rect 19760 12384 19766 12436
rect 21818 12424 21824 12436
rect 21560 12396 21824 12424
rect 21560 12368 21588 12396
rect 21818 12384 21824 12396
rect 21876 12384 21882 12436
rect 15194 12316 15200 12368
rect 15252 12356 15258 12368
rect 15562 12356 15568 12368
rect 15252 12328 15568 12356
rect 15252 12316 15258 12328
rect 15562 12316 15568 12328
rect 15620 12316 15626 12368
rect 15838 12356 15844 12368
rect 15764 12328 15844 12356
rect 14829 12291 14887 12297
rect 14829 12257 14841 12291
rect 14875 12257 14887 12291
rect 14829 12251 14887 12257
rect 14918 12248 14924 12300
rect 14976 12288 14982 12300
rect 15764 12297 15792 12328
rect 15838 12316 15844 12328
rect 15896 12316 15902 12368
rect 16025 12359 16083 12365
rect 16025 12325 16037 12359
rect 16071 12356 16083 12359
rect 16666 12356 16672 12368
rect 16071 12328 16672 12356
rect 16071 12325 16083 12328
rect 16025 12319 16083 12325
rect 16666 12316 16672 12328
rect 16724 12356 16730 12368
rect 16724 12328 16896 12356
rect 16724 12316 16730 12328
rect 15749 12291 15807 12297
rect 15749 12288 15761 12291
rect 14976 12260 15761 12288
rect 14976 12248 14982 12260
rect 15749 12257 15761 12260
rect 15795 12257 15807 12291
rect 15749 12251 15807 12257
rect 16574 12248 16580 12300
rect 16632 12288 16638 12300
rect 16632 12260 16804 12288
rect 16632 12248 16638 12260
rect 9125 12223 9183 12229
rect 9125 12189 9137 12223
rect 9171 12189 9183 12223
rect 9125 12183 9183 12189
rect 9582 12180 9588 12232
rect 9640 12220 9646 12232
rect 9677 12223 9735 12229
rect 9677 12220 9689 12223
rect 9640 12192 9689 12220
rect 9640 12180 9646 12192
rect 9677 12189 9689 12192
rect 9723 12189 9735 12223
rect 9677 12183 9735 12189
rect 9858 12180 9864 12232
rect 9916 12220 9922 12232
rect 11977 12223 12035 12229
rect 11977 12220 11989 12223
rect 9916 12192 11989 12220
rect 9916 12180 9922 12192
rect 11977 12189 11989 12192
rect 12023 12189 12035 12223
rect 11977 12183 12035 12189
rect 12066 12180 12072 12232
rect 12124 12220 12130 12232
rect 12161 12223 12219 12229
rect 12161 12220 12173 12223
rect 12124 12192 12173 12220
rect 12124 12180 12130 12192
rect 12161 12189 12173 12192
rect 12207 12189 12219 12223
rect 12161 12183 12219 12189
rect 12710 12180 12716 12232
rect 12768 12220 12774 12232
rect 13081 12223 13139 12229
rect 13081 12220 13093 12223
rect 12768 12192 13093 12220
rect 12768 12180 12774 12192
rect 13081 12189 13093 12192
rect 13127 12220 13139 12223
rect 13127 12192 13216 12220
rect 13127 12189 13139 12192
rect 13081 12183 13139 12189
rect 8478 12152 8484 12164
rect 8036 12124 8484 12152
rect 8478 12112 8484 12124
rect 8536 12112 8542 12164
rect 10226 12112 10232 12164
rect 10284 12152 10290 12164
rect 10689 12155 10747 12161
rect 10689 12152 10701 12155
rect 10284 12124 10701 12152
rect 10284 12112 10290 12124
rect 10689 12121 10701 12124
rect 10735 12121 10747 12155
rect 10689 12115 10747 12121
rect 10873 12155 10931 12161
rect 10873 12121 10885 12155
rect 10919 12152 10931 12155
rect 11882 12152 11888 12164
rect 10919 12124 11888 12152
rect 10919 12121 10931 12124
rect 10873 12115 10931 12121
rect 11882 12112 11888 12124
rect 11940 12112 11946 12164
rect 12621 12155 12679 12161
rect 12621 12121 12633 12155
rect 12667 12152 12679 12155
rect 12986 12152 12992 12164
rect 12667 12124 12992 12152
rect 12667 12121 12679 12124
rect 12621 12115 12679 12121
rect 12986 12112 12992 12124
rect 13044 12112 13050 12164
rect 6411 12056 7052 12084
rect 6411 12053 6423 12056
rect 6365 12047 6423 12053
rect 8570 12044 8576 12096
rect 8628 12044 8634 12096
rect 9214 12044 9220 12096
rect 9272 12044 9278 12096
rect 10502 12044 10508 12096
rect 10560 12044 10566 12096
rect 13188 12084 13216 12192
rect 13262 12180 13268 12232
rect 13320 12180 13326 12232
rect 13449 12223 13507 12229
rect 13449 12189 13461 12223
rect 13495 12220 13507 12223
rect 13722 12220 13728 12232
rect 13495 12192 13728 12220
rect 13495 12189 13507 12192
rect 13449 12183 13507 12189
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 14277 12223 14335 12229
rect 14277 12189 14289 12223
rect 14323 12220 14335 12223
rect 14366 12220 14372 12232
rect 14323 12192 14372 12220
rect 14323 12189 14335 12192
rect 14277 12183 14335 12189
rect 14366 12180 14372 12192
rect 14424 12180 14430 12232
rect 14458 12180 14464 12232
rect 14516 12180 14522 12232
rect 15562 12180 15568 12232
rect 15620 12180 15626 12232
rect 15654 12180 15660 12232
rect 15712 12180 15718 12232
rect 15838 12180 15844 12232
rect 15896 12220 15902 12232
rect 15896 12192 16436 12220
rect 15896 12180 15902 12192
rect 13357 12155 13415 12161
rect 13357 12121 13369 12155
rect 13403 12152 13415 12155
rect 13538 12152 13544 12164
rect 13403 12124 13544 12152
rect 13403 12121 13415 12124
rect 13357 12115 13415 12121
rect 13538 12112 13544 12124
rect 13596 12112 13602 12164
rect 15580 12152 15608 12180
rect 16022 12152 16028 12164
rect 15580 12124 16028 12152
rect 16022 12112 16028 12124
rect 16080 12112 16086 12164
rect 16408 12152 16436 12192
rect 16482 12180 16488 12232
rect 16540 12180 16546 12232
rect 16666 12180 16672 12232
rect 16724 12180 16730 12232
rect 16776 12229 16804 12260
rect 16868 12229 16896 12328
rect 17034 12316 17040 12368
rect 17092 12356 17098 12368
rect 19610 12356 19616 12368
rect 17092 12328 19616 12356
rect 17092 12316 17098 12328
rect 19610 12316 19616 12328
rect 19668 12316 19674 12368
rect 19720 12328 21220 12356
rect 17129 12291 17187 12297
rect 17129 12257 17141 12291
rect 17175 12288 17187 12291
rect 17681 12291 17739 12297
rect 17681 12288 17693 12291
rect 17175 12260 17693 12288
rect 17175 12257 17187 12260
rect 17129 12251 17187 12257
rect 17681 12257 17693 12260
rect 17727 12257 17739 12291
rect 17681 12251 17739 12257
rect 17770 12248 17776 12300
rect 17828 12248 17834 12300
rect 17862 12248 17868 12300
rect 17920 12248 17926 12300
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 19720 12288 19748 12328
rect 19392 12260 19748 12288
rect 19392 12248 19398 12260
rect 19794 12248 19800 12300
rect 19852 12288 19858 12300
rect 19852 12260 20208 12288
rect 19852 12248 19858 12260
rect 16761 12223 16819 12229
rect 16761 12189 16773 12223
rect 16807 12189 16819 12223
rect 16761 12183 16819 12189
rect 16853 12223 16911 12229
rect 16853 12189 16865 12223
rect 16899 12189 16911 12223
rect 16853 12183 16911 12189
rect 17402 12180 17408 12232
rect 17460 12220 17466 12232
rect 17957 12223 18015 12229
rect 17957 12220 17969 12223
rect 17460 12192 17969 12220
rect 17460 12180 17466 12192
rect 17957 12189 17969 12192
rect 18003 12189 18015 12223
rect 17957 12183 18015 12189
rect 19889 12223 19947 12229
rect 19889 12189 19901 12223
rect 19935 12189 19947 12223
rect 19889 12183 19947 12189
rect 19981 12223 20039 12229
rect 19981 12189 19993 12223
rect 20027 12189 20039 12223
rect 19981 12183 20039 12189
rect 19058 12152 19064 12164
rect 16408 12124 19064 12152
rect 19058 12112 19064 12124
rect 19116 12112 19122 12164
rect 14274 12084 14280 12096
rect 13188 12056 14280 12084
rect 14274 12044 14280 12056
rect 14332 12044 14338 12096
rect 17310 12044 17316 12096
rect 17368 12084 17374 12096
rect 17770 12084 17776 12096
rect 17368 12056 17776 12084
rect 17368 12044 17374 12056
rect 17770 12044 17776 12056
rect 17828 12084 17834 12096
rect 19904 12084 19932 12183
rect 19996 12152 20024 12183
rect 20070 12180 20076 12232
rect 20128 12180 20134 12232
rect 20180 12229 20208 12260
rect 21082 12248 21088 12300
rect 21140 12248 21146 12300
rect 21192 12288 21220 12328
rect 21266 12316 21272 12368
rect 21324 12356 21330 12368
rect 21450 12356 21456 12368
rect 21324 12328 21456 12356
rect 21324 12316 21330 12328
rect 21450 12316 21456 12328
rect 21508 12316 21514 12368
rect 21542 12316 21548 12368
rect 21600 12316 21606 12368
rect 22462 12356 22468 12368
rect 21744 12328 22468 12356
rect 21744 12297 21772 12328
rect 22462 12316 22468 12328
rect 22520 12316 22526 12368
rect 21729 12291 21787 12297
rect 21192 12260 21588 12288
rect 20165 12223 20223 12229
rect 20165 12189 20177 12223
rect 20211 12189 20223 12223
rect 20165 12183 20223 12189
rect 20346 12180 20352 12232
rect 20404 12180 20410 12232
rect 20714 12180 20720 12232
rect 20772 12220 20778 12232
rect 21174 12220 21180 12232
rect 20772 12192 21180 12220
rect 20772 12180 20778 12192
rect 21174 12180 21180 12192
rect 21232 12220 21238 12232
rect 21269 12223 21327 12229
rect 21269 12220 21281 12223
rect 21232 12192 21281 12220
rect 21232 12180 21238 12192
rect 21269 12189 21281 12192
rect 21315 12189 21327 12223
rect 21269 12183 21327 12189
rect 21450 12180 21456 12232
rect 21508 12180 21514 12232
rect 21560 12229 21588 12260
rect 21729 12257 21741 12291
rect 21775 12257 21787 12291
rect 21729 12251 21787 12257
rect 21910 12248 21916 12300
rect 21968 12288 21974 12300
rect 22922 12288 22928 12300
rect 21968 12260 22094 12288
rect 21968 12248 21974 12260
rect 21560 12223 21629 12229
rect 21560 12192 21583 12223
rect 21571 12189 21583 12192
rect 21617 12189 21629 12223
rect 22066 12220 22094 12260
rect 22296 12260 22928 12288
rect 22296 12229 22324 12260
rect 22922 12248 22928 12260
rect 22980 12248 22986 12300
rect 22281 12223 22339 12229
rect 22066 12192 22232 12220
rect 21571 12183 21629 12189
rect 21361 12155 21419 12161
rect 19996 12124 21220 12152
rect 20530 12084 20536 12096
rect 17828 12056 20536 12084
rect 17828 12044 17834 12056
rect 20530 12044 20536 12056
rect 20588 12044 20594 12096
rect 21192 12084 21220 12124
rect 21361 12121 21373 12155
rect 21407 12152 21419 12155
rect 22002 12152 22008 12164
rect 21407 12124 22008 12152
rect 21407 12121 21419 12124
rect 21361 12115 21419 12121
rect 22002 12112 22008 12124
rect 22060 12112 22066 12164
rect 22204 12152 22232 12192
rect 22281 12189 22293 12223
rect 22327 12189 22339 12223
rect 22281 12183 22339 12189
rect 22373 12223 22431 12229
rect 22373 12189 22385 12223
rect 22419 12220 22431 12223
rect 22738 12220 22744 12232
rect 22419 12192 22744 12220
rect 22419 12189 22431 12192
rect 22373 12183 22431 12189
rect 22388 12152 22416 12183
rect 22738 12180 22744 12192
rect 22796 12180 22802 12232
rect 23014 12180 23020 12232
rect 23072 12180 23078 12232
rect 23198 12180 23204 12232
rect 23256 12180 23262 12232
rect 22204 12124 22416 12152
rect 22462 12112 22468 12164
rect 22520 12152 22526 12164
rect 22557 12155 22615 12161
rect 22557 12152 22569 12155
rect 22520 12124 22569 12152
rect 22520 12112 22526 12124
rect 22557 12121 22569 12124
rect 22603 12152 22615 12155
rect 22646 12152 22652 12164
rect 22603 12124 22652 12152
rect 22603 12121 22615 12124
rect 22557 12115 22615 12121
rect 22646 12112 22652 12124
rect 22704 12112 22710 12164
rect 22370 12084 22376 12096
rect 21192 12056 22376 12084
rect 22370 12044 22376 12056
rect 22428 12084 22434 12096
rect 23109 12087 23167 12093
rect 23109 12084 23121 12087
rect 22428 12056 23121 12084
rect 22428 12044 22434 12056
rect 23109 12053 23121 12056
rect 23155 12053 23167 12087
rect 23109 12047 23167 12053
rect 1104 11994 23987 12016
rect 1104 11942 6630 11994
rect 6682 11942 6694 11994
rect 6746 11942 6758 11994
rect 6810 11942 6822 11994
rect 6874 11942 6886 11994
rect 6938 11942 12311 11994
rect 12363 11942 12375 11994
rect 12427 11942 12439 11994
rect 12491 11942 12503 11994
rect 12555 11942 12567 11994
rect 12619 11942 17992 11994
rect 18044 11942 18056 11994
rect 18108 11942 18120 11994
rect 18172 11942 18184 11994
rect 18236 11942 18248 11994
rect 18300 11942 23673 11994
rect 23725 11942 23737 11994
rect 23789 11942 23801 11994
rect 23853 11942 23865 11994
rect 23917 11942 23929 11994
rect 23981 11942 23987 11994
rect 1104 11920 23987 11942
rect 4338 11840 4344 11892
rect 4396 11840 4402 11892
rect 4798 11840 4804 11892
rect 4856 11880 4862 11892
rect 5074 11880 5080 11892
rect 4856 11852 5080 11880
rect 4856 11840 4862 11852
rect 5074 11840 5080 11852
rect 5132 11880 5138 11892
rect 5810 11880 5816 11892
rect 5132 11852 5816 11880
rect 5132 11840 5138 11852
rect 5810 11840 5816 11852
rect 5868 11840 5874 11892
rect 6178 11840 6184 11892
rect 6236 11880 6242 11892
rect 6549 11883 6607 11889
rect 6549 11880 6561 11883
rect 6236 11852 6561 11880
rect 6236 11840 6242 11852
rect 6549 11849 6561 11852
rect 6595 11849 6607 11883
rect 6549 11843 6607 11849
rect 7190 11840 7196 11892
rect 7248 11880 7254 11892
rect 8573 11883 8631 11889
rect 8573 11880 8585 11883
rect 7248 11852 8585 11880
rect 7248 11840 7254 11852
rect 8573 11849 8585 11852
rect 8619 11849 8631 11883
rect 8573 11843 8631 11849
rect 11422 11840 11428 11892
rect 11480 11880 11486 11892
rect 12066 11880 12072 11892
rect 11480 11852 12072 11880
rect 11480 11840 11486 11852
rect 12066 11840 12072 11852
rect 12124 11880 12130 11892
rect 12621 11883 12679 11889
rect 12621 11880 12633 11883
rect 12124 11852 12633 11880
rect 12124 11840 12130 11852
rect 12621 11849 12633 11852
rect 12667 11849 12679 11883
rect 12621 11843 12679 11849
rect 13262 11840 13268 11892
rect 13320 11880 13326 11892
rect 13320 11852 14504 11880
rect 13320 11840 13326 11852
rect 1854 11772 1860 11824
rect 1912 11812 1918 11824
rect 1912 11784 2774 11812
rect 1912 11772 1918 11784
rect 2746 11744 2774 11784
rect 3510 11772 3516 11824
rect 3568 11812 3574 11824
rect 5169 11815 5227 11821
rect 5169 11812 5181 11815
rect 3568 11784 5181 11812
rect 3568 11772 3574 11784
rect 5169 11781 5181 11784
rect 5215 11781 5227 11815
rect 5902 11812 5908 11824
rect 5169 11775 5227 11781
rect 5276 11784 5908 11812
rect 3927 11747 3985 11753
rect 3927 11744 3939 11747
rect 2746 11716 3939 11744
rect 3927 11713 3939 11716
rect 3973 11744 3985 11747
rect 5276 11744 5304 11784
rect 5902 11772 5908 11784
rect 5960 11772 5966 11824
rect 6454 11772 6460 11824
rect 6512 11812 6518 11824
rect 6825 11815 6883 11821
rect 6825 11812 6837 11815
rect 6512 11784 6837 11812
rect 6512 11772 6518 11784
rect 6825 11781 6837 11784
rect 6871 11781 6883 11815
rect 8941 11815 8999 11821
rect 6825 11775 6883 11781
rect 6932 11784 8800 11812
rect 6932 11756 6960 11784
rect 8772 11756 8800 11784
rect 8941 11781 8953 11815
rect 8987 11812 8999 11815
rect 10502 11812 10508 11824
rect 8987 11784 10508 11812
rect 8987 11781 8999 11784
rect 8941 11775 8999 11781
rect 10502 11772 10508 11784
rect 10560 11772 10566 11824
rect 12158 11772 12164 11824
rect 12216 11812 12222 11824
rect 12710 11812 12716 11824
rect 12216 11784 12716 11812
rect 12216 11772 12222 11784
rect 12710 11772 12716 11784
rect 12768 11812 12774 11824
rect 13541 11815 13599 11821
rect 13541 11812 13553 11815
rect 12768 11784 13553 11812
rect 12768 11772 12774 11784
rect 13541 11781 13553 11784
rect 13587 11781 13599 11815
rect 13541 11775 13599 11781
rect 13906 11772 13912 11824
rect 13964 11812 13970 11824
rect 14090 11812 14096 11824
rect 13964 11784 14096 11812
rect 13964 11772 13970 11784
rect 14090 11772 14096 11784
rect 14148 11772 14154 11824
rect 14182 11772 14188 11824
rect 14240 11812 14246 11824
rect 14369 11815 14427 11821
rect 14369 11812 14381 11815
rect 14240 11784 14381 11812
rect 14240 11772 14246 11784
rect 14369 11781 14381 11784
rect 14415 11781 14427 11815
rect 14476 11812 14504 11852
rect 14550 11840 14556 11892
rect 14608 11880 14614 11892
rect 15197 11883 15255 11889
rect 15197 11880 15209 11883
rect 14608 11852 15209 11880
rect 14608 11840 14614 11852
rect 15197 11849 15209 11852
rect 15243 11880 15255 11883
rect 15378 11880 15384 11892
rect 15243 11852 15384 11880
rect 15243 11849 15255 11852
rect 15197 11843 15255 11849
rect 15378 11840 15384 11852
rect 15436 11840 15442 11892
rect 15565 11883 15623 11889
rect 15565 11849 15577 11883
rect 15611 11880 15623 11883
rect 15930 11880 15936 11892
rect 15611 11852 15936 11880
rect 15611 11849 15623 11852
rect 15565 11843 15623 11849
rect 15930 11840 15936 11852
rect 15988 11840 15994 11892
rect 17310 11880 17316 11892
rect 16868 11852 17316 11880
rect 15289 11815 15347 11821
rect 15289 11812 15301 11815
rect 14476 11784 15301 11812
rect 14369 11775 14427 11781
rect 15289 11781 15301 11784
rect 15335 11812 15347 11815
rect 16574 11812 16580 11824
rect 15335 11784 16580 11812
rect 15335 11781 15347 11784
rect 15289 11775 15347 11781
rect 16574 11772 16580 11784
rect 16632 11772 16638 11824
rect 3973 11716 5304 11744
rect 3973 11713 3985 11716
rect 3927 11707 3985 11713
rect 5350 11704 5356 11756
rect 5408 11704 5414 11756
rect 5442 11704 5448 11756
rect 5500 11704 5506 11756
rect 5534 11704 5540 11756
rect 5592 11704 5598 11756
rect 5675 11747 5733 11753
rect 5675 11713 5687 11747
rect 5721 11744 5733 11747
rect 5721 11716 5948 11744
rect 5721 11713 5733 11716
rect 5675 11707 5733 11713
rect 5920 11688 5948 11716
rect 6730 11704 6736 11756
rect 6788 11704 6794 11756
rect 6914 11704 6920 11756
rect 6972 11704 6978 11756
rect 7035 11747 7093 11753
rect 7035 11713 7047 11747
rect 7081 11744 7093 11747
rect 7081 11716 8708 11744
rect 7081 11713 7093 11716
rect 7035 11707 7093 11713
rect 2774 11636 2780 11688
rect 2832 11676 2838 11688
rect 3694 11676 3700 11688
rect 2832 11648 3700 11676
rect 2832 11636 2838 11648
rect 3694 11636 3700 11648
rect 3752 11636 3758 11688
rect 3786 11636 3792 11688
rect 3844 11636 3850 11688
rect 4065 11679 4123 11685
rect 4065 11645 4077 11679
rect 4111 11645 4123 11679
rect 4065 11639 4123 11645
rect 3804 11608 3832 11636
rect 3712 11580 3832 11608
rect 4080 11608 4108 11639
rect 4154 11636 4160 11688
rect 4212 11636 4218 11688
rect 5810 11636 5816 11688
rect 5868 11636 5874 11688
rect 5902 11636 5908 11688
rect 5960 11676 5966 11688
rect 7050 11676 7078 11707
rect 5960 11648 7078 11676
rect 5960 11636 5966 11648
rect 7190 11636 7196 11688
rect 7248 11636 7254 11688
rect 8680 11676 8708 11716
rect 8754 11704 8760 11756
rect 8812 11704 8818 11756
rect 8846 11704 8852 11756
rect 8904 11704 8910 11756
rect 9059 11747 9117 11753
rect 9059 11713 9071 11747
rect 9105 11713 9117 11747
rect 9059 11707 9117 11713
rect 8938 11676 8944 11688
rect 8680 11648 8944 11676
rect 8938 11636 8944 11648
rect 8996 11676 9002 11688
rect 9074 11676 9102 11707
rect 10042 11704 10048 11756
rect 10100 11704 10106 11756
rect 10134 11704 10140 11756
rect 10192 11744 10198 11756
rect 10597 11747 10655 11753
rect 10597 11744 10609 11747
rect 10192 11716 10609 11744
rect 10192 11704 10198 11716
rect 10597 11713 10609 11716
rect 10643 11713 10655 11747
rect 10597 11707 10655 11713
rect 12066 11704 12072 11756
rect 12124 11744 12130 11756
rect 13449 11747 13507 11753
rect 13449 11744 13461 11747
rect 12124 11716 13461 11744
rect 12124 11704 12130 11716
rect 13449 11713 13461 11716
rect 13495 11713 13507 11747
rect 13449 11707 13507 11713
rect 13814 11704 13820 11756
rect 13872 11744 13878 11756
rect 14458 11744 14464 11756
rect 13872 11716 14464 11744
rect 13872 11704 13878 11716
rect 14458 11704 14464 11716
rect 14516 11704 14522 11756
rect 15010 11704 15016 11756
rect 15068 11704 15074 11756
rect 15381 11747 15439 11753
rect 15381 11713 15393 11747
rect 15427 11744 15439 11747
rect 15838 11744 15844 11756
rect 15427 11716 15844 11744
rect 15427 11713 15439 11716
rect 15381 11707 15439 11713
rect 15838 11704 15844 11716
rect 15896 11704 15902 11756
rect 16868 11753 16896 11852
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 17402 11840 17408 11892
rect 17460 11840 17466 11892
rect 19978 11840 19984 11892
rect 20036 11880 20042 11892
rect 20717 11883 20775 11889
rect 20717 11880 20729 11883
rect 20036 11852 20729 11880
rect 20036 11840 20042 11852
rect 20717 11849 20729 11852
rect 20763 11849 20775 11883
rect 20717 11843 20775 11849
rect 22002 11840 22008 11892
rect 22060 11880 22066 11892
rect 22189 11883 22247 11889
rect 22189 11880 22201 11883
rect 22060 11852 22201 11880
rect 22060 11840 22066 11852
rect 22189 11849 22201 11852
rect 22235 11849 22247 11883
rect 22189 11843 22247 11849
rect 22554 11812 22560 11824
rect 16960 11784 22560 11812
rect 16960 11753 16988 11784
rect 16853 11747 16911 11753
rect 16853 11713 16865 11747
rect 16899 11713 16911 11747
rect 16853 11707 16911 11713
rect 16945 11747 17003 11753
rect 16945 11713 16957 11747
rect 16991 11713 17003 11747
rect 16945 11707 17003 11713
rect 17034 11704 17040 11756
rect 17092 11744 17098 11756
rect 17129 11747 17187 11753
rect 17129 11744 17141 11747
rect 17092 11716 17141 11744
rect 17092 11704 17098 11716
rect 17129 11713 17141 11716
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 17221 11747 17279 11753
rect 17221 11713 17233 11747
rect 17267 11744 17279 11747
rect 17586 11744 17592 11756
rect 17267 11716 17592 11744
rect 17267 11713 17279 11716
rect 17221 11707 17279 11713
rect 8996 11648 9102 11676
rect 9217 11679 9275 11685
rect 8996 11636 9002 11648
rect 9217 11645 9229 11679
rect 9263 11645 9275 11679
rect 9217 11639 9275 11645
rect 9953 11679 10011 11685
rect 9953 11645 9965 11679
rect 9999 11676 10011 11679
rect 10226 11676 10232 11688
rect 9999 11648 10232 11676
rect 9999 11645 10011 11648
rect 9953 11639 10011 11645
rect 5166 11608 5172 11620
rect 4080 11580 5172 11608
rect 3712 11552 3740 11580
rect 5166 11568 5172 11580
rect 5224 11568 5230 11620
rect 5534 11568 5540 11620
rect 5592 11608 5598 11620
rect 6914 11608 6920 11620
rect 5592 11580 6920 11608
rect 5592 11568 5598 11580
rect 6914 11568 6920 11580
rect 6972 11568 6978 11620
rect 7282 11568 7288 11620
rect 7340 11608 7346 11620
rect 8021 11611 8079 11617
rect 8021 11608 8033 11611
rect 7340 11580 8033 11608
rect 7340 11568 7346 11580
rect 8021 11577 8033 11580
rect 8067 11608 8079 11611
rect 9232 11608 9260 11639
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 13354 11636 13360 11688
rect 13412 11636 13418 11688
rect 13998 11636 14004 11688
rect 14056 11676 14062 11688
rect 15028 11676 15056 11704
rect 14056 11648 16344 11676
rect 14056 11636 14062 11648
rect 8067 11580 9260 11608
rect 8067 11577 8079 11580
rect 8021 11571 8079 11577
rect 14274 11568 14280 11620
rect 14332 11608 14338 11620
rect 15013 11611 15071 11617
rect 15013 11608 15025 11611
rect 14332 11580 15025 11608
rect 14332 11568 14338 11580
rect 15013 11577 15025 11580
rect 15059 11577 15071 11611
rect 15013 11571 15071 11577
rect 16316 11552 16344 11648
rect 16758 11636 16764 11688
rect 16816 11676 16822 11688
rect 17236 11676 17264 11707
rect 17586 11704 17592 11716
rect 17644 11704 17650 11756
rect 20530 11704 20536 11756
rect 20588 11744 20594 11756
rect 21100 11753 21128 11784
rect 22554 11772 22560 11784
rect 22612 11772 22618 11824
rect 22738 11772 22744 11824
rect 22796 11772 22802 11824
rect 20901 11747 20959 11753
rect 20901 11744 20913 11747
rect 20588 11716 20913 11744
rect 20588 11704 20594 11716
rect 20901 11713 20913 11716
rect 20947 11713 20959 11747
rect 20901 11707 20959 11713
rect 21085 11747 21143 11753
rect 21085 11713 21097 11747
rect 21131 11713 21143 11747
rect 21085 11707 21143 11713
rect 21358 11704 21364 11756
rect 21416 11744 21422 11756
rect 22097 11747 22155 11753
rect 22097 11744 22109 11747
rect 21416 11716 22109 11744
rect 21416 11704 21422 11716
rect 22097 11713 22109 11716
rect 22143 11713 22155 11747
rect 22097 11707 22155 11713
rect 22281 11747 22339 11753
rect 22281 11713 22293 11747
rect 22327 11744 22339 11747
rect 22756 11744 22784 11772
rect 22327 11716 22784 11744
rect 22327 11713 22339 11716
rect 22281 11707 22339 11713
rect 16816 11648 17264 11676
rect 16816 11636 16822 11648
rect 17862 11636 17868 11688
rect 17920 11636 17926 11688
rect 20162 11636 20168 11688
rect 20220 11676 20226 11688
rect 20438 11676 20444 11688
rect 20220 11648 20444 11676
rect 20220 11636 20226 11648
rect 20438 11636 20444 11648
rect 20496 11676 20502 11688
rect 23014 11676 23020 11688
rect 20496 11648 23020 11676
rect 20496 11636 20502 11648
rect 23014 11636 23020 11648
rect 23072 11636 23078 11688
rect 16850 11568 16856 11620
rect 16908 11608 16914 11620
rect 19337 11611 19395 11617
rect 19337 11608 19349 11611
rect 16908 11580 19349 11608
rect 16908 11568 16914 11580
rect 19337 11577 19349 11580
rect 19383 11608 19395 11611
rect 19794 11608 19800 11620
rect 19383 11580 19800 11608
rect 19383 11577 19395 11580
rect 19337 11571 19395 11577
rect 19794 11568 19800 11580
rect 19852 11568 19858 11620
rect 20254 11568 20260 11620
rect 20312 11608 20318 11620
rect 21358 11608 21364 11620
rect 20312 11580 21364 11608
rect 20312 11568 20318 11580
rect 21358 11568 21364 11580
rect 21416 11568 21422 11620
rect 3694 11500 3700 11552
rect 3752 11500 3758 11552
rect 9122 11500 9128 11552
rect 9180 11540 9186 11552
rect 9582 11540 9588 11552
rect 9180 11512 9588 11540
rect 9180 11500 9186 11512
rect 9582 11500 9588 11512
rect 9640 11540 9646 11552
rect 9769 11543 9827 11549
rect 9769 11540 9781 11543
rect 9640 11512 9781 11540
rect 9640 11500 9646 11512
rect 9769 11509 9781 11512
rect 9815 11509 9827 11543
rect 9769 11503 9827 11509
rect 11238 11500 11244 11552
rect 11296 11540 11302 11552
rect 11698 11540 11704 11552
rect 11296 11512 11704 11540
rect 11296 11500 11302 11512
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 16206 11500 16212 11552
rect 16264 11500 16270 11552
rect 16298 11500 16304 11552
rect 16356 11540 16362 11552
rect 18509 11543 18567 11549
rect 18509 11540 18521 11543
rect 16356 11512 18521 11540
rect 16356 11500 16362 11512
rect 18509 11509 18521 11512
rect 18555 11540 18567 11543
rect 18690 11540 18696 11552
rect 18555 11512 18696 11540
rect 18555 11509 18567 11512
rect 18509 11503 18567 11509
rect 18690 11500 18696 11512
rect 18748 11540 18754 11552
rect 19702 11540 19708 11552
rect 18748 11512 19708 11540
rect 18748 11500 18754 11512
rect 19702 11500 19708 11512
rect 19760 11500 19766 11552
rect 20438 11500 20444 11552
rect 20496 11540 20502 11552
rect 20901 11543 20959 11549
rect 20901 11540 20913 11543
rect 20496 11512 20913 11540
rect 20496 11500 20502 11512
rect 20901 11509 20913 11512
rect 20947 11509 20959 11543
rect 20901 11503 20959 11509
rect 1104 11450 23828 11472
rect 1104 11398 3790 11450
rect 3842 11398 3854 11450
rect 3906 11398 3918 11450
rect 3970 11398 3982 11450
rect 4034 11398 4046 11450
rect 4098 11398 9471 11450
rect 9523 11398 9535 11450
rect 9587 11398 9599 11450
rect 9651 11398 9663 11450
rect 9715 11398 9727 11450
rect 9779 11398 15152 11450
rect 15204 11398 15216 11450
rect 15268 11398 15280 11450
rect 15332 11398 15344 11450
rect 15396 11398 15408 11450
rect 15460 11398 20833 11450
rect 20885 11398 20897 11450
rect 20949 11398 20961 11450
rect 21013 11398 21025 11450
rect 21077 11398 21089 11450
rect 21141 11398 23828 11450
rect 1104 11376 23828 11398
rect 1857 11339 1915 11345
rect 1857 11305 1869 11339
rect 1903 11336 1915 11339
rect 1946 11336 1952 11348
rect 1903 11308 1952 11336
rect 1903 11305 1915 11308
rect 1857 11299 1915 11305
rect 1946 11296 1952 11308
rect 2004 11296 2010 11348
rect 5442 11296 5448 11348
rect 5500 11336 5506 11348
rect 7926 11336 7932 11348
rect 5500 11308 7932 11336
rect 5500 11296 5506 11308
rect 7926 11296 7932 11308
rect 7984 11296 7990 11348
rect 11793 11339 11851 11345
rect 11793 11305 11805 11339
rect 11839 11336 11851 11339
rect 12621 11339 12679 11345
rect 12621 11336 12633 11339
rect 11839 11308 12633 11336
rect 11839 11305 11851 11308
rect 11793 11299 11851 11305
rect 12621 11305 12633 11308
rect 12667 11336 12679 11339
rect 13078 11336 13084 11348
rect 12667 11308 13084 11336
rect 12667 11305 12679 11308
rect 12621 11299 12679 11305
rect 13078 11296 13084 11308
rect 13136 11296 13142 11348
rect 13173 11339 13231 11345
rect 13173 11305 13185 11339
rect 13219 11336 13231 11339
rect 13538 11336 13544 11348
rect 13219 11308 13544 11336
rect 13219 11305 13231 11308
rect 13173 11299 13231 11305
rect 4154 11228 4160 11280
rect 4212 11268 4218 11280
rect 4525 11271 4583 11277
rect 4525 11268 4537 11271
rect 4212 11240 4537 11268
rect 4212 11228 4218 11240
rect 4525 11237 4537 11240
rect 4571 11268 4583 11271
rect 5626 11268 5632 11280
rect 4571 11240 5632 11268
rect 4571 11237 4583 11240
rect 4525 11231 4583 11237
rect 5626 11228 5632 11240
rect 5684 11228 5690 11280
rect 6638 11228 6644 11280
rect 6696 11268 6702 11280
rect 6696 11240 8248 11268
rect 6696 11228 6702 11240
rect 3694 11200 3700 11212
rect 2700 11172 3700 11200
rect 1578 11092 1584 11144
rect 1636 11092 1642 11144
rect 1854 11092 1860 11144
rect 1912 11132 1918 11144
rect 2700 11141 2728 11172
rect 3694 11160 3700 11172
rect 3752 11160 3758 11212
rect 4249 11203 4307 11209
rect 4249 11169 4261 11203
rect 4295 11200 4307 11203
rect 4430 11200 4436 11212
rect 4295 11172 4436 11200
rect 4295 11169 4307 11172
rect 4249 11163 4307 11169
rect 4430 11160 4436 11172
rect 4488 11160 4494 11212
rect 2133 11135 2191 11141
rect 2133 11132 2145 11135
rect 1912 11104 2145 11132
rect 1912 11092 1918 11104
rect 2133 11101 2145 11104
rect 2179 11101 2191 11135
rect 2133 11095 2191 11101
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11101 2743 11135
rect 2685 11095 2743 11101
rect 2774 11092 2780 11144
rect 2832 11132 2838 11144
rect 2961 11135 3019 11141
rect 2961 11132 2973 11135
rect 2832 11104 2973 11132
rect 2832 11092 2838 11104
rect 2961 11101 2973 11104
rect 3007 11101 3019 11135
rect 2961 11095 3019 11101
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 4522 11132 4528 11144
rect 4203 11104 4528 11132
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 4522 11092 4528 11104
rect 4580 11092 4586 11144
rect 5442 11092 5448 11144
rect 5500 11132 5506 11144
rect 6086 11132 6092 11144
rect 5500 11104 6092 11132
rect 5500 11092 5506 11104
rect 6086 11092 6092 11104
rect 6144 11132 6150 11144
rect 8220 11141 8248 11240
rect 11606 11228 11612 11280
rect 11664 11268 11670 11280
rect 13188 11268 13216 11299
rect 13538 11296 13544 11308
rect 13596 11336 13602 11348
rect 14369 11339 14427 11345
rect 14369 11336 14381 11339
rect 13596 11308 14381 11336
rect 13596 11296 13602 11308
rect 14369 11305 14381 11308
rect 14415 11336 14427 11339
rect 14550 11336 14556 11348
rect 14415 11308 14556 11336
rect 14415 11305 14427 11308
rect 14369 11299 14427 11305
rect 14550 11296 14556 11308
rect 14608 11296 14614 11348
rect 14734 11296 14740 11348
rect 14792 11336 14798 11348
rect 14829 11339 14887 11345
rect 14829 11336 14841 11339
rect 14792 11308 14841 11336
rect 14792 11296 14798 11308
rect 14829 11305 14841 11308
rect 14875 11305 14887 11339
rect 16482 11336 16488 11348
rect 14829 11299 14887 11305
rect 15212 11308 16488 11336
rect 11664 11240 13216 11268
rect 11664 11228 11670 11240
rect 8938 11160 8944 11212
rect 8996 11200 9002 11212
rect 9309 11203 9367 11209
rect 9309 11200 9321 11203
rect 8996 11172 9321 11200
rect 8996 11160 9002 11172
rect 9309 11169 9321 11172
rect 9355 11200 9367 11203
rect 10318 11200 10324 11212
rect 9355 11172 10324 11200
rect 9355 11169 9367 11172
rect 9309 11163 9367 11169
rect 10318 11160 10324 11172
rect 10376 11160 10382 11212
rect 10410 11160 10416 11212
rect 10468 11200 10474 11212
rect 14090 11200 14096 11212
rect 10468 11172 14096 11200
rect 10468 11160 10474 11172
rect 14090 11160 14096 11172
rect 14148 11160 14154 11212
rect 15212 11200 15240 11308
rect 16482 11296 16488 11308
rect 16540 11296 16546 11348
rect 16666 11296 16672 11348
rect 16724 11336 16730 11348
rect 16853 11339 16911 11345
rect 16853 11336 16865 11339
rect 16724 11308 16865 11336
rect 16724 11296 16730 11308
rect 16853 11305 16865 11308
rect 16899 11305 16911 11339
rect 16853 11299 16911 11305
rect 18322 11296 18328 11348
rect 18380 11336 18386 11348
rect 18509 11339 18567 11345
rect 18509 11336 18521 11339
rect 18380 11308 18521 11336
rect 18380 11296 18386 11308
rect 18509 11305 18521 11308
rect 18555 11305 18567 11339
rect 18509 11299 18567 11305
rect 20070 11296 20076 11348
rect 20128 11296 20134 11348
rect 20346 11296 20352 11348
rect 20404 11336 20410 11348
rect 22925 11339 22983 11345
rect 22925 11336 22937 11339
rect 20404 11308 22937 11336
rect 20404 11296 20410 11308
rect 22925 11305 22937 11308
rect 22971 11305 22983 11339
rect 22925 11299 22983 11305
rect 15654 11228 15660 11280
rect 15712 11268 15718 11280
rect 22370 11268 22376 11280
rect 15712 11240 17034 11268
rect 15712 11228 15718 11240
rect 15120 11172 15240 11200
rect 7469 11135 7527 11141
rect 7469 11132 7481 11135
rect 6144 11104 7481 11132
rect 6144 11092 6150 11104
rect 7469 11101 7481 11104
rect 7515 11101 7527 11135
rect 7469 11095 7527 11101
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11132 8263 11135
rect 9030 11132 9036 11144
rect 8251 11104 9036 11132
rect 8251 11101 8263 11104
rect 8205 11095 8263 11101
rect 6362 11024 6368 11076
rect 6420 11064 6426 11076
rect 7484 11064 7512 11095
rect 9030 11092 9036 11104
rect 9088 11092 9094 11144
rect 9398 11092 9404 11144
rect 9456 11132 9462 11144
rect 9585 11135 9643 11141
rect 9585 11132 9597 11135
rect 9456 11104 9597 11132
rect 9456 11092 9462 11104
rect 9585 11101 9597 11104
rect 9631 11101 9643 11135
rect 9585 11095 9643 11101
rect 11698 11092 11704 11144
rect 11756 11132 11762 11144
rect 15120 11141 15148 11172
rect 15746 11160 15752 11212
rect 15804 11200 15810 11212
rect 15933 11203 15991 11209
rect 15933 11200 15945 11203
rect 15804 11172 15945 11200
rect 15804 11160 15810 11172
rect 15933 11169 15945 11172
rect 15979 11169 15991 11203
rect 15933 11163 15991 11169
rect 16022 11160 16028 11212
rect 16080 11200 16086 11212
rect 17006 11200 17034 11240
rect 17144 11240 19334 11268
rect 17144 11200 17172 11240
rect 16080 11172 16160 11200
rect 17006 11172 17172 11200
rect 16080 11160 16086 11172
rect 12069 11135 12127 11141
rect 12069 11132 12081 11135
rect 11756 11104 12081 11132
rect 11756 11092 11762 11104
rect 12069 11101 12081 11104
rect 12115 11101 12127 11135
rect 12069 11095 12127 11101
rect 15105 11135 15163 11141
rect 15105 11101 15117 11135
rect 15151 11101 15163 11135
rect 15105 11095 15163 11101
rect 15197 11135 15255 11141
rect 15197 11101 15209 11135
rect 15243 11101 15255 11135
rect 15197 11095 15255 11101
rect 9858 11064 9864 11076
rect 6420 11036 6854 11064
rect 7484 11036 9864 11064
rect 6420 11024 6426 11036
rect 9858 11024 9864 11036
rect 9916 11024 9922 11076
rect 10134 11024 10140 11076
rect 10192 11024 10198 11076
rect 11606 11024 11612 11076
rect 11664 11024 11670 11076
rect 11790 11024 11796 11076
rect 11848 11064 11854 11076
rect 13262 11064 13268 11076
rect 11848 11036 13268 11064
rect 11848 11024 11854 11036
rect 13262 11024 13268 11036
rect 13320 11024 13326 11076
rect 13725 11067 13783 11073
rect 13725 11033 13737 11067
rect 13771 11064 13783 11067
rect 13814 11064 13820 11076
rect 13771 11036 13820 11064
rect 13771 11033 13783 11036
rect 13725 11027 13783 11033
rect 13814 11024 13820 11036
rect 13872 11024 13878 11076
rect 14918 11024 14924 11076
rect 14976 11064 14982 11076
rect 15212 11064 15240 11095
rect 15286 11092 15292 11144
rect 15344 11092 15350 11144
rect 16132 11141 16160 11172
rect 15473 11135 15531 11141
rect 15473 11101 15485 11135
rect 15519 11101 15531 11135
rect 15473 11095 15531 11101
rect 16117 11135 16175 11141
rect 16117 11101 16129 11135
rect 16163 11101 16175 11135
rect 16117 11095 16175 11101
rect 14976 11036 15240 11064
rect 15488 11064 15516 11095
rect 16298 11092 16304 11144
rect 16356 11092 16362 11144
rect 17034 11092 17040 11144
rect 17092 11092 17098 11144
rect 17144 11141 17172 11172
rect 17494 11160 17500 11212
rect 17552 11200 17558 11212
rect 18417 11203 18475 11209
rect 18417 11200 18429 11203
rect 17552 11172 18429 11200
rect 17552 11160 17558 11172
rect 18417 11169 18429 11172
rect 18463 11169 18475 11203
rect 18417 11163 18475 11169
rect 18506 11160 18512 11212
rect 18564 11200 18570 11212
rect 18601 11203 18659 11209
rect 18601 11200 18613 11203
rect 18564 11172 18613 11200
rect 18564 11160 18570 11172
rect 18601 11169 18613 11172
rect 18647 11169 18659 11203
rect 18601 11163 18659 11169
rect 17129 11135 17187 11141
rect 17129 11101 17141 11135
rect 17175 11101 17187 11135
rect 17129 11095 17187 11101
rect 17313 11135 17371 11141
rect 17313 11101 17325 11135
rect 17359 11101 17371 11135
rect 17313 11095 17371 11101
rect 17405 11135 17463 11141
rect 17405 11101 17417 11135
rect 17451 11132 17463 11135
rect 17770 11132 17776 11144
rect 17451 11104 17776 11132
rect 17451 11101 17463 11104
rect 17405 11095 17463 11101
rect 16206 11064 16212 11076
rect 15488 11036 16212 11064
rect 14976 11024 14982 11036
rect 5994 10956 6000 11008
rect 6052 10996 6058 11008
rect 6270 10996 6276 11008
rect 6052 10968 6276 10996
rect 6052 10956 6058 10968
rect 6270 10956 6276 10968
rect 6328 10996 6334 11008
rect 11238 10996 11244 11008
rect 6328 10968 11244 10996
rect 6328 10956 6334 10968
rect 11238 10956 11244 10968
rect 11296 10956 11302 11008
rect 15212 10996 15240 11036
rect 16206 11024 16212 11036
rect 16264 11024 16270 11076
rect 16482 11024 16488 11076
rect 16540 11064 16546 11076
rect 17328 11064 17356 11095
rect 17770 11092 17776 11104
rect 17828 11092 17834 11144
rect 18693 11135 18751 11141
rect 18693 11101 18705 11135
rect 18739 11101 18751 11135
rect 19306 11132 19334 11240
rect 19720 11240 22376 11268
rect 19720 11141 19748 11240
rect 22370 11228 22376 11240
rect 22428 11268 22434 11280
rect 23198 11268 23204 11280
rect 22428 11240 23204 11268
rect 22428 11228 22434 11240
rect 23198 11228 23204 11240
rect 23256 11228 23262 11280
rect 21910 11160 21916 11212
rect 21968 11160 21974 11212
rect 22278 11160 22284 11212
rect 22336 11200 22342 11212
rect 22336 11172 22784 11200
rect 22336 11160 22342 11172
rect 19705 11135 19763 11141
rect 19705 11132 19717 11135
rect 19306 11104 19717 11132
rect 18693 11095 18751 11101
rect 19705 11101 19717 11104
rect 19751 11101 19763 11135
rect 19705 11095 19763 11101
rect 18414 11064 18420 11076
rect 16540 11036 17080 11064
rect 17328 11036 18420 11064
rect 16540 11024 16546 11036
rect 16942 10996 16948 11008
rect 15212 10968 16948 10996
rect 16942 10956 16948 10968
rect 17000 10956 17006 11008
rect 17052 10996 17080 11036
rect 18414 11024 18420 11036
rect 18472 11024 18478 11076
rect 18506 11024 18512 11076
rect 18564 11064 18570 11076
rect 18708 11064 18736 11095
rect 19794 11092 19800 11144
rect 19852 11132 19858 11144
rect 21358 11132 21364 11144
rect 19852 11104 21364 11132
rect 19852 11092 19858 11104
rect 21358 11092 21364 11104
rect 21416 11132 21422 11144
rect 21726 11132 21732 11144
rect 21416 11104 21732 11132
rect 21416 11092 21422 11104
rect 21726 11092 21732 11104
rect 21784 11092 21790 11144
rect 22094 11092 22100 11144
rect 22152 11132 22158 11144
rect 22373 11135 22431 11141
rect 22373 11132 22385 11135
rect 22152 11104 22385 11132
rect 22152 11092 22158 11104
rect 22373 11101 22385 11104
rect 22419 11101 22431 11135
rect 22373 11095 22431 11101
rect 22462 11092 22468 11144
rect 22520 11092 22526 11144
rect 22646 11092 22652 11144
rect 22704 11092 22710 11144
rect 22756 11141 22784 11172
rect 22741 11135 22799 11141
rect 22741 11101 22753 11135
rect 22787 11101 22799 11135
rect 22741 11095 22799 11101
rect 18564 11036 18736 11064
rect 18564 11024 18570 11036
rect 18782 11024 18788 11076
rect 18840 11064 18846 11076
rect 19058 11064 19064 11076
rect 18840 11036 19064 11064
rect 18840 11024 18846 11036
rect 19058 11024 19064 11036
rect 19116 11064 19122 11076
rect 19116 11036 19472 11064
rect 19116 11024 19122 11036
rect 17865 10999 17923 11005
rect 17865 10996 17877 10999
rect 17052 10968 17877 10996
rect 17865 10965 17877 10968
rect 17911 10996 17923 10999
rect 19242 10996 19248 11008
rect 17911 10968 19248 10996
rect 17911 10965 17923 10968
rect 17865 10959 17923 10965
rect 19242 10956 19248 10968
rect 19300 10956 19306 11008
rect 19444 10996 19472 11036
rect 19518 11024 19524 11076
rect 19576 11024 19582 11076
rect 19889 11067 19947 11073
rect 19889 11064 19901 11067
rect 19628 11036 19901 11064
rect 19628 10996 19656 11036
rect 19889 11033 19901 11036
rect 19935 11033 19947 11067
rect 19889 11027 19947 11033
rect 19444 10968 19656 10996
rect 1104 10906 23987 10928
rect 1104 10854 6630 10906
rect 6682 10854 6694 10906
rect 6746 10854 6758 10906
rect 6810 10854 6822 10906
rect 6874 10854 6886 10906
rect 6938 10854 12311 10906
rect 12363 10854 12375 10906
rect 12427 10854 12439 10906
rect 12491 10854 12503 10906
rect 12555 10854 12567 10906
rect 12619 10854 17992 10906
rect 18044 10854 18056 10906
rect 18108 10854 18120 10906
rect 18172 10854 18184 10906
rect 18236 10854 18248 10906
rect 18300 10854 23673 10906
rect 23725 10854 23737 10906
rect 23789 10854 23801 10906
rect 23853 10854 23865 10906
rect 23917 10854 23929 10906
rect 23981 10854 23987 10906
rect 1104 10832 23987 10854
rect 1578 10752 1584 10804
rect 1636 10792 1642 10804
rect 1765 10795 1823 10801
rect 1765 10792 1777 10795
rect 1636 10764 1777 10792
rect 1636 10752 1642 10764
rect 1765 10761 1777 10764
rect 1811 10761 1823 10795
rect 2958 10792 2964 10804
rect 1765 10755 1823 10761
rect 1964 10764 2964 10792
rect 1964 10665 1992 10764
rect 2958 10752 2964 10764
rect 3016 10792 3022 10804
rect 5074 10792 5080 10804
rect 3016 10764 5080 10792
rect 3016 10752 3022 10764
rect 5074 10752 5080 10764
rect 5132 10752 5138 10804
rect 5350 10752 5356 10804
rect 5408 10792 5414 10804
rect 5445 10795 5503 10801
rect 5445 10792 5457 10795
rect 5408 10764 5457 10792
rect 5408 10752 5414 10764
rect 5445 10761 5457 10764
rect 5491 10761 5503 10795
rect 5445 10755 5503 10761
rect 6546 10752 6552 10804
rect 6604 10792 6610 10804
rect 6733 10795 6791 10801
rect 6733 10792 6745 10795
rect 6604 10764 6745 10792
rect 6604 10752 6610 10764
rect 6733 10761 6745 10764
rect 6779 10761 6791 10795
rect 6733 10755 6791 10761
rect 8754 10752 8760 10804
rect 8812 10792 8818 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 8812 10764 8953 10792
rect 8812 10752 8818 10764
rect 8941 10761 8953 10764
rect 8987 10792 8999 10795
rect 9306 10792 9312 10804
rect 8987 10764 9312 10792
rect 8987 10761 8999 10764
rect 8941 10755 8999 10761
rect 9306 10752 9312 10764
rect 9364 10752 9370 10804
rect 11698 10752 11704 10804
rect 11756 10792 11762 10804
rect 12710 10792 12716 10804
rect 11756 10764 12716 10792
rect 11756 10752 11762 10764
rect 12710 10752 12716 10764
rect 12768 10792 12774 10804
rect 12805 10795 12863 10801
rect 12805 10792 12817 10795
rect 12768 10764 12817 10792
rect 12768 10752 12774 10764
rect 12805 10761 12817 10764
rect 12851 10761 12863 10795
rect 12805 10755 12863 10761
rect 13722 10752 13728 10804
rect 13780 10792 13786 10804
rect 14737 10795 14795 10801
rect 13780 10764 14596 10792
rect 13780 10752 13786 10764
rect 2222 10684 2228 10736
rect 2280 10684 2286 10736
rect 2498 10684 2504 10736
rect 2556 10724 2562 10736
rect 3053 10727 3111 10733
rect 2556 10696 3004 10724
rect 2556 10684 2562 10696
rect 2976 10668 3004 10696
rect 3053 10693 3065 10727
rect 3099 10724 3111 10727
rect 4430 10724 4436 10736
rect 3099 10696 4436 10724
rect 3099 10693 3111 10696
rect 3053 10687 3111 10693
rect 4430 10684 4436 10696
rect 4488 10684 4494 10736
rect 7006 10724 7012 10736
rect 6932 10696 7012 10724
rect 1949 10659 2007 10665
rect 1949 10625 1961 10659
rect 1995 10625 2007 10659
rect 1949 10619 2007 10625
rect 2314 10616 2320 10668
rect 2372 10656 2378 10668
rect 2685 10659 2743 10665
rect 2685 10656 2697 10659
rect 2372 10628 2697 10656
rect 2372 10616 2378 10628
rect 2685 10625 2697 10628
rect 2731 10625 2743 10659
rect 2685 10619 2743 10625
rect 2958 10616 2964 10668
rect 3016 10616 3022 10668
rect 3142 10616 3148 10668
rect 3200 10656 3206 10668
rect 4525 10659 4583 10665
rect 4525 10656 4537 10659
rect 3200 10628 4537 10656
rect 3200 10616 3206 10628
rect 4525 10625 4537 10628
rect 4571 10625 4583 10659
rect 4525 10619 4583 10625
rect 5626 10616 5632 10668
rect 5684 10616 5690 10668
rect 5721 10659 5779 10665
rect 5721 10625 5733 10659
rect 5767 10656 5779 10659
rect 6178 10656 6184 10668
rect 5767 10628 6184 10656
rect 5767 10625 5779 10628
rect 5721 10619 5779 10625
rect 6178 10616 6184 10628
rect 6236 10616 6242 10668
rect 6932 10665 6960 10696
rect 7006 10684 7012 10696
rect 7064 10684 7070 10736
rect 10134 10724 10140 10736
rect 8956 10696 10140 10724
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 7098 10616 7104 10668
rect 7156 10616 7162 10668
rect 7650 10616 7656 10668
rect 7708 10656 7714 10668
rect 7745 10659 7803 10665
rect 7745 10656 7757 10659
rect 7708 10628 7757 10656
rect 7708 10616 7714 10628
rect 7745 10625 7757 10628
rect 7791 10625 7803 10659
rect 7745 10619 7803 10625
rect 7929 10659 7987 10665
rect 7929 10625 7941 10659
rect 7975 10656 7987 10659
rect 8662 10656 8668 10668
rect 7975 10628 8668 10656
rect 7975 10625 7987 10628
rect 7929 10619 7987 10625
rect 8662 10616 8668 10628
rect 8720 10616 8726 10668
rect 8956 10665 8984 10696
rect 10134 10684 10140 10696
rect 10192 10684 10198 10736
rect 11900 10696 12434 10724
rect 8941 10659 8999 10665
rect 8941 10625 8953 10659
rect 8987 10625 8999 10659
rect 8941 10619 8999 10625
rect 9122 10616 9128 10668
rect 9180 10616 9186 10668
rect 9861 10659 9919 10665
rect 9861 10625 9873 10659
rect 9907 10656 9919 10659
rect 9950 10656 9956 10668
rect 9907 10628 9956 10656
rect 9907 10625 9919 10628
rect 9861 10619 9919 10625
rect 9950 10616 9956 10628
rect 10008 10616 10014 10668
rect 10318 10616 10324 10668
rect 10376 10656 10382 10668
rect 11900 10665 11928 10696
rect 11885 10659 11943 10665
rect 11885 10656 11897 10659
rect 10376 10628 11897 10656
rect 10376 10616 10382 10628
rect 11885 10625 11897 10628
rect 11931 10625 11943 10659
rect 11885 10619 11943 10625
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 1670 10548 1676 10600
rect 1728 10588 1734 10600
rect 2041 10591 2099 10597
rect 2041 10588 2053 10591
rect 1728 10560 2053 10588
rect 1728 10548 1734 10560
rect 2041 10557 2053 10560
rect 2087 10588 2099 10591
rect 2406 10588 2412 10600
rect 2087 10560 2412 10588
rect 2087 10557 2099 10560
rect 2041 10551 2099 10557
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 4154 10548 4160 10600
rect 4212 10588 4218 10600
rect 4249 10591 4307 10597
rect 4249 10588 4261 10591
rect 4212 10560 4261 10588
rect 4212 10548 4218 10560
rect 4249 10557 4261 10560
rect 4295 10557 4307 10591
rect 4249 10551 4307 10557
rect 5810 10548 5816 10600
rect 5868 10548 5874 10600
rect 5905 10591 5963 10597
rect 5905 10557 5917 10591
rect 5951 10588 5963 10591
rect 5951 10560 6776 10588
rect 5951 10557 5963 10560
rect 5905 10551 5963 10557
rect 6748 10520 6776 10560
rect 7006 10548 7012 10600
rect 7064 10548 7070 10600
rect 7190 10548 7196 10600
rect 7248 10548 7254 10600
rect 9677 10591 9735 10597
rect 9677 10557 9689 10591
rect 9723 10588 9735 10591
rect 10594 10588 10600 10600
rect 9723 10560 10600 10588
rect 9723 10557 9735 10560
rect 9677 10551 9735 10557
rect 10594 10548 10600 10560
rect 10652 10548 10658 10600
rect 7208 10520 7236 10548
rect 6748 10492 7236 10520
rect 7466 10480 7472 10532
rect 7524 10520 7530 10532
rect 11701 10523 11759 10529
rect 11701 10520 11713 10523
rect 7524 10492 11713 10520
rect 7524 10480 7530 10492
rect 11701 10489 11713 10492
rect 11747 10489 11759 10523
rect 11701 10483 11759 10489
rect 2225 10455 2283 10461
rect 2225 10421 2237 10455
rect 2271 10452 2283 10455
rect 2590 10452 2596 10464
rect 2271 10424 2596 10452
rect 2271 10421 2283 10424
rect 2225 10415 2283 10421
rect 2590 10412 2596 10424
rect 2648 10412 2654 10464
rect 3605 10455 3663 10461
rect 3605 10421 3617 10455
rect 3651 10452 3663 10455
rect 3694 10452 3700 10464
rect 3651 10424 3700 10452
rect 3651 10421 3663 10424
rect 3605 10415 3663 10421
rect 3694 10412 3700 10424
rect 3752 10412 3758 10464
rect 5718 10412 5724 10464
rect 5776 10452 5782 10464
rect 7745 10455 7803 10461
rect 7745 10452 7757 10455
rect 5776 10424 7757 10452
rect 5776 10412 5782 10424
rect 7745 10421 7757 10424
rect 7791 10421 7803 10455
rect 7745 10415 7803 10421
rect 10045 10455 10103 10461
rect 10045 10421 10057 10455
rect 10091 10452 10103 10455
rect 10502 10452 10508 10464
rect 10091 10424 10508 10452
rect 10091 10421 10103 10424
rect 10045 10415 10103 10421
rect 10502 10412 10508 10424
rect 10560 10412 10566 10464
rect 10594 10412 10600 10464
rect 10652 10412 10658 10464
rect 10870 10412 10876 10464
rect 10928 10452 10934 10464
rect 11057 10455 11115 10461
rect 11057 10452 11069 10455
rect 10928 10424 11069 10452
rect 10928 10412 10934 10424
rect 11057 10421 11069 10424
rect 11103 10452 11115 10455
rect 11992 10452 12020 10619
rect 12066 10616 12072 10668
rect 12124 10616 12130 10668
rect 12250 10616 12256 10668
rect 12308 10616 12314 10668
rect 12406 10520 12434 10696
rect 13262 10684 13268 10736
rect 13320 10724 13326 10736
rect 14369 10727 14427 10733
rect 14369 10724 14381 10727
rect 13320 10696 14381 10724
rect 13320 10684 13326 10696
rect 14369 10693 14381 10696
rect 14415 10693 14427 10727
rect 14369 10687 14427 10693
rect 14461 10727 14519 10733
rect 14461 10693 14473 10727
rect 14507 10693 14519 10727
rect 14461 10687 14519 10693
rect 13998 10616 14004 10668
rect 14056 10656 14062 10668
rect 14274 10665 14280 10668
rect 14093 10659 14151 10665
rect 14093 10656 14105 10659
rect 14056 10628 14105 10656
rect 14056 10616 14062 10628
rect 14093 10625 14105 10628
rect 14139 10625 14151 10659
rect 14093 10619 14151 10625
rect 14241 10659 14280 10665
rect 14241 10625 14253 10659
rect 14241 10619 14280 10625
rect 14274 10616 14280 10619
rect 14332 10616 14338 10668
rect 13081 10591 13139 10597
rect 13081 10557 13093 10591
rect 13127 10588 13139 10591
rect 13262 10588 13268 10600
rect 13127 10560 13268 10588
rect 13127 10557 13139 10560
rect 13081 10551 13139 10557
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 14476 10588 14504 10687
rect 14568 10665 14596 10764
rect 14737 10761 14749 10795
rect 14783 10792 14795 10795
rect 15286 10792 15292 10804
rect 14783 10764 15292 10792
rect 14783 10761 14795 10764
rect 14737 10755 14795 10761
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 15562 10752 15568 10804
rect 15620 10792 15626 10804
rect 15620 10764 15976 10792
rect 15620 10752 15626 10764
rect 14558 10659 14616 10665
rect 14558 10625 14570 10659
rect 14604 10625 14616 10659
rect 14558 10619 14616 10625
rect 15194 10616 15200 10668
rect 15252 10656 15258 10668
rect 15565 10659 15623 10665
rect 15565 10656 15577 10659
rect 15252 10628 15577 10656
rect 15252 10616 15258 10628
rect 15565 10625 15577 10628
rect 15611 10625 15623 10659
rect 15565 10619 15623 10625
rect 15657 10659 15715 10665
rect 15657 10625 15669 10659
rect 15703 10625 15715 10659
rect 15657 10619 15715 10625
rect 15672 10588 15700 10619
rect 15838 10616 15844 10668
rect 15896 10616 15902 10668
rect 15948 10665 15976 10764
rect 17126 10752 17132 10804
rect 17184 10792 17190 10804
rect 18325 10795 18383 10801
rect 17184 10764 17540 10792
rect 17184 10752 17190 10764
rect 16574 10684 16580 10736
rect 16632 10724 16638 10736
rect 17512 10733 17540 10764
rect 18325 10761 18337 10795
rect 18371 10792 18383 10795
rect 18414 10792 18420 10804
rect 18371 10764 18420 10792
rect 18371 10761 18383 10764
rect 18325 10755 18383 10761
rect 18414 10752 18420 10764
rect 18472 10752 18478 10804
rect 21358 10752 21364 10804
rect 21416 10752 21422 10804
rect 17497 10727 17555 10733
rect 16632 10696 17448 10724
rect 16632 10684 16638 10696
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10625 15991 10659
rect 15933 10619 15991 10625
rect 16850 10616 16856 10668
rect 16908 10616 16914 10668
rect 17052 10665 17080 10696
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 17129 10659 17187 10665
rect 17129 10625 17141 10659
rect 17175 10625 17187 10659
rect 17129 10619 17187 10625
rect 17222 10659 17280 10665
rect 17222 10625 17234 10659
rect 17268 10656 17280 10659
rect 17310 10656 17316 10668
rect 17268 10628 17316 10656
rect 17268 10625 17280 10628
rect 17222 10619 17280 10625
rect 14476 10560 16528 10588
rect 13170 10520 13176 10532
rect 12406 10492 13176 10520
rect 13170 10480 13176 10492
rect 13228 10480 13234 10532
rect 13633 10523 13691 10529
rect 13633 10489 13645 10523
rect 13679 10520 13691 10523
rect 14182 10520 14188 10532
rect 13679 10492 14188 10520
rect 13679 10489 13691 10492
rect 13633 10483 13691 10489
rect 14182 10480 14188 10492
rect 14240 10480 14246 10532
rect 11103 10424 12020 10452
rect 13265 10455 13323 10461
rect 11103 10421 11115 10424
rect 11057 10415 11115 10421
rect 13265 10421 13277 10455
rect 13311 10452 13323 10455
rect 14366 10452 14372 10464
rect 13311 10424 14372 10452
rect 13311 10421 13323 10424
rect 13265 10415 13323 10421
rect 14366 10412 14372 10424
rect 14424 10412 14430 10464
rect 15381 10455 15439 10461
rect 15381 10421 15393 10455
rect 15427 10452 15439 10455
rect 15562 10452 15568 10464
rect 15427 10424 15568 10452
rect 15427 10421 15439 10424
rect 15381 10415 15439 10421
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 16500 10452 16528 10560
rect 17144 10520 17172 10619
rect 17310 10616 17316 10628
rect 17368 10616 17374 10668
rect 17420 10656 17448 10696
rect 17497 10693 17509 10727
rect 17543 10693 17555 10727
rect 19426 10724 19432 10736
rect 17497 10687 17555 10693
rect 17604 10696 19432 10724
rect 17604 10656 17632 10696
rect 19426 10684 19432 10696
rect 19484 10684 19490 10736
rect 17420 10628 17632 10656
rect 18509 10659 18567 10665
rect 18509 10625 18521 10659
rect 18555 10625 18567 10659
rect 18509 10619 18567 10625
rect 18524 10588 18552 10619
rect 18598 10616 18604 10668
rect 18656 10616 18662 10668
rect 18690 10616 18696 10668
rect 18748 10656 18754 10668
rect 18877 10659 18935 10665
rect 18877 10656 18889 10659
rect 18748 10628 18889 10656
rect 18748 10616 18754 10628
rect 18877 10625 18889 10628
rect 18923 10625 18935 10659
rect 18877 10619 18935 10625
rect 21174 10616 21180 10668
rect 21232 10656 21238 10668
rect 22373 10659 22431 10665
rect 22373 10656 22385 10659
rect 21232 10628 22385 10656
rect 21232 10616 21238 10628
rect 22373 10625 22385 10628
rect 22419 10625 22431 10659
rect 22373 10619 22431 10625
rect 18524 10560 19472 10588
rect 17144 10492 18368 10520
rect 18340 10464 18368 10492
rect 18046 10452 18052 10464
rect 16500 10424 18052 10452
rect 18046 10412 18052 10424
rect 18104 10412 18110 10464
rect 18322 10412 18328 10464
rect 18380 10452 18386 10464
rect 18785 10455 18843 10461
rect 18785 10452 18797 10455
rect 18380 10424 18797 10452
rect 18380 10412 18386 10424
rect 18785 10421 18797 10424
rect 18831 10452 18843 10455
rect 19242 10452 19248 10464
rect 18831 10424 19248 10452
rect 18831 10421 18843 10424
rect 18785 10415 18843 10421
rect 19242 10412 19248 10424
rect 19300 10412 19306 10464
rect 19444 10461 19472 10560
rect 22094 10548 22100 10600
rect 22152 10548 22158 10600
rect 22189 10591 22247 10597
rect 22189 10557 22201 10591
rect 22235 10557 22247 10591
rect 22189 10551 22247 10557
rect 22281 10591 22339 10597
rect 22281 10557 22293 10591
rect 22327 10588 22339 10591
rect 22327 10560 22508 10588
rect 22327 10557 22339 10560
rect 22281 10551 22339 10557
rect 22204 10520 22232 10551
rect 22370 10520 22376 10532
rect 22204 10492 22376 10520
rect 22370 10480 22376 10492
rect 22428 10480 22434 10532
rect 19429 10455 19487 10461
rect 19429 10421 19441 10455
rect 19475 10452 19487 10455
rect 19610 10452 19616 10464
rect 19475 10424 19616 10452
rect 19475 10421 19487 10424
rect 19429 10415 19487 10421
rect 19610 10412 19616 10424
rect 19668 10452 19674 10464
rect 20714 10452 20720 10464
rect 19668 10424 20720 10452
rect 19668 10412 19674 10424
rect 20714 10412 20720 10424
rect 20772 10412 20778 10464
rect 21726 10412 21732 10464
rect 21784 10452 21790 10464
rect 22480 10452 22508 10560
rect 21784 10424 22508 10452
rect 21784 10412 21790 10424
rect 22554 10412 22560 10464
rect 22612 10412 22618 10464
rect 1104 10362 23828 10384
rect 1104 10310 3790 10362
rect 3842 10310 3854 10362
rect 3906 10310 3918 10362
rect 3970 10310 3982 10362
rect 4034 10310 4046 10362
rect 4098 10310 9471 10362
rect 9523 10310 9535 10362
rect 9587 10310 9599 10362
rect 9651 10310 9663 10362
rect 9715 10310 9727 10362
rect 9779 10310 15152 10362
rect 15204 10310 15216 10362
rect 15268 10310 15280 10362
rect 15332 10310 15344 10362
rect 15396 10310 15408 10362
rect 15460 10310 20833 10362
rect 20885 10310 20897 10362
rect 20949 10310 20961 10362
rect 21013 10310 21025 10362
rect 21077 10310 21089 10362
rect 21141 10310 23828 10362
rect 1104 10288 23828 10310
rect 4246 10208 4252 10260
rect 4304 10248 4310 10260
rect 4525 10251 4583 10257
rect 4525 10248 4537 10251
rect 4304 10220 4537 10248
rect 4304 10208 4310 10220
rect 4525 10217 4537 10220
rect 4571 10217 4583 10251
rect 4525 10211 4583 10217
rect 5626 10208 5632 10260
rect 5684 10248 5690 10260
rect 6181 10251 6239 10257
rect 6181 10248 6193 10251
rect 5684 10220 6193 10248
rect 5684 10208 5690 10220
rect 6181 10217 6193 10220
rect 6227 10217 6239 10251
rect 6181 10211 6239 10217
rect 7374 10208 7380 10260
rect 7432 10248 7438 10260
rect 8573 10251 8631 10257
rect 8573 10248 8585 10251
rect 7432 10220 8585 10248
rect 7432 10208 7438 10220
rect 8573 10217 8585 10220
rect 8619 10248 8631 10251
rect 10134 10248 10140 10260
rect 8619 10220 10140 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 10134 10208 10140 10220
rect 10192 10208 10198 10260
rect 13630 10208 13636 10260
rect 13688 10248 13694 10260
rect 15473 10251 15531 10257
rect 15473 10248 15485 10251
rect 13688 10220 15485 10248
rect 13688 10208 13694 10220
rect 15473 10217 15485 10220
rect 15519 10217 15531 10251
rect 15473 10211 15531 10217
rect 15657 10251 15715 10257
rect 15657 10217 15669 10251
rect 15703 10248 15715 10251
rect 17862 10248 17868 10260
rect 15703 10220 17868 10248
rect 15703 10217 15715 10220
rect 15657 10211 15715 10217
rect 17862 10208 17868 10220
rect 17920 10208 17926 10260
rect 18046 10208 18052 10260
rect 18104 10248 18110 10260
rect 18690 10248 18696 10260
rect 18104 10220 18696 10248
rect 18104 10208 18110 10220
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 21637 10251 21695 10257
rect 21637 10217 21649 10251
rect 21683 10248 21695 10251
rect 22462 10248 22468 10260
rect 21683 10220 22468 10248
rect 21683 10217 21695 10220
rect 21637 10211 21695 10217
rect 22462 10208 22468 10220
rect 22520 10208 22526 10260
rect 2498 10180 2504 10192
rect 2056 10152 2504 10180
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10044 2007 10047
rect 2056 10044 2084 10152
rect 2498 10140 2504 10152
rect 2556 10140 2562 10192
rect 3234 10140 3240 10192
rect 3292 10140 3298 10192
rect 5445 10183 5503 10189
rect 5445 10149 5457 10183
rect 5491 10180 5503 10183
rect 7392 10180 7420 10208
rect 10870 10180 10876 10192
rect 5491 10152 7420 10180
rect 9600 10152 10876 10180
rect 5491 10149 5503 10152
rect 5445 10143 5503 10149
rect 2225 10115 2283 10121
rect 2225 10081 2237 10115
rect 2271 10112 2283 10115
rect 2774 10112 2780 10124
rect 2271 10084 2780 10112
rect 2271 10081 2283 10084
rect 2225 10075 2283 10081
rect 2774 10072 2780 10084
rect 2832 10072 2838 10124
rect 4430 10112 4436 10124
rect 2884 10084 3096 10112
rect 1995 10016 2084 10044
rect 2133 10047 2191 10053
rect 1995 10013 2007 10016
rect 1949 10007 2007 10013
rect 2133 10013 2145 10047
rect 2179 10013 2191 10047
rect 2133 10007 2191 10013
rect 2148 9976 2176 10007
rect 2314 9976 2320 9988
rect 2148 9948 2320 9976
rect 2314 9936 2320 9948
rect 2372 9976 2378 9988
rect 2884 9976 2912 10084
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10013 3019 10047
rect 2961 10007 3019 10013
rect 2372 9948 2912 9976
rect 2372 9936 2378 9948
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 2976 9908 3004 10007
rect 3068 9976 3096 10084
rect 3252 10084 4436 10112
rect 3252 10053 3280 10084
rect 4430 10072 4436 10084
rect 4488 10072 4494 10124
rect 5810 10072 5816 10124
rect 5868 10112 5874 10124
rect 5868 10084 6500 10112
rect 5868 10072 5874 10084
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10013 3295 10047
rect 3237 10007 3295 10013
rect 4062 10004 4068 10056
rect 4120 10004 4126 10056
rect 4154 10004 4160 10056
rect 4212 10004 4218 10056
rect 4249 10047 4307 10053
rect 4249 10013 4261 10047
rect 4295 10013 4307 10047
rect 4249 10007 4307 10013
rect 4341 10047 4399 10053
rect 4341 10013 4353 10047
rect 4387 10044 4399 10047
rect 4614 10044 4620 10056
rect 4387 10016 4620 10044
rect 4387 10013 4399 10016
rect 4341 10007 4399 10013
rect 4264 9976 4292 10007
rect 4614 10004 4620 10016
rect 4672 10004 4678 10056
rect 4982 10004 4988 10056
rect 5040 10004 5046 10056
rect 5166 10004 5172 10056
rect 5224 10044 5230 10056
rect 6472 10044 6500 10084
rect 6546 10072 6552 10124
rect 6604 10112 6610 10124
rect 9600 10112 9628 10152
rect 10870 10140 10876 10152
rect 10928 10140 10934 10192
rect 13262 10140 13268 10192
rect 13320 10140 13326 10192
rect 14274 10140 14280 10192
rect 14332 10180 14338 10192
rect 14332 10152 15056 10180
rect 14332 10140 14338 10152
rect 6604 10084 9628 10112
rect 9677 10115 9735 10121
rect 6604 10072 6610 10084
rect 9677 10081 9689 10115
rect 9723 10112 9735 10115
rect 9858 10112 9864 10124
rect 9723 10084 9864 10112
rect 9723 10081 9735 10084
rect 9677 10075 9735 10081
rect 9858 10072 9864 10084
rect 9916 10112 9922 10124
rect 10042 10112 10048 10124
rect 9916 10084 10048 10112
rect 9916 10072 9922 10084
rect 10042 10072 10048 10084
rect 10100 10072 10106 10124
rect 13170 10072 13176 10124
rect 13228 10112 13234 10124
rect 15028 10121 15056 10152
rect 16206 10140 16212 10192
rect 16264 10180 16270 10192
rect 17405 10183 17463 10189
rect 17405 10180 17417 10183
rect 16264 10152 17417 10180
rect 16264 10140 16270 10152
rect 17405 10149 17417 10152
rect 17451 10149 17463 10183
rect 17405 10143 17463 10149
rect 17586 10140 17592 10192
rect 17644 10180 17650 10192
rect 19889 10183 19947 10189
rect 19889 10180 19901 10183
rect 17644 10152 19901 10180
rect 17644 10140 17650 10152
rect 19889 10149 19901 10152
rect 19935 10149 19947 10183
rect 19889 10143 19947 10149
rect 15013 10115 15071 10121
rect 13228 10084 14596 10112
rect 13228 10072 13234 10084
rect 6917 10047 6975 10053
rect 6917 10044 6929 10047
rect 5224 10016 6132 10044
rect 6472 10016 6929 10044
rect 5224 10004 5230 10016
rect 5997 9979 6055 9985
rect 5997 9976 6009 9979
rect 3068 9948 6009 9976
rect 5997 9945 6009 9948
rect 6043 9945 6055 9979
rect 6104 9976 6132 10016
rect 6917 10013 6929 10016
rect 6963 10044 6975 10047
rect 7098 10044 7104 10056
rect 6963 10016 7104 10044
rect 6963 10013 6975 10016
rect 6917 10007 6975 10013
rect 7098 10004 7104 10016
rect 7156 10044 7162 10056
rect 7377 10047 7435 10053
rect 7377 10044 7389 10047
rect 7156 10016 7389 10044
rect 7156 10004 7162 10016
rect 7377 10013 7389 10016
rect 7423 10044 7435 10047
rect 8938 10044 8944 10056
rect 7423 10016 8944 10044
rect 7423 10013 7435 10016
rect 7377 10007 7435 10013
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 9122 10004 9128 10056
rect 9180 10044 9186 10056
rect 9217 10047 9275 10053
rect 9217 10044 9229 10047
rect 9180 10016 9229 10044
rect 9180 10004 9186 10016
rect 9217 10013 9229 10016
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 11698 10004 11704 10056
rect 11756 10004 11762 10056
rect 11974 10004 11980 10056
rect 12032 10004 12038 10056
rect 14274 10004 14280 10056
rect 14332 10004 14338 10056
rect 14366 10004 14372 10056
rect 14424 10004 14430 10056
rect 14568 10053 14596 10084
rect 15013 10081 15025 10115
rect 15059 10112 15071 10115
rect 19150 10112 19156 10124
rect 15059 10084 16344 10112
rect 15059 10081 15071 10084
rect 15013 10075 15071 10081
rect 14553 10047 14611 10053
rect 14553 10013 14565 10047
rect 14599 10044 14611 10047
rect 15102 10044 15108 10056
rect 14599 10016 15108 10044
rect 14599 10013 14611 10016
rect 14553 10007 14611 10013
rect 15102 10004 15108 10016
rect 15160 10004 15166 10056
rect 15470 10004 15476 10056
rect 15528 10044 15534 10056
rect 15528 10016 15884 10044
rect 15528 10004 15534 10016
rect 11796 9988 11848 9994
rect 6197 9979 6255 9985
rect 6197 9976 6209 9979
rect 6104 9948 6209 9976
rect 5997 9939 6055 9945
rect 6197 9945 6209 9948
rect 6243 9945 6255 9979
rect 7558 9976 7564 9988
rect 6197 9939 6255 9945
rect 6288 9948 7564 9976
rect 2832 9880 3004 9908
rect 6012 9908 6040 9939
rect 6288 9908 6316 9948
rect 7558 9936 7564 9948
rect 7616 9936 7622 9988
rect 14384 9976 14412 10004
rect 14826 9976 14832 9988
rect 14384 9948 14832 9976
rect 14826 9936 14832 9948
rect 14884 9936 14890 9988
rect 15562 9936 15568 9988
rect 15620 9985 15626 9988
rect 15856 9985 15884 10016
rect 15620 9979 15683 9985
rect 15620 9945 15637 9979
rect 15671 9945 15683 9979
rect 15620 9939 15683 9945
rect 15841 9979 15899 9985
rect 15841 9945 15853 9979
rect 15887 9976 15899 9979
rect 16206 9976 16212 9988
rect 15887 9948 16212 9976
rect 15887 9945 15899 9948
rect 15841 9939 15899 9945
rect 15620 9936 15626 9939
rect 16206 9936 16212 9948
rect 16264 9936 16270 9988
rect 16316 9976 16344 10084
rect 16408 10084 19156 10112
rect 16408 10053 16436 10084
rect 19150 10072 19156 10084
rect 19208 10072 19214 10124
rect 20806 10072 20812 10124
rect 20864 10112 20870 10124
rect 20864 10084 21312 10112
rect 20864 10072 20870 10084
rect 16393 10047 16451 10053
rect 16393 10013 16405 10047
rect 16439 10013 16451 10047
rect 16393 10007 16451 10013
rect 16574 10004 16580 10056
rect 16632 10004 16638 10056
rect 16850 10004 16856 10056
rect 16908 10044 16914 10056
rect 18049 10047 18107 10053
rect 18049 10044 18061 10047
rect 16908 10016 18061 10044
rect 16908 10004 16914 10016
rect 18049 10013 18061 10016
rect 18095 10013 18107 10047
rect 18049 10007 18107 10013
rect 18233 10047 18291 10053
rect 18233 10013 18245 10047
rect 18279 10013 18291 10047
rect 18233 10007 18291 10013
rect 16868 9976 16896 10004
rect 16316 9948 16896 9976
rect 16942 9936 16948 9988
rect 17000 9936 17006 9988
rect 18248 9976 18276 10007
rect 18322 10004 18328 10056
rect 18380 10004 18386 10056
rect 18414 10004 18420 10056
rect 18472 10004 18478 10056
rect 18506 10004 18512 10056
rect 18564 10004 18570 10056
rect 19426 10044 19432 10056
rect 18616 10016 19432 10044
rect 18616 9976 18644 10016
rect 19426 10004 19432 10016
rect 19484 10004 19490 10056
rect 20073 10047 20131 10053
rect 20073 10013 20085 10047
rect 20119 10044 20131 10047
rect 20254 10044 20260 10056
rect 20119 10016 20260 10044
rect 20119 10013 20131 10016
rect 20073 10007 20131 10013
rect 20254 10004 20260 10016
rect 20312 10004 20318 10056
rect 20533 10047 20591 10053
rect 20533 10013 20545 10047
rect 20579 10044 20591 10047
rect 20622 10044 20628 10056
rect 20579 10016 20628 10044
rect 20579 10013 20591 10016
rect 20533 10007 20591 10013
rect 20622 10004 20628 10016
rect 20680 10044 20686 10056
rect 20993 10047 21051 10053
rect 20993 10044 21005 10047
rect 20680 10016 21005 10044
rect 20680 10004 20686 10016
rect 20993 10013 21005 10016
rect 21039 10013 21051 10047
rect 20993 10007 21051 10013
rect 21082 10004 21088 10056
rect 21140 10044 21146 10056
rect 21284 10053 21312 10084
rect 21177 10047 21235 10053
rect 21177 10044 21189 10047
rect 21140 10016 21189 10044
rect 21140 10004 21146 10016
rect 21177 10013 21189 10016
rect 21223 10013 21235 10047
rect 21177 10007 21235 10013
rect 21269 10047 21327 10053
rect 21269 10013 21281 10047
rect 21315 10013 21327 10047
rect 21269 10007 21327 10013
rect 21358 10004 21364 10056
rect 21416 10004 21422 10056
rect 18248 9948 18644 9976
rect 18693 9979 18751 9985
rect 18693 9945 18705 9979
rect 18739 9976 18751 9979
rect 18739 9948 21956 9976
rect 18739 9945 18751 9948
rect 18693 9939 18751 9945
rect 11796 9930 11848 9936
rect 6012 9880 6316 9908
rect 2832 9868 2838 9880
rect 6362 9868 6368 9920
rect 6420 9868 6426 9920
rect 8938 9868 8944 9920
rect 8996 9908 9002 9920
rect 9401 9911 9459 9917
rect 9401 9908 9413 9911
rect 8996 9880 9413 9908
rect 8996 9868 9002 9880
rect 9401 9877 9413 9880
rect 9447 9908 9459 9911
rect 10229 9911 10287 9917
rect 10229 9908 10241 9911
rect 9447 9880 10241 9908
rect 9447 9877 9459 9880
rect 9401 9871 9459 9877
rect 10229 9877 10241 9880
rect 10275 9877 10287 9911
rect 10229 9871 10287 9877
rect 13262 9868 13268 9920
rect 13320 9908 13326 9920
rect 16574 9908 16580 9920
rect 13320 9880 16580 9908
rect 13320 9868 13326 9880
rect 16574 9868 16580 9880
rect 16632 9868 16638 9920
rect 16960 9908 16988 9936
rect 20162 9908 20168 9920
rect 16960 9880 20168 9908
rect 20162 9868 20168 9880
rect 20220 9868 20226 9920
rect 21928 9908 21956 9948
rect 22278 9908 22284 9920
rect 21928 9880 22284 9908
rect 22278 9868 22284 9880
rect 22336 9868 22342 9920
rect 1104 9818 23987 9840
rect 1104 9766 6630 9818
rect 6682 9766 6694 9818
rect 6746 9766 6758 9818
rect 6810 9766 6822 9818
rect 6874 9766 6886 9818
rect 6938 9766 12311 9818
rect 12363 9766 12375 9818
rect 12427 9766 12439 9818
rect 12491 9766 12503 9818
rect 12555 9766 12567 9818
rect 12619 9766 17992 9818
rect 18044 9766 18056 9818
rect 18108 9766 18120 9818
rect 18172 9766 18184 9818
rect 18236 9766 18248 9818
rect 18300 9766 23673 9818
rect 23725 9766 23737 9818
rect 23789 9766 23801 9818
rect 23853 9766 23865 9818
rect 23917 9766 23929 9818
rect 23981 9766 23987 9818
rect 1104 9744 23987 9766
rect 2222 9664 2228 9716
rect 2280 9664 2286 9716
rect 3145 9707 3203 9713
rect 3145 9673 3157 9707
rect 3191 9704 3203 9707
rect 4062 9704 4068 9716
rect 3191 9676 4068 9704
rect 3191 9673 3203 9676
rect 3145 9667 3203 9673
rect 4062 9664 4068 9676
rect 4120 9664 4126 9716
rect 6178 9664 6184 9716
rect 6236 9704 6242 9716
rect 7006 9704 7012 9716
rect 6236 9676 7012 9704
rect 6236 9664 6242 9676
rect 7006 9664 7012 9676
rect 7064 9664 7070 9716
rect 8205 9707 8263 9713
rect 7208 9676 7512 9704
rect 3602 9596 3608 9648
rect 3660 9636 3666 9648
rect 4893 9639 4951 9645
rect 4893 9636 4905 9639
rect 3660 9608 4905 9636
rect 3660 9596 3666 9608
rect 4893 9605 4905 9608
rect 4939 9605 4951 9639
rect 4893 9599 4951 9605
rect 5169 9639 5227 9645
rect 5169 9605 5181 9639
rect 5215 9636 5227 9639
rect 5534 9636 5540 9648
rect 5215 9608 5540 9636
rect 5215 9605 5227 9608
rect 5169 9599 5227 9605
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 2130 9528 2136 9580
rect 2188 9568 2194 9580
rect 2188 9540 2233 9568
rect 2188 9528 2194 9540
rect 2314 9528 2320 9580
rect 2372 9568 2378 9580
rect 2409 9571 2467 9577
rect 2409 9568 2421 9571
rect 2372 9540 2421 9568
rect 2372 9528 2378 9540
rect 2409 9537 2421 9540
rect 2455 9537 2467 9571
rect 2409 9531 2467 9537
rect 2590 9528 2596 9580
rect 2648 9568 2654 9580
rect 3053 9571 3111 9577
rect 3053 9568 3065 9571
rect 2648 9540 3065 9568
rect 2648 9528 2654 9540
rect 3053 9537 3065 9540
rect 3099 9537 3111 9571
rect 3053 9531 3111 9537
rect 3234 9528 3240 9580
rect 3292 9528 3298 9580
rect 3881 9571 3939 9577
rect 3881 9537 3893 9571
rect 3927 9568 3939 9571
rect 4706 9568 4712 9580
rect 3927 9540 4712 9568
rect 3927 9537 3939 9540
rect 3881 9531 3939 9537
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 4982 9528 4988 9580
rect 5040 9568 5046 9580
rect 5077 9571 5135 9577
rect 5077 9568 5089 9571
rect 5040 9540 5089 9568
rect 5040 9528 5046 9540
rect 5077 9537 5089 9540
rect 5123 9537 5135 9571
rect 5077 9531 5135 9537
rect 5258 9528 5264 9580
rect 5316 9528 5322 9580
rect 5399 9571 5457 9577
rect 5399 9537 5411 9571
rect 5445 9568 5457 9571
rect 5902 9568 5908 9580
rect 5445 9540 5908 9568
rect 5445 9537 5457 9540
rect 5399 9531 5457 9537
rect 5902 9528 5908 9540
rect 5960 9528 5966 9580
rect 7098 9528 7104 9580
rect 7156 9568 7162 9580
rect 7208 9577 7236 9676
rect 7484 9636 7512 9676
rect 8205 9673 8217 9707
rect 8251 9704 8263 9707
rect 8478 9704 8484 9716
rect 8251 9676 8484 9704
rect 8251 9673 8263 9676
rect 8205 9667 8263 9673
rect 8478 9664 8484 9676
rect 8536 9664 8542 9716
rect 9398 9664 9404 9716
rect 9456 9664 9462 9716
rect 11238 9664 11244 9716
rect 11296 9704 11302 9716
rect 11514 9704 11520 9716
rect 11296 9676 11520 9704
rect 11296 9664 11302 9676
rect 11514 9664 11520 9676
rect 11572 9704 11578 9716
rect 13262 9704 13268 9716
rect 11572 9676 13268 9704
rect 11572 9664 11578 9676
rect 13262 9664 13268 9676
rect 13320 9664 13326 9716
rect 14182 9664 14188 9716
rect 14240 9704 14246 9716
rect 14277 9707 14335 9713
rect 14277 9704 14289 9707
rect 14240 9676 14289 9704
rect 14240 9664 14246 9676
rect 14277 9673 14289 9676
rect 14323 9673 14335 9707
rect 21082 9704 21088 9716
rect 14277 9667 14335 9673
rect 17604 9676 21088 9704
rect 8297 9639 8355 9645
rect 8297 9636 8309 9639
rect 7484 9608 8309 9636
rect 8297 9605 8309 9608
rect 8343 9636 8355 9639
rect 9416 9636 9444 9664
rect 8343 9608 9168 9636
rect 9416 9608 10916 9636
rect 8343 9605 8355 9608
rect 8297 9599 8355 9605
rect 7193 9571 7251 9577
rect 7193 9568 7205 9571
rect 7156 9540 7205 9568
rect 7156 9528 7162 9540
rect 7193 9537 7205 9540
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 5537 9503 5595 9509
rect 5537 9469 5549 9503
rect 5583 9500 5595 9503
rect 5718 9500 5724 9512
rect 5583 9472 5724 9500
rect 5583 9469 5595 9472
rect 5537 9463 5595 9469
rect 5718 9460 5724 9472
rect 5776 9460 5782 9512
rect 4154 9392 4160 9444
rect 4212 9432 4218 9444
rect 7006 9432 7012 9444
rect 4212 9404 7012 9432
rect 4212 9392 4218 9404
rect 7006 9392 7012 9404
rect 7064 9392 7070 9444
rect 7300 9432 7328 9531
rect 7374 9528 7380 9580
rect 7432 9577 7438 9580
rect 9140 9577 9168 9608
rect 7432 9571 7471 9577
rect 7459 9537 7471 9571
rect 7432 9531 7471 9537
rect 9125 9571 9183 9577
rect 9125 9537 9137 9571
rect 9171 9537 9183 9571
rect 9125 9531 9183 9537
rect 7432 9528 7438 9531
rect 9306 9528 9312 9580
rect 9364 9528 9370 9580
rect 9401 9571 9459 9577
rect 9401 9537 9413 9571
rect 9447 9537 9459 9571
rect 9401 9531 9459 9537
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9537 9551 9571
rect 9493 9531 9551 9537
rect 7650 9460 7656 9512
rect 7708 9500 7714 9512
rect 8021 9503 8079 9509
rect 8021 9500 8033 9503
rect 7708 9472 8033 9500
rect 7708 9460 7714 9472
rect 8021 9469 8033 9472
rect 8067 9469 8079 9503
rect 9416 9500 9444 9531
rect 8021 9463 8079 9469
rect 8128 9472 9444 9500
rect 8128 9444 8156 9472
rect 8110 9432 8116 9444
rect 7300 9404 8116 9432
rect 8110 9392 8116 9404
rect 8168 9392 8174 9444
rect 8665 9435 8723 9441
rect 8665 9401 8677 9435
rect 8711 9432 8723 9435
rect 8846 9432 8852 9444
rect 8711 9404 8852 9432
rect 8711 9401 8723 9404
rect 8665 9395 8723 9401
rect 8846 9392 8852 9404
rect 8904 9392 8910 9444
rect 8938 9392 8944 9444
rect 8996 9432 9002 9444
rect 9306 9432 9312 9444
rect 8996 9404 9312 9432
rect 8996 9392 9002 9404
rect 9306 9392 9312 9404
rect 9364 9432 9370 9444
rect 9508 9432 9536 9531
rect 9858 9528 9864 9580
rect 9916 9568 9922 9580
rect 10229 9571 10287 9577
rect 10229 9568 10241 9571
rect 9916 9540 10241 9568
rect 9916 9528 9922 9540
rect 10229 9537 10241 9540
rect 10275 9537 10287 9571
rect 10229 9531 10287 9537
rect 9766 9460 9772 9512
rect 9824 9460 9830 9512
rect 10318 9460 10324 9512
rect 10376 9460 10382 9512
rect 10502 9432 10508 9444
rect 9364 9404 9536 9432
rect 10336 9404 10508 9432
rect 9364 9392 9370 9404
rect 1670 9324 1676 9376
rect 1728 9324 1734 9376
rect 2593 9367 2651 9373
rect 2593 9333 2605 9367
rect 2639 9364 2651 9367
rect 2958 9364 2964 9376
rect 2639 9336 2964 9364
rect 2639 9333 2651 9336
rect 2593 9327 2651 9333
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 3326 9324 3332 9376
rect 3384 9364 3390 9376
rect 4341 9367 4399 9373
rect 4341 9364 4353 9367
rect 3384 9336 4353 9364
rect 3384 9324 3390 9336
rect 4341 9333 4353 9336
rect 4387 9364 4399 9367
rect 4890 9364 4896 9376
rect 4387 9336 4896 9364
rect 4387 9333 4399 9336
rect 4341 9327 4399 9333
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 5350 9324 5356 9376
rect 5408 9364 5414 9376
rect 7742 9364 7748 9376
rect 5408 9336 7748 9364
rect 5408 9324 5414 9336
rect 7742 9324 7748 9336
rect 7800 9324 7806 9376
rect 7926 9324 7932 9376
rect 7984 9364 7990 9376
rect 10226 9364 10232 9376
rect 7984 9336 10232 9364
rect 7984 9324 7990 9336
rect 10226 9324 10232 9336
rect 10284 9324 10290 9376
rect 10336 9373 10364 9404
rect 10502 9392 10508 9404
rect 10560 9392 10566 9444
rect 10888 9432 10916 9608
rect 11054 9596 11060 9648
rect 11112 9636 11118 9648
rect 11112 9608 11928 9636
rect 11112 9596 11118 9608
rect 10962 9528 10968 9580
rect 11020 9568 11026 9580
rect 11900 9577 11928 9608
rect 12710 9596 12716 9648
rect 12768 9636 12774 9648
rect 12768 9608 12940 9636
rect 12768 9596 12774 9608
rect 12912 9577 12940 9608
rect 13722 9596 13728 9648
rect 13780 9596 13786 9648
rect 13814 9596 13820 9648
rect 13872 9636 13878 9648
rect 14918 9636 14924 9648
rect 13872 9608 14924 9636
rect 13872 9596 13878 9608
rect 11701 9571 11759 9577
rect 11701 9568 11713 9571
rect 11020 9540 11713 9568
rect 11020 9528 11026 9540
rect 11701 9537 11713 9540
rect 11747 9537 11759 9571
rect 11701 9531 11759 9537
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 12897 9571 12955 9577
rect 12897 9537 12909 9571
rect 12943 9537 12955 9571
rect 12897 9531 12955 9537
rect 13081 9571 13139 9577
rect 13081 9537 13093 9571
rect 13127 9537 13139 9571
rect 13081 9531 13139 9537
rect 13265 9571 13323 9577
rect 13265 9537 13277 9571
rect 13311 9568 13323 9571
rect 13906 9568 13912 9580
rect 13311 9540 13912 9568
rect 13311 9537 13323 9540
rect 13265 9531 13323 9537
rect 13096 9500 13124 9531
rect 13906 9528 13912 9540
rect 13964 9528 13970 9580
rect 14292 9577 14320 9608
rect 14918 9596 14924 9608
rect 14976 9596 14982 9648
rect 15933 9639 15991 9645
rect 15933 9605 15945 9639
rect 15979 9636 15991 9639
rect 16298 9636 16304 9648
rect 15979 9608 16304 9636
rect 15979 9605 15991 9608
rect 15933 9599 15991 9605
rect 16298 9596 16304 9608
rect 16356 9596 16362 9648
rect 17218 9596 17224 9648
rect 17276 9636 17282 9648
rect 17604 9645 17632 9676
rect 21082 9664 21088 9676
rect 21140 9664 21146 9716
rect 22094 9664 22100 9716
rect 22152 9664 22158 9716
rect 17589 9639 17647 9645
rect 17589 9636 17601 9639
rect 17276 9608 17601 9636
rect 17276 9596 17282 9608
rect 17589 9605 17601 9608
rect 17635 9605 17647 9639
rect 17589 9599 17647 9605
rect 17678 9596 17684 9648
rect 17736 9636 17742 9648
rect 18049 9639 18107 9645
rect 18049 9636 18061 9639
rect 17736 9608 18061 9636
rect 17736 9596 17742 9608
rect 18049 9605 18061 9608
rect 18095 9636 18107 9639
rect 20349 9639 20407 9645
rect 18095 9608 19104 9636
rect 18095 9605 18107 9608
rect 18049 9599 18107 9605
rect 14277 9571 14335 9577
rect 14277 9537 14289 9571
rect 14323 9537 14335 9571
rect 14277 9531 14335 9537
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9568 14519 9571
rect 14734 9568 14740 9580
rect 14507 9540 14740 9568
rect 14507 9537 14519 9540
rect 14461 9531 14519 9537
rect 14734 9528 14740 9540
rect 14792 9568 14798 9580
rect 15013 9571 15071 9577
rect 15013 9568 15025 9571
rect 14792 9540 15025 9568
rect 14792 9528 14798 9540
rect 15013 9537 15025 9540
rect 15059 9537 15071 9571
rect 15013 9531 15071 9537
rect 15102 9528 15108 9580
rect 15160 9528 15166 9580
rect 16758 9528 16764 9580
rect 16816 9568 16822 9580
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16816 9540 16865 9568
rect 16816 9528 16822 9540
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 18233 9571 18291 9577
rect 18233 9537 18245 9571
rect 18279 9537 18291 9571
rect 18233 9531 18291 9537
rect 13354 9500 13360 9512
rect 13096 9472 13360 9500
rect 13354 9460 13360 9472
rect 13412 9460 13418 9512
rect 13924 9500 13952 9528
rect 13924 9472 15332 9500
rect 14458 9432 14464 9444
rect 10888 9404 14464 9432
rect 14458 9392 14464 9404
rect 14516 9392 14522 9444
rect 10321 9367 10379 9373
rect 10321 9333 10333 9367
rect 10367 9333 10379 9367
rect 10321 9327 10379 9333
rect 10597 9367 10655 9373
rect 10597 9333 10609 9367
rect 10643 9364 10655 9367
rect 10870 9364 10876 9376
rect 10643 9336 10876 9364
rect 10643 9333 10655 9336
rect 10597 9327 10655 9333
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 11793 9367 11851 9373
rect 11793 9333 11805 9367
rect 11839 9364 11851 9367
rect 12526 9364 12532 9376
rect 11839 9336 12532 9364
rect 11839 9333 11851 9336
rect 11793 9327 11851 9333
rect 12526 9324 12532 9336
rect 12584 9324 12590 9376
rect 14826 9324 14832 9376
rect 14884 9364 14890 9376
rect 15013 9367 15071 9373
rect 15013 9364 15025 9367
rect 14884 9336 15025 9364
rect 14884 9324 14890 9336
rect 15013 9333 15025 9336
rect 15059 9333 15071 9367
rect 15304 9364 15332 9472
rect 16022 9460 16028 9512
rect 16080 9500 16086 9512
rect 16390 9500 16396 9512
rect 16080 9472 16396 9500
rect 16080 9460 16086 9472
rect 16390 9460 16396 9472
rect 16448 9500 16454 9512
rect 17221 9503 17279 9509
rect 17221 9500 17233 9503
rect 16448 9472 17233 9500
rect 16448 9460 16454 9472
rect 17221 9469 17233 9472
rect 17267 9469 17279 9503
rect 18248 9500 18276 9531
rect 18414 9528 18420 9580
rect 18472 9528 18478 9580
rect 19076 9577 19104 9608
rect 20349 9605 20361 9639
rect 20395 9636 20407 9639
rect 21174 9636 21180 9648
rect 20395 9608 21180 9636
rect 20395 9605 20407 9608
rect 20349 9599 20407 9605
rect 21174 9596 21180 9608
rect 21232 9596 21238 9648
rect 21266 9596 21272 9648
rect 21324 9636 21330 9648
rect 21542 9636 21548 9648
rect 21324 9608 21548 9636
rect 21324 9596 21330 9608
rect 21542 9596 21548 9608
rect 21600 9596 21606 9648
rect 22112 9636 22140 9664
rect 22112 9608 22324 9636
rect 19061 9571 19119 9577
rect 19061 9537 19073 9571
rect 19107 9537 19119 9571
rect 19061 9531 19119 9537
rect 19334 9528 19340 9580
rect 19392 9528 19398 9580
rect 20073 9571 20131 9577
rect 20073 9537 20085 9571
rect 20119 9537 20131 9571
rect 20073 9531 20131 9537
rect 20257 9571 20315 9577
rect 20257 9537 20269 9571
rect 20303 9568 20315 9571
rect 20622 9568 20628 9580
rect 20303 9540 20628 9568
rect 20303 9537 20315 9540
rect 20257 9531 20315 9537
rect 18322 9500 18328 9512
rect 18248 9472 18328 9500
rect 17221 9463 17279 9469
rect 18322 9460 18328 9472
rect 18380 9500 18386 9512
rect 18874 9500 18880 9512
rect 18380 9472 18880 9500
rect 18380 9460 18386 9472
rect 18874 9460 18880 9472
rect 18932 9460 18938 9512
rect 19153 9503 19211 9509
rect 19153 9469 19165 9503
rect 19199 9500 19211 9503
rect 19242 9500 19248 9512
rect 19199 9472 19248 9500
rect 19199 9469 19211 9472
rect 19153 9463 19211 9469
rect 19242 9460 19248 9472
rect 19300 9500 19306 9512
rect 20088 9500 20116 9531
rect 20622 9528 20628 9540
rect 20680 9528 20686 9580
rect 20806 9528 20812 9580
rect 20864 9568 20870 9580
rect 21726 9568 21732 9580
rect 20864 9540 21732 9568
rect 20864 9528 20870 9540
rect 21726 9528 21732 9540
rect 21784 9528 21790 9580
rect 22002 9528 22008 9580
rect 22060 9528 22066 9580
rect 22296 9577 22324 9608
rect 22097 9571 22155 9577
rect 22097 9537 22109 9571
rect 22143 9537 22155 9571
rect 22097 9531 22155 9537
rect 22281 9571 22339 9577
rect 22281 9537 22293 9571
rect 22327 9537 22339 9571
rect 22281 9531 22339 9537
rect 20438 9500 20444 9512
rect 19300 9472 20444 9500
rect 19300 9460 19306 9472
rect 20438 9460 20444 9472
rect 20496 9460 20502 9512
rect 21174 9460 21180 9512
rect 21232 9500 21238 9512
rect 22112 9500 22140 9531
rect 21232 9472 22140 9500
rect 21232 9460 21238 9472
rect 15381 9435 15439 9441
rect 15381 9401 15393 9435
rect 15427 9432 15439 9435
rect 19521 9435 19579 9441
rect 15427 9404 17264 9432
rect 15427 9401 15439 9404
rect 15381 9395 15439 9401
rect 17236 9376 17264 9404
rect 19521 9401 19533 9435
rect 19567 9432 19579 9435
rect 22278 9432 22284 9444
rect 19567 9404 22284 9432
rect 19567 9401 19579 9404
rect 19521 9395 19579 9401
rect 22278 9392 22284 9404
rect 22336 9392 22342 9444
rect 16850 9364 16856 9376
rect 15304 9336 16856 9364
rect 15013 9327 15071 9333
rect 16850 9324 16856 9336
rect 16908 9364 16914 9376
rect 16991 9367 17049 9373
rect 16991 9364 17003 9367
rect 16908 9336 17003 9364
rect 16908 9324 16914 9336
rect 16991 9333 17003 9336
rect 17037 9333 17049 9367
rect 16991 9327 17049 9333
rect 17126 9324 17132 9376
rect 17184 9324 17190 9376
rect 17218 9324 17224 9376
rect 17276 9324 17282 9376
rect 18598 9324 18604 9376
rect 18656 9364 18662 9376
rect 19426 9364 19432 9376
rect 18656 9336 19432 9364
rect 18656 9324 18662 9336
rect 19426 9324 19432 9336
rect 19484 9364 19490 9376
rect 21634 9364 21640 9376
rect 19484 9336 21640 9364
rect 19484 9324 19490 9336
rect 21634 9324 21640 9336
rect 21692 9324 21698 9376
rect 22094 9324 22100 9376
rect 22152 9364 22158 9376
rect 22370 9364 22376 9376
rect 22152 9336 22376 9364
rect 22152 9324 22158 9336
rect 22370 9324 22376 9336
rect 22428 9324 22434 9376
rect 22465 9367 22523 9373
rect 22465 9333 22477 9367
rect 22511 9364 22523 9367
rect 22646 9364 22652 9376
rect 22511 9336 22652 9364
rect 22511 9333 22523 9336
rect 22465 9327 22523 9333
rect 22646 9324 22652 9336
rect 22704 9324 22710 9376
rect 1104 9274 23828 9296
rect 1104 9222 3790 9274
rect 3842 9222 3854 9274
rect 3906 9222 3918 9274
rect 3970 9222 3982 9274
rect 4034 9222 4046 9274
rect 4098 9222 9471 9274
rect 9523 9222 9535 9274
rect 9587 9222 9599 9274
rect 9651 9222 9663 9274
rect 9715 9222 9727 9274
rect 9779 9222 15152 9274
rect 15204 9222 15216 9274
rect 15268 9222 15280 9274
rect 15332 9222 15344 9274
rect 15396 9222 15408 9274
rect 15460 9222 20833 9274
rect 20885 9222 20897 9274
rect 20949 9222 20961 9274
rect 21013 9222 21025 9274
rect 21077 9222 21089 9274
rect 21141 9222 23828 9274
rect 1104 9200 23828 9222
rect 5166 9120 5172 9172
rect 5224 9120 5230 9172
rect 5350 9120 5356 9172
rect 5408 9120 5414 9172
rect 6822 9120 6828 9172
rect 6880 9120 6886 9172
rect 7009 9163 7067 9169
rect 7009 9129 7021 9163
rect 7055 9160 7067 9163
rect 7190 9160 7196 9172
rect 7055 9132 7196 9160
rect 7055 9129 7067 9132
rect 7009 9123 7067 9129
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 9214 9120 9220 9172
rect 9272 9160 9278 9172
rect 9272 9132 14228 9160
rect 9272 9120 9278 9132
rect 4522 9052 4528 9104
rect 4580 9092 4586 9104
rect 5261 9095 5319 9101
rect 5261 9092 5273 9095
rect 4580 9064 5273 9092
rect 4580 9052 4586 9064
rect 5261 9061 5273 9064
rect 5307 9061 5319 9095
rect 5261 9055 5319 9061
rect 2222 9024 2228 9036
rect 1872 8996 2228 9024
rect 1872 8965 1900 8996
rect 2222 8984 2228 8996
rect 2280 8984 2286 9036
rect 2406 8984 2412 9036
rect 2464 9024 2470 9036
rect 2464 8996 4016 9024
rect 2464 8984 2470 8996
rect 1857 8959 1915 8965
rect 1857 8925 1869 8959
rect 1903 8925 1915 8959
rect 1857 8919 1915 8925
rect 2041 8959 2099 8965
rect 2041 8925 2053 8959
rect 2087 8956 2099 8959
rect 2130 8956 2136 8968
rect 2087 8928 2136 8956
rect 2087 8925 2099 8928
rect 2041 8919 2099 8925
rect 2130 8916 2136 8928
rect 2188 8956 2194 8968
rect 2188 8928 2820 8956
rect 2188 8916 2194 8928
rect 2498 8848 2504 8900
rect 2556 8888 2562 8900
rect 2685 8891 2743 8897
rect 2685 8888 2697 8891
rect 2556 8860 2697 8888
rect 2556 8848 2562 8860
rect 2685 8857 2697 8860
rect 2731 8857 2743 8891
rect 2792 8888 2820 8928
rect 2866 8916 2872 8968
rect 2924 8956 2930 8968
rect 3988 8965 4016 8996
rect 5166 8984 5172 9036
rect 5224 9024 5230 9036
rect 5368 9024 5396 9120
rect 6840 9092 6868 9120
rect 11517 9095 11575 9101
rect 11517 9092 11529 9095
rect 6840 9064 11529 9092
rect 11517 9061 11529 9064
rect 11563 9061 11575 9095
rect 13998 9092 14004 9104
rect 11517 9055 11575 9061
rect 13188 9064 14004 9092
rect 5224 8996 5396 9024
rect 5224 8984 5230 8996
rect 6178 8984 6184 9036
rect 6236 9024 6242 9036
rect 6733 9027 6791 9033
rect 6733 9024 6745 9027
rect 6236 8996 6745 9024
rect 6236 8984 6242 8996
rect 6733 8993 6745 8996
rect 6779 8993 6791 9027
rect 6733 8987 6791 8993
rect 6822 8984 6828 9036
rect 6880 9024 6886 9036
rect 7650 9024 7656 9036
rect 6880 8996 7656 9024
rect 6880 8984 6886 8996
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 7834 8984 7840 9036
rect 7892 9024 7898 9036
rect 10318 9024 10324 9036
rect 7892 8996 10324 9024
rect 7892 8984 7898 8996
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 10594 8984 10600 9036
rect 10652 9024 10658 9036
rect 11057 9027 11115 9033
rect 11057 9024 11069 9027
rect 10652 8996 11069 9024
rect 10652 8984 10658 8996
rect 11057 8993 11069 8996
rect 11103 9024 11115 9027
rect 12158 9024 12164 9036
rect 11103 8996 12164 9024
rect 11103 8993 11115 8996
rect 11057 8987 11115 8993
rect 2961 8959 3019 8965
rect 2961 8956 2973 8959
rect 2924 8928 2973 8956
rect 2924 8916 2930 8928
rect 2961 8925 2973 8928
rect 3007 8925 3019 8959
rect 2961 8919 3019 8925
rect 3973 8959 4031 8965
rect 3973 8925 3985 8959
rect 4019 8925 4031 8959
rect 3973 8919 4031 8925
rect 5353 8959 5411 8965
rect 5353 8925 5365 8959
rect 5399 8956 5411 8959
rect 6454 8956 6460 8968
rect 5399 8928 6460 8956
rect 5399 8925 5411 8928
rect 5353 8919 5411 8925
rect 6454 8916 6460 8928
rect 6512 8916 6518 8968
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8925 6607 8959
rect 6549 8919 6607 8925
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8956 6699 8959
rect 7006 8956 7012 8968
rect 6687 8928 7012 8956
rect 6687 8925 6699 8928
rect 6641 8919 6699 8925
rect 4154 8888 4160 8900
rect 2792 8860 4160 8888
rect 2685 8851 2743 8857
rect 4154 8848 4160 8860
rect 4212 8848 4218 8900
rect 4246 8848 4252 8900
rect 4304 8848 4310 8900
rect 5074 8848 5080 8900
rect 5132 8848 5138 8900
rect 5258 8848 5264 8900
rect 5316 8888 5322 8900
rect 5442 8888 5448 8900
rect 5316 8860 5448 8888
rect 5316 8848 5322 8860
rect 5442 8848 5448 8860
rect 5500 8888 5506 8900
rect 6564 8888 6592 8919
rect 7006 8916 7012 8928
rect 7064 8916 7070 8968
rect 9122 8916 9128 8968
rect 9180 8916 9186 8968
rect 10042 8916 10048 8968
rect 10100 8916 10106 8968
rect 8018 8888 8024 8900
rect 5500 8860 8024 8888
rect 5500 8848 5506 8860
rect 8018 8848 8024 8860
rect 8076 8848 8082 8900
rect 9582 8848 9588 8900
rect 9640 8848 9646 8900
rect 10336 8888 10364 8984
rect 11698 8916 11704 8968
rect 11756 8916 11762 8968
rect 11808 8965 11836 8996
rect 12158 8984 12164 8996
rect 12216 8984 12222 9036
rect 11793 8959 11851 8965
rect 11793 8925 11805 8959
rect 11839 8925 11851 8959
rect 11793 8919 11851 8925
rect 11974 8916 11980 8968
rect 12032 8916 12038 8968
rect 12069 8959 12127 8965
rect 12069 8925 12081 8959
rect 12115 8925 12127 8959
rect 12069 8919 12127 8925
rect 12084 8888 12112 8919
rect 12526 8916 12532 8968
rect 12584 8916 12590 8968
rect 13188 8965 13216 9064
rect 13998 9052 14004 9064
rect 14056 9052 14062 9104
rect 14200 9092 14228 9132
rect 17862 9120 17868 9172
rect 17920 9160 17926 9172
rect 20073 9163 20131 9169
rect 20073 9160 20085 9163
rect 17920 9132 20085 9160
rect 17920 9120 17926 9132
rect 20073 9129 20085 9132
rect 20119 9129 20131 9163
rect 20990 9160 20996 9172
rect 20073 9123 20131 9129
rect 20180 9132 20996 9160
rect 15562 9092 15568 9104
rect 14200 9064 15568 9092
rect 15562 9052 15568 9064
rect 15620 9052 15626 9104
rect 18598 9092 18604 9104
rect 16592 9064 18604 9092
rect 13354 8984 13360 9036
rect 13412 9024 13418 9036
rect 14366 9024 14372 9036
rect 13412 8996 14372 9024
rect 13412 8984 13418 8996
rect 14366 8984 14372 8996
rect 14424 8984 14430 9036
rect 14550 8984 14556 9036
rect 14608 9024 14614 9036
rect 14826 9024 14832 9036
rect 14608 8996 14832 9024
rect 14608 8984 14614 8996
rect 14826 8984 14832 8996
rect 14884 8984 14890 9036
rect 15473 9027 15531 9033
rect 15473 8993 15485 9027
rect 15519 9024 15531 9027
rect 16482 9024 16488 9036
rect 15519 8996 16488 9024
rect 15519 8993 15531 8996
rect 15473 8987 15531 8993
rect 16482 8984 16488 8996
rect 16540 8984 16546 9036
rect 13173 8959 13231 8965
rect 13173 8925 13185 8959
rect 13219 8925 13231 8959
rect 13173 8919 13231 8925
rect 13262 8916 13268 8968
rect 13320 8916 13326 8968
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8925 13507 8959
rect 13449 8919 13507 8925
rect 13541 8959 13599 8965
rect 13541 8925 13553 8959
rect 13587 8956 13599 8959
rect 13814 8956 13820 8968
rect 13587 8928 13820 8956
rect 13587 8925 13599 8928
rect 13541 8919 13599 8925
rect 12802 8888 12808 8900
rect 10336 8860 12808 8888
rect 12802 8848 12808 8860
rect 12860 8848 12866 8900
rect 13464 8888 13492 8919
rect 13814 8916 13820 8928
rect 13872 8956 13878 8968
rect 14274 8956 14280 8968
rect 13872 8928 14280 8956
rect 13872 8916 13878 8928
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 14458 8916 14464 8968
rect 14516 8916 14522 8968
rect 14734 8916 14740 8968
rect 14792 8916 14798 8968
rect 14918 8916 14924 8968
rect 14976 8956 14982 8968
rect 14976 8928 15976 8956
rect 14976 8916 14982 8928
rect 14752 8888 14780 8916
rect 13464 8860 14780 8888
rect 15948 8888 15976 8928
rect 16022 8916 16028 8968
rect 16080 8956 16086 8968
rect 16592 8965 16620 9064
rect 18598 9052 18604 9064
rect 18656 9052 18662 9104
rect 18785 9095 18843 9101
rect 18785 9061 18797 9095
rect 18831 9092 18843 9095
rect 19150 9092 19156 9104
rect 18831 9064 19156 9092
rect 18831 9061 18843 9064
rect 18785 9055 18843 9061
rect 19150 9052 19156 9064
rect 19208 9052 19214 9104
rect 19521 9095 19579 9101
rect 19521 9061 19533 9095
rect 19567 9092 19579 9095
rect 19610 9092 19616 9104
rect 19567 9064 19616 9092
rect 19567 9061 19579 9064
rect 19521 9055 19579 9061
rect 19610 9052 19616 9064
rect 19668 9052 19674 9104
rect 16850 8984 16856 9036
rect 16908 8984 16914 9036
rect 17586 8984 17592 9036
rect 17644 9024 17650 9036
rect 20180 9024 20208 9132
rect 20990 9120 20996 9132
rect 21048 9160 21054 9172
rect 22097 9163 22155 9169
rect 21048 9132 21404 9160
rect 21048 9120 21054 9132
rect 20530 9052 20536 9104
rect 20588 9092 20594 9104
rect 21082 9092 21088 9104
rect 20588 9064 21088 9092
rect 20588 9052 20594 9064
rect 21082 9052 21088 9064
rect 21140 9052 21146 9104
rect 20806 9024 20812 9036
rect 17644 8996 20208 9024
rect 20364 8996 20812 9024
rect 17644 8984 17650 8996
rect 16577 8959 16635 8965
rect 16577 8956 16589 8959
rect 16080 8928 16589 8956
rect 16080 8916 16086 8928
rect 16577 8925 16589 8928
rect 16623 8925 16635 8959
rect 16868 8956 16896 8984
rect 18046 8956 18052 8968
rect 16868 8928 18052 8956
rect 16577 8919 16635 8925
rect 18046 8916 18052 8928
rect 18104 8916 18110 8968
rect 18141 8959 18199 8965
rect 18141 8925 18153 8959
rect 18187 8956 18199 8959
rect 18690 8956 18696 8968
rect 18187 8928 18696 8956
rect 18187 8925 18199 8928
rect 18141 8919 18199 8925
rect 18690 8916 18696 8928
rect 18748 8916 18754 8968
rect 20364 8965 20392 8996
rect 20806 8984 20812 8996
rect 20864 9024 20870 9036
rect 21266 9024 21272 9036
rect 20864 8996 21272 9024
rect 20864 8984 20870 8996
rect 21266 8984 21272 8996
rect 21324 8984 21330 9036
rect 21376 9024 21404 9132
rect 22097 9129 22109 9163
rect 22143 9160 22155 9163
rect 22186 9160 22192 9172
rect 22143 9132 22192 9160
rect 22143 9129 22155 9132
rect 22097 9123 22155 9129
rect 22186 9120 22192 9132
rect 22244 9120 22250 9172
rect 22830 9160 22836 9172
rect 22480 9132 22836 9160
rect 21818 9024 21824 9036
rect 21376 8996 21824 9024
rect 20257 8959 20315 8965
rect 20257 8925 20269 8959
rect 20303 8925 20315 8959
rect 20257 8919 20315 8925
rect 20349 8959 20407 8965
rect 20349 8925 20361 8959
rect 20395 8925 20407 8959
rect 20349 8919 20407 8925
rect 15948 8860 16068 8888
rect 1949 8823 2007 8829
rect 1949 8789 1961 8823
rect 1995 8820 2007 8823
rect 3050 8820 3056 8832
rect 1995 8792 3056 8820
rect 1995 8789 2007 8792
rect 1949 8783 2007 8789
rect 3050 8780 3056 8792
rect 3108 8780 3114 8832
rect 3694 8780 3700 8832
rect 3752 8820 3758 8832
rect 4062 8820 4068 8832
rect 3752 8792 4068 8820
rect 3752 8780 3758 8792
rect 4062 8780 4068 8792
rect 4120 8820 4126 8832
rect 10594 8820 10600 8832
rect 4120 8792 10600 8820
rect 4120 8780 4126 8792
rect 10594 8780 10600 8792
rect 10652 8780 10658 8832
rect 11330 8780 11336 8832
rect 11388 8820 11394 8832
rect 12621 8823 12679 8829
rect 12621 8820 12633 8823
rect 11388 8792 12633 8820
rect 11388 8780 11394 8792
rect 12621 8789 12633 8792
rect 12667 8789 12679 8823
rect 12621 8783 12679 8789
rect 13725 8823 13783 8829
rect 13725 8789 13737 8823
rect 13771 8820 13783 8823
rect 15654 8820 15660 8832
rect 13771 8792 15660 8820
rect 13771 8789 13783 8792
rect 13725 8783 13783 8789
rect 15654 8780 15660 8792
rect 15712 8780 15718 8832
rect 16040 8829 16068 8860
rect 18322 8848 18328 8900
rect 18380 8888 18386 8900
rect 19794 8888 19800 8900
rect 18380 8860 19800 8888
rect 18380 8848 18386 8860
rect 19794 8848 19800 8860
rect 19852 8848 19858 8900
rect 20272 8888 20300 8919
rect 20530 8916 20536 8968
rect 20588 8916 20594 8968
rect 20625 8959 20683 8965
rect 20625 8925 20637 8959
rect 20671 8956 20683 8959
rect 21082 8956 21088 8968
rect 20671 8928 21088 8956
rect 20671 8925 20683 8928
rect 20625 8919 20683 8925
rect 21082 8916 21088 8928
rect 21140 8956 21146 8968
rect 21376 8965 21404 8996
rect 21818 8984 21824 8996
rect 21876 8984 21882 9036
rect 22480 8968 22508 9132
rect 22830 9120 22836 9132
rect 22888 9120 22894 9172
rect 22738 9052 22744 9104
rect 22796 9092 22802 9104
rect 23201 9095 23259 9101
rect 23201 9092 23213 9095
rect 22796 9064 23213 9092
rect 22796 9052 22802 9064
rect 23201 9061 23213 9064
rect 23247 9061 23259 9095
rect 23201 9055 23259 9061
rect 22756 9024 22784 9052
rect 22572 8996 22784 9024
rect 21177 8959 21235 8965
rect 21177 8956 21189 8959
rect 21140 8928 21189 8956
rect 21140 8916 21146 8928
rect 21177 8925 21189 8928
rect 21223 8925 21235 8959
rect 21177 8919 21235 8925
rect 21361 8959 21419 8965
rect 21361 8925 21373 8959
rect 21407 8925 21419 8959
rect 21361 8919 21419 8925
rect 21450 8916 21456 8968
rect 21508 8916 21514 8968
rect 22373 8959 22431 8965
rect 22373 8925 22385 8959
rect 22419 8925 22431 8959
rect 22373 8919 22431 8925
rect 22388 8888 22416 8919
rect 22462 8916 22468 8968
rect 22520 8916 22526 8968
rect 22572 8965 22600 8996
rect 22557 8959 22615 8965
rect 22557 8925 22569 8959
rect 22603 8925 22615 8959
rect 22557 8919 22615 8925
rect 22741 8959 22799 8965
rect 22741 8925 22753 8959
rect 22787 8956 22799 8959
rect 23198 8956 23204 8968
rect 22787 8928 23204 8956
rect 22787 8925 22799 8928
rect 22741 8919 22799 8925
rect 23198 8916 23204 8928
rect 23256 8916 23262 8968
rect 22830 8888 22836 8900
rect 20272 8860 22836 8888
rect 22830 8848 22836 8860
rect 22888 8848 22894 8900
rect 16025 8823 16083 8829
rect 16025 8789 16037 8823
rect 16071 8820 16083 8823
rect 16942 8820 16948 8832
rect 16071 8792 16948 8820
rect 16071 8789 16083 8792
rect 16025 8783 16083 8789
rect 16942 8780 16948 8792
rect 17000 8780 17006 8832
rect 17862 8780 17868 8832
rect 17920 8780 17926 8832
rect 18046 8780 18052 8832
rect 18104 8820 18110 8832
rect 21358 8820 21364 8832
rect 18104 8792 21364 8820
rect 18104 8780 18110 8792
rect 21358 8780 21364 8792
rect 21416 8780 21422 8832
rect 21634 8780 21640 8832
rect 21692 8780 21698 8832
rect 1104 8730 23987 8752
rect 1104 8678 6630 8730
rect 6682 8678 6694 8730
rect 6746 8678 6758 8730
rect 6810 8678 6822 8730
rect 6874 8678 6886 8730
rect 6938 8678 12311 8730
rect 12363 8678 12375 8730
rect 12427 8678 12439 8730
rect 12491 8678 12503 8730
rect 12555 8678 12567 8730
rect 12619 8678 17992 8730
rect 18044 8678 18056 8730
rect 18108 8678 18120 8730
rect 18172 8678 18184 8730
rect 18236 8678 18248 8730
rect 18300 8678 23673 8730
rect 23725 8678 23737 8730
rect 23789 8678 23801 8730
rect 23853 8678 23865 8730
rect 23917 8678 23929 8730
rect 23981 8678 23987 8730
rect 1104 8656 23987 8678
rect 3513 8619 3571 8625
rect 3513 8585 3525 8619
rect 3559 8616 3571 8619
rect 7098 8616 7104 8628
rect 3559 8588 7104 8616
rect 3559 8585 3571 8588
rect 3513 8579 3571 8585
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 9309 8619 9367 8625
rect 9309 8616 9321 8619
rect 7800 8588 9321 8616
rect 7800 8576 7806 8588
rect 9309 8585 9321 8588
rect 9355 8585 9367 8619
rect 9309 8579 9367 8585
rect 2746 8520 3372 8548
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8480 2467 8483
rect 2590 8480 2596 8492
rect 2455 8452 2596 8480
rect 2455 8449 2467 8452
rect 2409 8443 2467 8449
rect 2332 8412 2360 8443
rect 2590 8440 2596 8452
rect 2648 8480 2654 8492
rect 2746 8480 2774 8520
rect 2648 8452 2774 8480
rect 2648 8440 2654 8452
rect 2958 8440 2964 8492
rect 3016 8480 3022 8492
rect 3344 8489 3372 8520
rect 4062 8508 4068 8560
rect 4120 8548 4126 8560
rect 4249 8551 4307 8557
rect 4249 8548 4261 8551
rect 4120 8520 4261 8548
rect 4120 8508 4126 8520
rect 4249 8517 4261 8520
rect 4295 8517 4307 8551
rect 4249 8511 4307 8517
rect 5166 8508 5172 8560
rect 5224 8508 5230 8560
rect 6454 8508 6460 8560
rect 6512 8548 6518 8560
rect 6733 8551 6791 8557
rect 6733 8548 6745 8551
rect 6512 8520 6745 8548
rect 6512 8508 6518 8520
rect 6733 8517 6745 8520
rect 6779 8548 6791 8551
rect 7285 8551 7343 8557
rect 6779 8520 7052 8548
rect 6779 8517 6791 8520
rect 6733 8511 6791 8517
rect 3053 8483 3111 8489
rect 3053 8480 3065 8483
rect 3016 8452 3065 8480
rect 3016 8440 3022 8452
rect 3053 8449 3065 8452
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 3329 8483 3387 8489
rect 3329 8449 3341 8483
rect 3375 8449 3387 8483
rect 3329 8443 3387 8449
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8449 4215 8483
rect 4157 8443 4215 8449
rect 4617 8483 4675 8489
rect 4617 8449 4629 8483
rect 4663 8480 4675 8483
rect 5350 8480 5356 8492
rect 4663 8452 5356 8480
rect 4663 8449 4675 8452
rect 4617 8443 4675 8449
rect 2498 8412 2504 8424
rect 2332 8384 2504 8412
rect 2498 8372 2504 8384
rect 2556 8372 2562 8424
rect 3234 8372 3240 8424
rect 3292 8372 3298 8424
rect 4172 8412 4200 8443
rect 5350 8440 5356 8452
rect 5408 8440 5414 8492
rect 6845 8483 6903 8489
rect 6845 8480 6857 8483
rect 6840 8449 6857 8480
rect 6891 8449 6903 8483
rect 6840 8443 6903 8449
rect 4172 8384 6500 8412
rect 2593 8347 2651 8353
rect 2593 8313 2605 8347
rect 2639 8344 2651 8347
rect 2682 8344 2688 8356
rect 2639 8316 2688 8344
rect 2639 8313 2651 8316
rect 2593 8307 2651 8313
rect 2682 8304 2688 8316
rect 2740 8344 2746 8356
rect 4522 8344 4528 8356
rect 2740 8316 4528 8344
rect 2740 8304 2746 8316
rect 4522 8304 4528 8316
rect 4580 8304 4586 8356
rect 4706 8304 4712 8356
rect 4764 8344 4770 8356
rect 5721 8347 5779 8353
rect 5721 8344 5733 8347
rect 4764 8316 5733 8344
rect 4764 8304 4770 8316
rect 5721 8313 5733 8316
rect 5767 8313 5779 8347
rect 6472 8344 6500 8384
rect 6546 8372 6552 8424
rect 6604 8412 6610 8424
rect 6840 8412 6868 8443
rect 6604 8384 6868 8412
rect 7024 8412 7052 8520
rect 7285 8517 7297 8551
rect 7331 8548 7343 8551
rect 8202 8548 8208 8560
rect 7331 8520 8208 8548
rect 7331 8517 7343 8520
rect 7285 8511 7343 8517
rect 8202 8508 8208 8520
rect 8260 8508 8266 8560
rect 7650 8440 7656 8492
rect 7708 8480 7714 8492
rect 7929 8483 7987 8489
rect 7929 8480 7941 8483
rect 7708 8452 7941 8480
rect 7708 8440 7714 8452
rect 7929 8449 7941 8452
rect 7975 8449 7987 8483
rect 7929 8443 7987 8449
rect 8294 8440 8300 8492
rect 8352 8480 8358 8492
rect 8389 8483 8447 8489
rect 8389 8480 8401 8483
rect 8352 8452 8401 8480
rect 8352 8440 8358 8452
rect 8389 8449 8401 8452
rect 8435 8449 8447 8483
rect 9324 8480 9352 8579
rect 10134 8576 10140 8628
rect 10192 8616 10198 8628
rect 11701 8619 11759 8625
rect 11701 8616 11713 8619
rect 10192 8588 11713 8616
rect 10192 8576 10198 8588
rect 11701 8585 11713 8588
rect 11747 8616 11759 8619
rect 12526 8616 12532 8628
rect 11747 8588 12532 8616
rect 11747 8585 11759 8588
rect 11701 8579 11759 8585
rect 12526 8576 12532 8588
rect 12584 8576 12590 8628
rect 13081 8619 13139 8625
rect 13081 8585 13093 8619
rect 13127 8616 13139 8619
rect 14458 8616 14464 8628
rect 13127 8588 14464 8616
rect 13127 8585 13139 8588
rect 13081 8579 13139 8585
rect 12158 8508 12164 8560
rect 12216 8548 12222 8560
rect 12345 8551 12403 8557
rect 12345 8548 12357 8551
rect 12216 8520 12357 8548
rect 12216 8508 12222 8520
rect 12345 8517 12357 8520
rect 12391 8548 12403 8551
rect 13096 8548 13124 8579
rect 14458 8576 14464 8588
rect 14516 8576 14522 8628
rect 15470 8576 15476 8628
rect 15528 8576 15534 8628
rect 15562 8576 15568 8628
rect 15620 8576 15626 8628
rect 16206 8576 16212 8628
rect 16264 8576 16270 8628
rect 16574 8576 16580 8628
rect 16632 8616 16638 8628
rect 16853 8619 16911 8625
rect 16853 8616 16865 8619
rect 16632 8588 16865 8616
rect 16632 8576 16638 8588
rect 16853 8585 16865 8588
rect 16899 8585 16911 8619
rect 16853 8579 16911 8585
rect 16942 8576 16948 8628
rect 17000 8616 17006 8628
rect 18322 8616 18328 8628
rect 17000 8588 18328 8616
rect 17000 8576 17006 8588
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 18966 8576 18972 8628
rect 19024 8616 19030 8628
rect 19337 8619 19395 8625
rect 19337 8616 19349 8619
rect 19024 8588 19349 8616
rect 19024 8576 19030 8588
rect 19337 8585 19349 8588
rect 19383 8585 19395 8619
rect 19337 8579 19395 8585
rect 19886 8576 19892 8628
rect 19944 8616 19950 8628
rect 20073 8619 20131 8625
rect 20073 8616 20085 8619
rect 19944 8588 20085 8616
rect 19944 8576 19950 8588
rect 20073 8585 20085 8588
rect 20119 8585 20131 8619
rect 20073 8579 20131 8585
rect 12391 8520 13124 8548
rect 12391 8517 12403 8520
rect 12345 8511 12403 8517
rect 14366 8508 14372 8560
rect 14424 8548 14430 8560
rect 15197 8551 15255 8557
rect 15197 8548 15209 8551
rect 14424 8520 15209 8548
rect 14424 8508 14430 8520
rect 15197 8517 15209 8520
rect 15243 8517 15255 8551
rect 15197 8511 15255 8517
rect 15749 8551 15807 8557
rect 15749 8517 15761 8551
rect 15795 8548 15807 8551
rect 16390 8548 16396 8560
rect 15795 8520 16396 8548
rect 15795 8517 15807 8520
rect 15749 8511 15807 8517
rect 16390 8508 16396 8520
rect 16448 8508 16454 8560
rect 19058 8508 19064 8560
rect 19116 8548 19122 8560
rect 19610 8548 19616 8560
rect 19116 8520 19616 8548
rect 19116 8508 19122 8520
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 9324 8452 9873 8480
rect 8389 8443 8447 8449
rect 9861 8449 9873 8452
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8480 10287 8483
rect 10965 8483 11023 8489
rect 10275 8452 10364 8480
rect 10275 8449 10287 8452
rect 10229 8443 10287 8449
rect 8021 8415 8079 8421
rect 8021 8412 8033 8415
rect 7024 8384 8033 8412
rect 6604 8372 6610 8384
rect 8021 8381 8033 8384
rect 8067 8381 8079 8415
rect 8021 8375 8079 8381
rect 6822 8344 6828 8356
rect 6472 8316 6828 8344
rect 5721 8307 5779 8313
rect 6822 8304 6828 8316
rect 6880 8304 6886 8356
rect 9953 8347 10011 8353
rect 9953 8313 9965 8347
rect 9999 8344 10011 8347
rect 10042 8344 10048 8356
rect 9999 8316 10048 8344
rect 9999 8313 10011 8316
rect 9953 8307 10011 8313
rect 10042 8304 10048 8316
rect 10100 8304 10106 8356
rect 10336 8344 10364 8452
rect 10965 8449 10977 8483
rect 11011 8480 11023 8483
rect 11146 8480 11152 8492
rect 11011 8452 11152 8480
rect 11011 8449 11023 8452
rect 10965 8443 11023 8449
rect 11146 8440 11152 8452
rect 11204 8480 11210 8492
rect 11422 8480 11428 8492
rect 11204 8452 11428 8480
rect 11204 8440 11210 8452
rect 11422 8440 11428 8452
rect 11480 8440 11486 8492
rect 11790 8440 11796 8492
rect 11848 8480 11854 8492
rect 12253 8483 12311 8489
rect 12253 8480 12265 8483
rect 11848 8452 12265 8480
rect 11848 8440 11854 8452
rect 12253 8449 12265 8452
rect 12299 8449 12311 8483
rect 12253 8443 12311 8449
rect 12526 8440 12532 8492
rect 12584 8480 12590 8492
rect 13170 8480 13176 8492
rect 12584 8452 13176 8480
rect 12584 8440 12590 8452
rect 13170 8440 13176 8452
rect 13228 8440 13234 8492
rect 13262 8440 13268 8492
rect 13320 8480 13326 8492
rect 13541 8483 13599 8489
rect 13541 8480 13553 8483
rect 13320 8452 13553 8480
rect 13320 8440 13326 8452
rect 13541 8449 13553 8452
rect 13587 8449 13599 8483
rect 13541 8443 13599 8449
rect 13725 8483 13783 8489
rect 13725 8449 13737 8483
rect 13771 8480 13783 8483
rect 13906 8480 13912 8492
rect 13771 8452 13912 8480
rect 13771 8449 13783 8452
rect 13725 8443 13783 8449
rect 10410 8372 10416 8424
rect 10468 8372 10474 8424
rect 10594 8372 10600 8424
rect 10652 8412 10658 8424
rect 11057 8415 11115 8421
rect 11057 8412 11069 8415
rect 10652 8384 11069 8412
rect 10652 8372 10658 8384
rect 11057 8381 11069 8384
rect 11103 8412 11115 8415
rect 13740 8412 13768 8443
rect 13906 8440 13912 8452
rect 13964 8440 13970 8492
rect 13998 8440 14004 8492
rect 14056 8440 14062 8492
rect 14090 8440 14096 8492
rect 14148 8440 14154 8492
rect 14182 8440 14188 8492
rect 14240 8480 14246 8492
rect 15381 8483 15439 8489
rect 15381 8480 15393 8483
rect 14240 8452 15393 8480
rect 14240 8440 14246 8452
rect 15381 8449 15393 8452
rect 15427 8449 15439 8483
rect 15381 8443 15439 8449
rect 11103 8384 12388 8412
rect 11103 8381 11115 8384
rect 11057 8375 11115 8381
rect 11606 8344 11612 8356
rect 10336 8316 11612 8344
rect 11606 8304 11612 8316
rect 11664 8304 11670 8356
rect 12360 8344 12388 8384
rect 12452 8384 13768 8412
rect 14016 8412 14044 8440
rect 14550 8412 14556 8424
rect 14016 8384 14556 8412
rect 12452 8344 12480 8384
rect 14550 8372 14556 8384
rect 14608 8372 14614 8424
rect 14737 8415 14795 8421
rect 14737 8381 14749 8415
rect 14783 8381 14795 8415
rect 15396 8412 15424 8443
rect 15654 8440 15660 8492
rect 15712 8480 15718 8492
rect 17405 8483 17463 8489
rect 17405 8480 17417 8483
rect 15712 8452 17417 8480
rect 15712 8440 15718 8452
rect 17405 8449 17417 8452
rect 17451 8449 17463 8483
rect 17405 8443 17463 8449
rect 16942 8412 16948 8424
rect 15396 8384 16948 8412
rect 14737 8375 14795 8381
rect 12360 8316 12480 8344
rect 12529 8347 12587 8353
rect 12529 8313 12541 8347
rect 12575 8344 12587 8347
rect 13814 8344 13820 8356
rect 12575 8316 13820 8344
rect 12575 8313 12587 8316
rect 12529 8307 12587 8313
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 14752 8344 14780 8375
rect 16942 8372 16948 8384
rect 17000 8372 17006 8424
rect 17420 8412 17448 8443
rect 17494 8440 17500 8492
rect 17552 8480 17558 8492
rect 17589 8483 17647 8489
rect 17589 8480 17601 8483
rect 17552 8452 17601 8480
rect 17552 8440 17558 8452
rect 17589 8449 17601 8452
rect 17635 8449 17647 8483
rect 17589 8443 17647 8449
rect 18138 8440 18144 8492
rect 18196 8440 18202 8492
rect 18325 8483 18383 8489
rect 18325 8449 18337 8483
rect 18371 8480 18383 8483
rect 19150 8480 19156 8492
rect 18371 8452 19156 8480
rect 18371 8449 18383 8452
rect 18325 8443 18383 8449
rect 19150 8440 19156 8452
rect 19208 8440 19214 8492
rect 19260 8489 19288 8520
rect 19610 8508 19616 8520
rect 19668 8508 19674 8560
rect 19245 8483 19303 8489
rect 19245 8449 19257 8483
rect 19291 8449 19303 8483
rect 19245 8443 19303 8449
rect 19426 8440 19432 8492
rect 19484 8440 19490 8492
rect 17770 8412 17776 8424
rect 17420 8384 17776 8412
rect 17770 8372 17776 8384
rect 17828 8372 17834 8424
rect 19886 8412 19892 8424
rect 18524 8384 19892 8412
rect 16758 8344 16764 8356
rect 14752 8316 16764 8344
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 17954 8304 17960 8356
rect 18012 8344 18018 8356
rect 18524 8344 18552 8384
rect 19886 8372 19892 8384
rect 19944 8372 19950 8424
rect 20088 8412 20116 8579
rect 20714 8576 20720 8628
rect 20772 8616 20778 8628
rect 22005 8619 22063 8625
rect 22005 8616 22017 8619
rect 20772 8588 22017 8616
rect 20772 8576 20778 8588
rect 22005 8585 22017 8588
rect 22051 8585 22063 8619
rect 22005 8579 22063 8585
rect 20441 8551 20499 8557
rect 20441 8517 20453 8551
rect 20487 8548 20499 8551
rect 20622 8548 20628 8560
rect 20487 8520 20628 8548
rect 20487 8517 20499 8520
rect 20441 8511 20499 8517
rect 20622 8508 20628 8520
rect 20680 8508 20686 8560
rect 20990 8508 20996 8560
rect 21048 8508 21054 8560
rect 21082 8508 21088 8560
rect 21140 8548 21146 8560
rect 21140 8520 22094 8548
rect 21140 8508 21146 8520
rect 20254 8440 20260 8492
rect 20312 8440 20318 8492
rect 20346 8440 20352 8492
rect 20404 8480 20410 8492
rect 20533 8483 20591 8489
rect 20533 8480 20545 8483
rect 20404 8452 20545 8480
rect 20404 8440 20410 8452
rect 20533 8449 20545 8452
rect 20579 8480 20591 8483
rect 21542 8480 21548 8492
rect 20579 8452 21548 8480
rect 20579 8449 20591 8452
rect 20533 8443 20591 8449
rect 21542 8440 21548 8452
rect 21600 8440 21606 8492
rect 22066 8480 22094 8520
rect 22189 8483 22247 8489
rect 22189 8480 22201 8483
rect 22066 8452 22201 8480
rect 22189 8449 22201 8452
rect 22235 8449 22247 8483
rect 22189 8443 22247 8449
rect 22278 8440 22284 8492
rect 22336 8440 22342 8492
rect 22465 8483 22523 8489
rect 22465 8449 22477 8483
rect 22511 8480 22523 8483
rect 22554 8480 22560 8492
rect 22511 8452 22560 8480
rect 22511 8449 22523 8452
rect 22465 8443 22523 8449
rect 22554 8440 22560 8452
rect 22612 8440 22618 8492
rect 22649 8483 22707 8489
rect 22649 8449 22661 8483
rect 22695 8480 22707 8483
rect 23014 8480 23020 8492
rect 22695 8452 23020 8480
rect 22695 8449 22707 8452
rect 22649 8443 22707 8449
rect 23014 8440 23020 8452
rect 23072 8440 23078 8492
rect 21174 8412 21180 8424
rect 20088 8384 21180 8412
rect 21174 8372 21180 8384
rect 21232 8372 21238 8424
rect 22370 8372 22376 8424
rect 22428 8372 22434 8424
rect 18012 8316 18552 8344
rect 18601 8347 18659 8353
rect 18012 8304 18018 8316
rect 18601 8313 18613 8347
rect 18647 8344 18659 8347
rect 18647 8316 19334 8344
rect 18647 8313 18659 8316
rect 18601 8307 18659 8313
rect 2038 8236 2044 8288
rect 2096 8276 2102 8288
rect 2133 8279 2191 8285
rect 2133 8276 2145 8279
rect 2096 8248 2145 8276
rect 2096 8236 2102 8248
rect 2133 8245 2145 8248
rect 2179 8245 2191 8279
rect 2133 8239 2191 8245
rect 3050 8236 3056 8288
rect 3108 8236 3114 8288
rect 3694 8236 3700 8288
rect 3752 8276 3758 8288
rect 4154 8276 4160 8288
rect 3752 8248 4160 8276
rect 3752 8236 3758 8248
rect 4154 8236 4160 8248
rect 4212 8236 4218 8288
rect 5902 8236 5908 8288
rect 5960 8276 5966 8288
rect 6549 8279 6607 8285
rect 6549 8276 6561 8279
rect 5960 8248 6561 8276
rect 5960 8236 5966 8248
rect 6549 8245 6561 8248
rect 6595 8276 6607 8279
rect 7650 8276 7656 8288
rect 6595 8248 7656 8276
rect 6595 8245 6607 8248
rect 6549 8239 6607 8245
rect 7650 8236 7656 8248
rect 7708 8236 7714 8288
rect 7742 8236 7748 8288
rect 7800 8236 7806 8288
rect 8297 8279 8355 8285
rect 8297 8245 8309 8279
rect 8343 8276 8355 8279
rect 8478 8276 8484 8288
rect 8343 8248 8484 8276
rect 8343 8245 8355 8248
rect 8297 8239 8355 8245
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 8846 8236 8852 8288
rect 8904 8276 8910 8288
rect 9582 8276 9588 8288
rect 8904 8248 9588 8276
rect 8904 8236 8910 8248
rect 9582 8236 9588 8248
rect 9640 8276 9646 8288
rect 10778 8276 10784 8288
rect 9640 8248 10784 8276
rect 9640 8236 9646 8248
rect 10778 8236 10784 8248
rect 10836 8276 10842 8288
rect 11054 8276 11060 8288
rect 10836 8248 11060 8276
rect 10836 8236 10842 8248
rect 11054 8236 11060 8248
rect 11112 8236 11118 8288
rect 19306 8276 19334 8316
rect 19518 8276 19524 8288
rect 19306 8248 19524 8276
rect 19518 8236 19524 8248
rect 19576 8276 19582 8288
rect 20346 8276 20352 8288
rect 19576 8248 20352 8276
rect 19576 8236 19582 8248
rect 20346 8236 20352 8248
rect 20404 8236 20410 8288
rect 1104 8186 23828 8208
rect 1104 8134 3790 8186
rect 3842 8134 3854 8186
rect 3906 8134 3918 8186
rect 3970 8134 3982 8186
rect 4034 8134 4046 8186
rect 4098 8134 9471 8186
rect 9523 8134 9535 8186
rect 9587 8134 9599 8186
rect 9651 8134 9663 8186
rect 9715 8134 9727 8186
rect 9779 8134 15152 8186
rect 15204 8134 15216 8186
rect 15268 8134 15280 8186
rect 15332 8134 15344 8186
rect 15396 8134 15408 8186
rect 15460 8134 20833 8186
rect 20885 8134 20897 8186
rect 20949 8134 20961 8186
rect 21013 8134 21025 8186
rect 21077 8134 21089 8186
rect 21141 8134 23828 8186
rect 1104 8112 23828 8134
rect 2225 8075 2283 8081
rect 2225 8041 2237 8075
rect 2271 8072 2283 8075
rect 2774 8072 2780 8084
rect 2271 8044 2780 8072
rect 2271 8041 2283 8044
rect 2225 8035 2283 8041
rect 2774 8032 2780 8044
rect 2832 8072 2838 8084
rect 3050 8072 3056 8084
rect 2832 8044 3056 8072
rect 2832 8032 2838 8044
rect 3050 8032 3056 8044
rect 3108 8032 3114 8084
rect 4246 8032 4252 8084
rect 4304 8072 4310 8084
rect 4617 8075 4675 8081
rect 4617 8072 4629 8075
rect 4304 8044 4629 8072
rect 4304 8032 4310 8044
rect 4617 8041 4629 8044
rect 4663 8041 4675 8075
rect 4617 8035 4675 8041
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7432 8044 7757 8072
rect 7432 8032 7438 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 7745 8035 7803 8041
rect 8110 8032 8116 8084
rect 8168 8032 8174 8084
rect 9766 8072 9772 8084
rect 9324 8044 9772 8072
rect 4065 8007 4123 8013
rect 4065 7973 4077 8007
rect 4111 8004 4123 8007
rect 4154 8004 4160 8016
rect 4111 7976 4160 8004
rect 4111 7973 4123 7976
rect 4065 7967 4123 7973
rect 4154 7964 4160 7976
rect 4212 8004 4218 8016
rect 5166 8004 5172 8016
rect 4212 7976 5172 8004
rect 4212 7964 4218 7976
rect 5166 7964 5172 7976
rect 5224 7964 5230 8016
rect 6914 7964 6920 8016
rect 6972 8004 6978 8016
rect 9122 8004 9128 8016
rect 6972 7976 9128 8004
rect 6972 7964 6978 7976
rect 9122 7964 9128 7976
rect 9180 7964 9186 8016
rect 4801 7939 4859 7945
rect 4801 7905 4813 7939
rect 4847 7905 4859 7939
rect 4801 7899 4859 7905
rect 7837 7939 7895 7945
rect 7837 7905 7849 7939
rect 7883 7936 7895 7939
rect 8110 7936 8116 7948
rect 7883 7908 8116 7936
rect 7883 7905 7895 7908
rect 7837 7899 7895 7905
rect 2133 7871 2191 7877
rect 2133 7837 2145 7871
rect 2179 7837 2191 7871
rect 2133 7831 2191 7837
rect 2317 7871 2375 7877
rect 2317 7837 2329 7871
rect 2363 7868 2375 7871
rect 2498 7868 2504 7880
rect 2363 7840 2504 7868
rect 2363 7837 2375 7840
rect 2317 7831 2375 7837
rect 2148 7800 2176 7831
rect 2498 7828 2504 7840
rect 2556 7828 2562 7880
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7868 3295 7871
rect 3418 7868 3424 7880
rect 3283 7840 3424 7868
rect 3283 7837 3295 7840
rect 3237 7831 3295 7837
rect 3418 7828 3424 7840
rect 3476 7828 3482 7880
rect 4522 7828 4528 7880
rect 4580 7828 4586 7880
rect 2590 7800 2596 7812
rect 2148 7772 2596 7800
rect 2590 7760 2596 7772
rect 2648 7760 2654 7812
rect 2774 7760 2780 7812
rect 2832 7800 2838 7812
rect 2961 7803 3019 7809
rect 2961 7800 2973 7803
rect 2832 7772 2973 7800
rect 2832 7760 2838 7772
rect 2961 7769 2973 7772
rect 3007 7769 3019 7803
rect 4816 7800 4844 7899
rect 8110 7896 8116 7908
rect 8168 7936 8174 7948
rect 9324 7936 9352 8044
rect 9766 8032 9772 8044
rect 9824 8072 9830 8084
rect 10594 8072 10600 8084
rect 9824 8044 10600 8072
rect 9824 8032 9830 8044
rect 10594 8032 10600 8044
rect 10652 8032 10658 8084
rect 11609 8075 11667 8081
rect 11609 8041 11621 8075
rect 11655 8072 11667 8075
rect 11698 8072 11704 8084
rect 11655 8044 11704 8072
rect 11655 8041 11667 8044
rect 11609 8035 11667 8041
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 12066 8032 12072 8084
rect 12124 8072 12130 8084
rect 12621 8075 12679 8081
rect 12621 8072 12633 8075
rect 12124 8044 12633 8072
rect 12124 8032 12130 8044
rect 12621 8041 12633 8044
rect 12667 8041 12679 8075
rect 12621 8035 12679 8041
rect 12805 8075 12863 8081
rect 12805 8041 12817 8075
rect 12851 8041 12863 8075
rect 12805 8035 12863 8041
rect 10042 7964 10048 8016
rect 10100 8004 10106 8016
rect 11057 8007 11115 8013
rect 10100 7976 11008 8004
rect 10100 7964 10106 7976
rect 10226 7936 10232 7948
rect 8168 7908 9352 7936
rect 9416 7908 10232 7936
rect 8168 7896 8174 7908
rect 5074 7828 5080 7880
rect 5132 7868 5138 7880
rect 5261 7871 5319 7877
rect 5261 7868 5273 7871
rect 5132 7840 5273 7868
rect 5132 7828 5138 7840
rect 5261 7837 5273 7840
rect 5307 7837 5319 7871
rect 5261 7831 5319 7837
rect 5350 7828 5356 7880
rect 5408 7868 5414 7880
rect 6273 7871 6331 7877
rect 6273 7868 6285 7871
rect 5408 7840 6285 7868
rect 5408 7828 5414 7840
rect 6273 7837 6285 7840
rect 6319 7837 6331 7871
rect 6273 7831 6331 7837
rect 6914 7828 6920 7880
rect 6972 7828 6978 7880
rect 7742 7828 7748 7880
rect 7800 7828 7806 7880
rect 9122 7868 9128 7880
rect 7852 7840 9128 7868
rect 5537 7803 5595 7809
rect 5537 7800 5549 7803
rect 4816 7772 5549 7800
rect 2961 7763 3019 7769
rect 5537 7769 5549 7772
rect 5583 7800 5595 7803
rect 5902 7800 5908 7812
rect 5583 7772 5908 7800
rect 5583 7769 5595 7772
rect 5537 7763 5595 7769
rect 5902 7760 5908 7772
rect 5960 7760 5966 7812
rect 6178 7760 6184 7812
rect 6236 7800 6242 7812
rect 6733 7803 6791 7809
rect 6733 7800 6745 7803
rect 6236 7772 6745 7800
rect 6236 7760 6242 7772
rect 6733 7769 6745 7772
rect 6779 7769 6791 7803
rect 6733 7763 6791 7769
rect 4801 7735 4859 7741
rect 4801 7701 4813 7735
rect 4847 7732 4859 7735
rect 5350 7732 5356 7744
rect 4847 7704 5356 7732
rect 4847 7701 4859 7704
rect 4801 7695 4859 7701
rect 5350 7692 5356 7704
rect 5408 7692 5414 7744
rect 6748 7732 6776 7763
rect 7374 7760 7380 7812
rect 7432 7800 7438 7812
rect 7852 7800 7880 7840
rect 9122 7828 9128 7840
rect 9180 7828 9186 7880
rect 9416 7877 9444 7908
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 10980 7936 11008 7976
rect 11057 7973 11069 8007
rect 11103 8004 11115 8007
rect 12820 8004 12848 8035
rect 13722 8032 13728 8084
rect 13780 8032 13786 8084
rect 14553 8075 14611 8081
rect 14553 8041 14565 8075
rect 14599 8072 14611 8075
rect 14734 8072 14740 8084
rect 14599 8044 14740 8072
rect 14599 8041 14611 8044
rect 14553 8035 14611 8041
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 15470 8032 15476 8084
rect 15528 8072 15534 8084
rect 15838 8072 15844 8084
rect 15528 8044 15844 8072
rect 15528 8032 15534 8044
rect 15838 8032 15844 8044
rect 15896 8032 15902 8084
rect 16025 8075 16083 8081
rect 16025 8041 16037 8075
rect 16071 8072 16083 8075
rect 17126 8072 17132 8084
rect 16071 8044 17132 8072
rect 16071 8041 16083 8044
rect 16025 8035 16083 8041
rect 17126 8032 17132 8044
rect 17184 8032 17190 8084
rect 18414 8032 18420 8084
rect 18472 8032 18478 8084
rect 18601 8075 18659 8081
rect 18601 8041 18613 8075
rect 18647 8041 18659 8075
rect 18601 8035 18659 8041
rect 11103 7976 12848 8004
rect 11103 7973 11115 7976
rect 11057 7967 11115 7973
rect 16850 7964 16856 8016
rect 16908 8004 16914 8016
rect 17034 8004 17040 8016
rect 16908 7976 17040 8004
rect 16908 7964 16914 7976
rect 17034 7964 17040 7976
rect 17092 7964 17098 8016
rect 17402 7964 17408 8016
rect 17460 8004 17466 8016
rect 18616 8004 18644 8035
rect 20530 8032 20536 8084
rect 20588 8072 20594 8084
rect 20809 8075 20867 8081
rect 20809 8072 20821 8075
rect 20588 8044 20821 8072
rect 20588 8032 20594 8044
rect 20809 8041 20821 8044
rect 20855 8041 20867 8075
rect 20809 8035 20867 8041
rect 22738 8032 22744 8084
rect 22796 8032 22802 8084
rect 22278 8004 22284 8016
rect 17460 7976 18644 8004
rect 19076 7976 22284 8004
rect 17460 7964 17466 7976
rect 11863 7939 11921 7945
rect 11863 7936 11875 7939
rect 10704 7908 10916 7936
rect 10980 7908 11875 7936
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7837 9551 7871
rect 9493 7831 9551 7837
rect 7432 7772 7880 7800
rect 7432 7760 7438 7772
rect 8386 7760 8392 7812
rect 8444 7800 8450 7812
rect 9309 7803 9367 7809
rect 9309 7800 9321 7803
rect 8444 7772 9321 7800
rect 8444 7760 8450 7772
rect 9309 7769 9321 7772
rect 9355 7769 9367 7803
rect 9508 7800 9536 7831
rect 10318 7828 10324 7880
rect 10376 7828 10382 7880
rect 10704 7877 10732 7908
rect 10413 7871 10471 7877
rect 10413 7837 10425 7871
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7837 10747 7871
rect 10689 7831 10747 7837
rect 10428 7800 10456 7831
rect 10778 7828 10784 7880
rect 10836 7828 10842 7880
rect 10888 7868 10916 7908
rect 11863 7905 11875 7908
rect 11909 7905 11921 7939
rect 11863 7899 11921 7905
rect 12989 7939 13047 7945
rect 12989 7905 13001 7939
rect 13035 7936 13047 7939
rect 15654 7936 15660 7948
rect 13035 7908 15660 7936
rect 13035 7905 13047 7908
rect 12989 7899 13047 7905
rect 15654 7896 15660 7908
rect 15712 7896 15718 7948
rect 16485 7939 16543 7945
rect 16485 7905 16497 7939
rect 16531 7936 16543 7939
rect 16868 7936 16896 7964
rect 16531 7908 16896 7936
rect 16531 7905 16543 7908
rect 16485 7899 16543 7905
rect 17310 7896 17316 7948
rect 17368 7936 17374 7948
rect 17865 7939 17923 7945
rect 17865 7936 17877 7939
rect 17368 7908 17877 7936
rect 17368 7896 17374 7908
rect 17865 7905 17877 7908
rect 17911 7936 17923 7939
rect 19076 7936 19104 7976
rect 22278 7964 22284 7976
rect 22336 7964 22342 8016
rect 17911 7908 19104 7936
rect 17911 7905 17923 7908
rect 17865 7899 17923 7905
rect 20254 7896 20260 7948
rect 20312 7936 20318 7948
rect 20312 7908 22140 7936
rect 20312 7896 20318 7908
rect 11422 7868 11428 7880
rect 10888 7840 11428 7868
rect 11422 7828 11428 7840
rect 11480 7828 11486 7880
rect 11780 7871 11838 7877
rect 11780 7868 11792 7871
rect 11716 7840 11792 7868
rect 9508 7772 10732 7800
rect 9309 7763 9367 7769
rect 8938 7732 8944 7744
rect 6748 7704 8944 7732
rect 8938 7692 8944 7704
rect 8996 7692 9002 7744
rect 9677 7735 9735 7741
rect 9677 7701 9689 7735
rect 9723 7732 9735 7735
rect 10597 7735 10655 7741
rect 10597 7732 10609 7735
rect 9723 7704 10609 7732
rect 9723 7701 9735 7704
rect 9677 7695 9735 7701
rect 10597 7701 10609 7704
rect 10643 7701 10655 7735
rect 10704 7732 10732 7772
rect 11330 7760 11336 7812
rect 11388 7800 11394 7812
rect 11716 7800 11744 7840
rect 11780 7837 11792 7840
rect 11826 7837 11838 7871
rect 11780 7831 11838 7837
rect 11977 7871 12035 7877
rect 11977 7837 11989 7871
rect 12023 7837 12035 7871
rect 11977 7831 12035 7837
rect 12069 7871 12127 7877
rect 12069 7837 12081 7871
rect 12115 7868 12127 7871
rect 12158 7868 12164 7880
rect 12115 7840 12164 7868
rect 12115 7837 12127 7840
rect 12069 7831 12127 7837
rect 11388 7772 11744 7800
rect 11992 7800 12020 7831
rect 12158 7828 12164 7840
rect 12216 7828 12222 7880
rect 12802 7828 12808 7880
rect 12860 7828 12866 7880
rect 14461 7871 14519 7877
rect 14461 7837 14473 7871
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 12710 7800 12716 7812
rect 11992 7772 12716 7800
rect 11388 7760 11394 7772
rect 12710 7760 12716 7772
rect 12768 7760 12774 7812
rect 13078 7760 13084 7812
rect 13136 7760 13142 7812
rect 14476 7800 14504 7831
rect 14642 7828 14648 7880
rect 14700 7828 14706 7880
rect 15194 7828 15200 7880
rect 15252 7868 15258 7880
rect 15562 7868 15568 7880
rect 15252 7840 15568 7868
rect 15252 7828 15258 7840
rect 15562 7828 15568 7840
rect 15620 7868 15626 7880
rect 15930 7868 15936 7880
rect 15620 7840 15936 7868
rect 15620 7828 15626 7840
rect 15672 7809 15700 7840
rect 15930 7828 15936 7840
rect 15988 7828 15994 7880
rect 16850 7828 16856 7880
rect 16908 7828 16914 7880
rect 17037 7871 17095 7877
rect 17037 7837 17049 7871
rect 17083 7837 17095 7871
rect 17037 7831 17095 7837
rect 15657 7803 15715 7809
rect 14476 7772 15056 7800
rect 15028 7744 15056 7772
rect 15657 7769 15669 7803
rect 15703 7769 15715 7803
rect 15657 7763 15715 7769
rect 16482 7760 16488 7812
rect 16540 7800 16546 7812
rect 17052 7800 17080 7831
rect 17218 7828 17224 7880
rect 17276 7828 17282 7880
rect 17402 7828 17408 7880
rect 17460 7828 17466 7880
rect 17770 7828 17776 7880
rect 17828 7868 17834 7880
rect 17828 7840 18628 7868
rect 17828 7828 17834 7840
rect 18555 7837 18628 7840
rect 18138 7800 18144 7812
rect 16540 7772 18144 7800
rect 16540 7760 16546 7772
rect 18138 7760 18144 7772
rect 18196 7760 18202 7812
rect 18555 7803 18567 7837
rect 18601 7806 18628 7837
rect 18690 7828 18696 7880
rect 18748 7868 18754 7880
rect 19429 7871 19487 7877
rect 19429 7868 19441 7871
rect 18748 7840 19441 7868
rect 18748 7828 18754 7840
rect 19429 7837 19441 7840
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 19610 7828 19616 7880
rect 19668 7828 19674 7880
rect 20073 7871 20131 7877
rect 20073 7837 20085 7871
rect 20119 7837 20131 7871
rect 20073 7831 20131 7837
rect 18601 7803 18613 7806
rect 18555 7797 18613 7803
rect 18785 7803 18843 7809
rect 18785 7769 18797 7803
rect 18831 7800 18843 7803
rect 19978 7800 19984 7812
rect 18831 7772 19984 7800
rect 18831 7769 18843 7772
rect 18785 7763 18843 7769
rect 19978 7760 19984 7772
rect 20036 7760 20042 7812
rect 12986 7732 12992 7744
rect 10704 7704 12992 7732
rect 10597 7695 10655 7701
rect 12986 7692 12992 7704
rect 13044 7692 13050 7744
rect 15010 7692 15016 7744
rect 15068 7732 15074 7744
rect 15105 7735 15163 7741
rect 15105 7732 15117 7735
rect 15068 7704 15117 7732
rect 15068 7692 15074 7704
rect 15105 7701 15117 7704
rect 15151 7701 15163 7735
rect 15105 7695 15163 7701
rect 15562 7692 15568 7744
rect 15620 7732 15626 7744
rect 15857 7735 15915 7741
rect 15857 7732 15869 7735
rect 15620 7704 15869 7732
rect 15620 7692 15626 7704
rect 15857 7701 15869 7704
rect 15903 7701 15915 7735
rect 15857 7695 15915 7701
rect 16758 7692 16764 7744
rect 16816 7732 16822 7744
rect 19426 7732 19432 7744
rect 16816 7704 19432 7732
rect 16816 7692 16822 7704
rect 19426 7692 19432 7704
rect 19484 7732 19490 7744
rect 20088 7732 20116 7831
rect 20714 7828 20720 7880
rect 20772 7868 20778 7880
rect 20809 7871 20867 7877
rect 20809 7868 20821 7871
rect 20772 7840 20821 7868
rect 20772 7828 20778 7840
rect 20809 7837 20821 7840
rect 20855 7837 20867 7871
rect 20809 7831 20867 7837
rect 21085 7871 21143 7877
rect 21085 7837 21097 7871
rect 21131 7868 21143 7871
rect 21174 7868 21180 7880
rect 21131 7840 21180 7868
rect 21131 7837 21143 7840
rect 21085 7831 21143 7837
rect 21174 7828 21180 7840
rect 21232 7828 21238 7880
rect 22112 7877 22140 7908
rect 22097 7871 22155 7877
rect 22097 7837 22109 7871
rect 22143 7837 22155 7871
rect 22097 7831 22155 7837
rect 20162 7760 20168 7812
rect 20220 7800 20226 7812
rect 20993 7803 21051 7809
rect 20993 7800 21005 7803
rect 20220 7772 21005 7800
rect 20220 7760 20226 7772
rect 20993 7769 21005 7772
rect 21039 7769 21051 7803
rect 20993 7763 21051 7769
rect 19484 7704 20116 7732
rect 22189 7735 22247 7741
rect 19484 7692 19490 7704
rect 22189 7701 22201 7735
rect 22235 7732 22247 7735
rect 22554 7732 22560 7744
rect 22235 7704 22560 7732
rect 22235 7701 22247 7704
rect 22189 7695 22247 7701
rect 22554 7692 22560 7704
rect 22612 7692 22618 7744
rect 1104 7642 23987 7664
rect 1104 7590 6630 7642
rect 6682 7590 6694 7642
rect 6746 7590 6758 7642
rect 6810 7590 6822 7642
rect 6874 7590 6886 7642
rect 6938 7590 12311 7642
rect 12363 7590 12375 7642
rect 12427 7590 12439 7642
rect 12491 7590 12503 7642
rect 12555 7590 12567 7642
rect 12619 7590 17992 7642
rect 18044 7590 18056 7642
rect 18108 7590 18120 7642
rect 18172 7590 18184 7642
rect 18236 7590 18248 7642
rect 18300 7590 23673 7642
rect 23725 7590 23737 7642
rect 23789 7590 23801 7642
rect 23853 7590 23865 7642
rect 23917 7590 23929 7642
rect 23981 7590 23987 7642
rect 1104 7568 23987 7590
rect 2130 7528 2136 7540
rect 1964 7500 2136 7528
rect 1964 7401 1992 7500
rect 2130 7488 2136 7500
rect 2188 7488 2194 7540
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 4580 7500 4844 7528
rect 4580 7488 4586 7500
rect 2314 7460 2320 7472
rect 2056 7432 2320 7460
rect 2056 7401 2084 7432
rect 2314 7420 2320 7432
rect 2372 7460 2378 7472
rect 2372 7432 4660 7460
rect 2372 7420 2378 7432
rect 1948 7395 2006 7401
rect 1948 7361 1960 7395
rect 1994 7361 2006 7395
rect 1948 7355 2006 7361
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7361 2099 7395
rect 2041 7355 2099 7361
rect 2774 7352 2780 7404
rect 2832 7352 2838 7404
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7392 3019 7395
rect 3881 7395 3939 7401
rect 3881 7392 3893 7395
rect 3007 7364 3893 7392
rect 3007 7361 3019 7364
rect 2961 7355 3019 7361
rect 3881 7361 3893 7364
rect 3927 7392 3939 7395
rect 4154 7392 4160 7404
rect 3927 7364 4160 7392
rect 3927 7361 3939 7364
rect 3881 7355 3939 7361
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 1854 7284 1860 7336
rect 1912 7324 1918 7336
rect 2593 7327 2651 7333
rect 2593 7324 2605 7327
rect 1912 7296 2605 7324
rect 1912 7284 1918 7296
rect 2593 7293 2605 7296
rect 2639 7293 2651 7327
rect 2593 7287 2651 7293
rect 3142 7284 3148 7336
rect 3200 7324 3206 7336
rect 4632 7333 4660 7432
rect 4816 7401 4844 7500
rect 8386 7488 8392 7540
rect 8444 7488 8450 7540
rect 9122 7488 9128 7540
rect 9180 7488 9186 7540
rect 9493 7531 9551 7537
rect 9493 7497 9505 7531
rect 9539 7528 9551 7531
rect 9858 7528 9864 7540
rect 9539 7500 9864 7528
rect 9539 7497 9551 7500
rect 9493 7491 9551 7497
rect 9858 7488 9864 7500
rect 9916 7488 9922 7540
rect 10226 7488 10232 7540
rect 10284 7488 10290 7540
rect 10318 7488 10324 7540
rect 10376 7528 10382 7540
rect 12069 7531 12127 7537
rect 12069 7528 12081 7531
rect 10376 7500 12081 7528
rect 10376 7488 10382 7500
rect 12069 7497 12081 7500
rect 12115 7497 12127 7531
rect 12069 7491 12127 7497
rect 15010 7488 15016 7540
rect 15068 7528 15074 7540
rect 15105 7531 15163 7537
rect 15105 7528 15117 7531
rect 15068 7500 15117 7528
rect 15068 7488 15074 7500
rect 15105 7497 15117 7500
rect 15151 7497 15163 7531
rect 15105 7491 15163 7497
rect 15194 7488 15200 7540
rect 15252 7488 15258 7540
rect 21453 7531 21511 7537
rect 21453 7497 21465 7531
rect 21499 7528 21511 7531
rect 21726 7528 21732 7540
rect 21499 7500 21732 7528
rect 21499 7497 21511 7500
rect 21453 7491 21511 7497
rect 21726 7488 21732 7500
rect 21784 7488 21790 7540
rect 22738 7488 22744 7540
rect 22796 7488 22802 7540
rect 5350 7420 5356 7472
rect 5408 7460 5414 7472
rect 8478 7460 8484 7472
rect 5408 7432 5580 7460
rect 5408 7420 5414 7432
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 4801 7355 4859 7361
rect 4890 7352 4896 7404
rect 4948 7392 4954 7404
rect 5552 7401 5580 7432
rect 7116 7432 8484 7460
rect 5445 7395 5503 7401
rect 5445 7392 5457 7395
rect 4948 7364 5457 7392
rect 4948 7352 4954 7364
rect 5445 7361 5457 7364
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7392 5963 7395
rect 6546 7392 6552 7404
rect 5951 7364 6552 7392
rect 5951 7361 5963 7364
rect 5905 7355 5963 7361
rect 6546 7352 6552 7364
rect 6604 7352 6610 7404
rect 7006 7352 7012 7404
rect 7064 7390 7070 7404
rect 7116 7390 7144 7432
rect 8478 7420 8484 7432
rect 8536 7420 8542 7472
rect 9140 7460 9168 7488
rect 10244 7460 10272 7488
rect 10962 7460 10968 7472
rect 9140 7432 10180 7460
rect 10244 7432 10968 7460
rect 7064 7362 7144 7390
rect 7064 7352 7070 7362
rect 7742 7352 7748 7404
rect 7800 7392 7806 7404
rect 8021 7395 8079 7401
rect 8021 7392 8033 7395
rect 7800 7364 8033 7392
rect 7800 7352 7806 7364
rect 8021 7361 8033 7364
rect 8067 7361 8079 7395
rect 8021 7355 8079 7361
rect 8110 7352 8116 7404
rect 8168 7352 8174 7404
rect 8846 7352 8852 7404
rect 8904 7352 8910 7404
rect 9030 7352 9036 7404
rect 9088 7352 9094 7404
rect 9122 7352 9128 7404
rect 9180 7352 9186 7404
rect 10152 7401 10180 7432
rect 10962 7420 10968 7432
rect 11020 7420 11026 7472
rect 11146 7420 11152 7472
rect 11204 7460 11210 7472
rect 12250 7460 12256 7472
rect 11204 7432 12256 7460
rect 11204 7420 11210 7432
rect 12250 7420 12256 7432
rect 12308 7420 12314 7472
rect 14369 7463 14427 7469
rect 14369 7429 14381 7463
rect 14415 7460 14427 7463
rect 14642 7460 14648 7472
rect 14415 7432 14648 7460
rect 14415 7429 14427 7432
rect 14369 7423 14427 7429
rect 14642 7420 14648 7432
rect 14700 7460 14706 7472
rect 14921 7463 14979 7469
rect 14921 7460 14933 7463
rect 14700 7432 14933 7460
rect 14700 7420 14706 7432
rect 14921 7429 14933 7432
rect 14967 7429 14979 7463
rect 14921 7423 14979 7429
rect 15473 7463 15531 7469
rect 15473 7429 15485 7463
rect 15519 7460 15531 7463
rect 17402 7460 17408 7472
rect 15519 7432 17408 7460
rect 15519 7429 15531 7432
rect 15473 7423 15531 7429
rect 17402 7420 17408 7432
rect 17460 7420 17466 7472
rect 17586 7420 17592 7472
rect 17644 7420 17650 7472
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7361 9275 7395
rect 9217 7355 9275 7361
rect 10137 7395 10195 7401
rect 10137 7361 10149 7395
rect 10183 7361 10195 7395
rect 10137 7355 10195 7361
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7392 10379 7395
rect 10410 7392 10416 7404
rect 10367 7364 10416 7392
rect 10367 7361 10379 7364
rect 10321 7355 10379 7361
rect 3605 7327 3663 7333
rect 3605 7324 3617 7327
rect 3200 7296 3617 7324
rect 3200 7284 3206 7296
rect 3605 7293 3617 7296
rect 3651 7293 3663 7327
rect 3605 7287 3663 7293
rect 4617 7327 4675 7333
rect 4617 7293 4629 7327
rect 4663 7324 4675 7327
rect 6917 7327 6975 7333
rect 6917 7324 6929 7327
rect 4663 7296 6929 7324
rect 4663 7293 4675 7296
rect 4617 7287 4675 7293
rect 6917 7293 6929 7296
rect 6963 7293 6975 7327
rect 6917 7287 6975 7293
rect 7926 7284 7932 7336
rect 7984 7324 7990 7336
rect 8128 7324 8156 7352
rect 7984 7296 8156 7324
rect 7984 7284 7990 7296
rect 8938 7284 8944 7336
rect 8996 7324 9002 7336
rect 9232 7324 9260 7355
rect 10410 7352 10416 7364
rect 10468 7352 10474 7404
rect 11977 7395 12035 7401
rect 11977 7361 11989 7395
rect 12023 7392 12035 7395
rect 12066 7392 12072 7404
rect 12023 7364 12072 7392
rect 12023 7361 12035 7364
rect 11977 7355 12035 7361
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 14090 7352 14096 7404
rect 14148 7392 14154 7404
rect 14274 7392 14280 7404
rect 14148 7364 14280 7392
rect 14148 7352 14154 7364
rect 14274 7352 14280 7364
rect 14332 7352 14338 7404
rect 15289 7395 15347 7401
rect 15289 7361 15301 7395
rect 15335 7392 15347 7395
rect 15838 7392 15844 7404
rect 15335 7364 15844 7392
rect 15335 7361 15347 7364
rect 15289 7355 15347 7361
rect 15838 7352 15844 7364
rect 15896 7352 15902 7404
rect 16758 7352 16764 7404
rect 16816 7392 16822 7404
rect 17034 7401 17040 7404
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 16816 7364 16865 7392
rect 16816 7352 16822 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 17000 7395 17040 7401
rect 17000 7361 17012 7395
rect 17000 7355 17040 7361
rect 17034 7352 17040 7355
rect 17092 7352 17098 7404
rect 18322 7352 18328 7404
rect 18380 7392 18386 7404
rect 18785 7395 18843 7401
rect 18785 7392 18797 7395
rect 18380 7364 18797 7392
rect 18380 7352 18386 7364
rect 18785 7361 18797 7364
rect 18831 7392 18843 7395
rect 18966 7392 18972 7404
rect 18831 7364 18972 7392
rect 18831 7361 18843 7364
rect 18785 7355 18843 7361
rect 18966 7352 18972 7364
rect 19024 7352 19030 7404
rect 19150 7352 19156 7404
rect 19208 7392 19214 7404
rect 19429 7395 19487 7401
rect 19429 7392 19441 7395
rect 19208 7364 19441 7392
rect 19208 7352 19214 7364
rect 19429 7361 19441 7364
rect 19475 7361 19487 7395
rect 21744 7392 21772 7488
rect 22756 7460 22784 7488
rect 22572 7432 22784 7460
rect 22572 7401 22600 7432
rect 22373 7395 22431 7401
rect 22373 7392 22385 7395
rect 21744 7364 22385 7392
rect 19429 7355 19487 7361
rect 22373 7361 22385 7364
rect 22419 7361 22431 7395
rect 22373 7355 22431 7361
rect 22557 7395 22615 7401
rect 22557 7361 22569 7395
rect 22603 7361 22615 7395
rect 22557 7355 22615 7361
rect 22649 7395 22707 7401
rect 22649 7361 22661 7395
rect 22695 7361 22707 7395
rect 22649 7355 22707 7361
rect 22741 7395 22799 7401
rect 22741 7361 22753 7395
rect 22787 7392 22799 7395
rect 22830 7392 22836 7404
rect 22787 7364 22836 7392
rect 22787 7361 22799 7364
rect 22741 7355 22799 7361
rect 11422 7324 11428 7336
rect 8996 7296 11428 7324
rect 8996 7284 9002 7296
rect 11422 7284 11428 7296
rect 11480 7284 11486 7336
rect 16574 7284 16580 7336
rect 16632 7324 16638 7336
rect 17221 7327 17279 7333
rect 17221 7324 17233 7327
rect 16632 7296 17233 7324
rect 16632 7284 16638 7296
rect 17221 7293 17233 7296
rect 17267 7293 17279 7327
rect 17221 7287 17279 7293
rect 19702 7284 19708 7336
rect 19760 7324 19766 7336
rect 20073 7327 20131 7333
rect 20073 7324 20085 7327
rect 19760 7296 20085 7324
rect 19760 7284 19766 7296
rect 20073 7293 20085 7296
rect 20119 7324 20131 7327
rect 20254 7324 20260 7336
rect 20119 7296 20260 7324
rect 20119 7293 20131 7296
rect 20073 7287 20131 7293
rect 20254 7284 20260 7296
rect 20312 7284 20318 7336
rect 20438 7284 20444 7336
rect 20496 7324 20502 7336
rect 22572 7324 22600 7355
rect 20496 7296 22600 7324
rect 20496 7284 20502 7296
rect 8294 7256 8300 7268
rect 7024 7228 8300 7256
rect 1857 7191 1915 7197
rect 1857 7157 1869 7191
rect 1903 7188 1915 7191
rect 2406 7188 2412 7200
rect 1903 7160 2412 7188
rect 1903 7157 1915 7160
rect 1857 7151 1915 7157
rect 2406 7148 2412 7160
rect 2464 7148 2470 7200
rect 5258 7148 5264 7200
rect 5316 7148 5322 7200
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 6270 7188 6276 7200
rect 5868 7160 6276 7188
rect 5868 7148 5874 7160
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 6546 7148 6552 7200
rect 6604 7188 6610 7200
rect 7024 7197 7052 7228
rect 8294 7216 8300 7228
rect 8352 7256 8358 7268
rect 8846 7256 8852 7268
rect 8352 7228 8852 7256
rect 8352 7216 8358 7228
rect 8846 7216 8852 7228
rect 8904 7216 8910 7268
rect 17126 7216 17132 7268
rect 17184 7216 17190 7268
rect 22462 7216 22468 7268
rect 22520 7256 22526 7268
rect 22664 7256 22692 7355
rect 22830 7352 22836 7364
rect 22888 7352 22894 7404
rect 22520 7228 22692 7256
rect 22520 7216 22526 7228
rect 6641 7191 6699 7197
rect 6641 7188 6653 7191
rect 6604 7160 6653 7188
rect 6604 7148 6610 7160
rect 6641 7157 6653 7160
rect 6687 7157 6699 7191
rect 6641 7151 6699 7157
rect 7009 7191 7067 7197
rect 7009 7157 7021 7191
rect 7055 7157 7067 7191
rect 7009 7151 7067 7157
rect 8110 7148 8116 7200
rect 8168 7148 8174 7200
rect 10318 7148 10324 7200
rect 10376 7188 10382 7200
rect 12710 7188 12716 7200
rect 10376 7160 12716 7188
rect 10376 7148 10382 7160
rect 12710 7148 12716 7160
rect 12768 7188 12774 7200
rect 13354 7188 13360 7200
rect 12768 7160 13360 7188
rect 12768 7148 12774 7160
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 15010 7148 15016 7200
rect 15068 7188 15074 7200
rect 15933 7191 15991 7197
rect 15933 7188 15945 7191
rect 15068 7160 15945 7188
rect 15068 7148 15074 7160
rect 15933 7157 15945 7160
rect 15979 7157 15991 7191
rect 15933 7151 15991 7157
rect 22738 7148 22744 7200
rect 22796 7188 22802 7200
rect 23017 7191 23075 7197
rect 23017 7188 23029 7191
rect 22796 7160 23029 7188
rect 22796 7148 22802 7160
rect 23017 7157 23029 7160
rect 23063 7157 23075 7191
rect 23017 7151 23075 7157
rect 1104 7098 23828 7120
rect 1104 7046 3790 7098
rect 3842 7046 3854 7098
rect 3906 7046 3918 7098
rect 3970 7046 3982 7098
rect 4034 7046 4046 7098
rect 4098 7046 9471 7098
rect 9523 7046 9535 7098
rect 9587 7046 9599 7098
rect 9651 7046 9663 7098
rect 9715 7046 9727 7098
rect 9779 7046 15152 7098
rect 15204 7046 15216 7098
rect 15268 7046 15280 7098
rect 15332 7046 15344 7098
rect 15396 7046 15408 7098
rect 15460 7046 20833 7098
rect 20885 7046 20897 7098
rect 20949 7046 20961 7098
rect 21013 7046 21025 7098
rect 21077 7046 21089 7098
rect 21141 7046 23828 7098
rect 1104 7024 23828 7046
rect 2317 6987 2375 6993
rect 2317 6953 2329 6987
rect 2363 6984 2375 6987
rect 2774 6984 2780 6996
rect 2363 6956 2780 6984
rect 2363 6953 2375 6956
rect 2317 6947 2375 6953
rect 2774 6944 2780 6956
rect 2832 6984 2838 6996
rect 8573 6987 8631 6993
rect 2832 6956 3280 6984
rect 2832 6944 2838 6956
rect 3252 6848 3280 6956
rect 8573 6953 8585 6987
rect 8619 6984 8631 6987
rect 9030 6984 9036 6996
rect 8619 6956 9036 6984
rect 8619 6953 8631 6956
rect 8573 6947 8631 6953
rect 9030 6944 9036 6956
rect 9088 6944 9094 6996
rect 10410 6944 10416 6996
rect 10468 6944 10474 6996
rect 13078 6944 13084 6996
rect 13136 6984 13142 6996
rect 13265 6987 13323 6993
rect 13265 6984 13277 6987
rect 13136 6956 13277 6984
rect 13136 6944 13142 6956
rect 13265 6953 13277 6956
rect 13311 6953 13323 6987
rect 13265 6947 13323 6953
rect 16574 6944 16580 6996
rect 16632 6984 16638 6996
rect 16669 6987 16727 6993
rect 16669 6984 16681 6987
rect 16632 6956 16681 6984
rect 16632 6944 16638 6956
rect 16669 6953 16681 6956
rect 16715 6953 16727 6987
rect 16669 6947 16727 6953
rect 8386 6916 8392 6928
rect 5184 6888 6224 6916
rect 4522 6848 4528 6860
rect 3252 6820 4528 6848
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6780 2007 6783
rect 2130 6780 2136 6792
rect 1995 6752 2136 6780
rect 1995 6749 2007 6752
rect 1949 6743 2007 6749
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 3252 6789 3280 6820
rect 4522 6808 4528 6820
rect 4580 6808 4586 6860
rect 4614 6808 4620 6860
rect 4672 6848 4678 6860
rect 4709 6851 4767 6857
rect 4709 6848 4721 6851
rect 4672 6820 4721 6848
rect 4672 6808 4678 6820
rect 4709 6817 4721 6820
rect 4755 6817 4767 6851
rect 4709 6811 4767 6817
rect 2317 6783 2375 6789
rect 2317 6749 2329 6783
rect 2363 6780 2375 6783
rect 3053 6783 3111 6789
rect 3053 6780 3065 6783
rect 2363 6752 3065 6780
rect 2363 6749 2375 6752
rect 2317 6743 2375 6749
rect 3053 6749 3065 6752
rect 3099 6749 3111 6783
rect 3053 6743 3111 6749
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6749 3295 6783
rect 3237 6743 3295 6749
rect 3329 6783 3387 6789
rect 3329 6749 3341 6783
rect 3375 6780 3387 6783
rect 4249 6783 4307 6789
rect 4249 6780 4261 6783
rect 3375 6752 4261 6780
rect 3375 6749 3387 6752
rect 3329 6743 3387 6749
rect 4249 6749 4261 6752
rect 4295 6780 4307 6783
rect 4295 6752 4568 6780
rect 4295 6749 4307 6752
rect 4249 6743 4307 6749
rect 3068 6712 3096 6743
rect 4157 6715 4215 6721
rect 3068 6684 3188 6712
rect 3160 6656 3188 6684
rect 4157 6681 4169 6715
rect 4203 6681 4215 6715
rect 4157 6675 4215 6681
rect 2501 6647 2559 6653
rect 2501 6613 2513 6647
rect 2547 6644 2559 6647
rect 2682 6644 2688 6656
rect 2547 6616 2688 6644
rect 2547 6613 2559 6616
rect 2501 6607 2559 6613
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 3142 6604 3148 6656
rect 3200 6604 3206 6656
rect 4172 6644 4200 6675
rect 4246 6644 4252 6656
rect 4172 6616 4252 6644
rect 4246 6604 4252 6616
rect 4304 6604 4310 6656
rect 4540 6644 4568 6752
rect 4617 6715 4675 6721
rect 4617 6681 4629 6715
rect 4663 6712 4675 6715
rect 5184 6712 5212 6888
rect 5258 6808 5264 6860
rect 5316 6848 5322 6860
rect 6089 6851 6147 6857
rect 6089 6848 6101 6851
rect 5316 6820 6101 6848
rect 5316 6808 5322 6820
rect 6089 6817 6101 6820
rect 6135 6817 6147 6851
rect 6196 6848 6224 6888
rect 8128 6888 8392 6916
rect 7469 6851 7527 6857
rect 6196 6820 7420 6848
rect 6089 6811 6147 6817
rect 5629 6783 5687 6789
rect 5629 6749 5641 6783
rect 5675 6780 5687 6783
rect 5718 6780 5724 6792
rect 5675 6752 5724 6780
rect 5675 6749 5687 6752
rect 5629 6743 5687 6749
rect 5718 6740 5724 6752
rect 5776 6740 5782 6792
rect 5810 6740 5816 6792
rect 5868 6740 5874 6792
rect 6181 6783 6239 6789
rect 6181 6749 6193 6783
rect 6227 6749 6239 6783
rect 7392 6780 7420 6820
rect 7469 6817 7481 6851
rect 7515 6848 7527 6851
rect 8128 6848 8156 6888
rect 8386 6876 8392 6888
rect 8444 6876 8450 6928
rect 10428 6916 10456 6944
rect 9232 6888 10456 6916
rect 7515 6820 8156 6848
rect 7515 6817 7527 6820
rect 7469 6811 7527 6817
rect 7834 6780 7840 6792
rect 7392 6752 7840 6780
rect 6181 6743 6239 6749
rect 4663 6684 5212 6712
rect 4663 6681 4675 6684
rect 4617 6675 4675 6681
rect 5442 6672 5448 6724
rect 5500 6712 5506 6724
rect 6196 6712 6224 6743
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 7944 6789 7972 6820
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 9232 6848 9260 6888
rect 11698 6876 11704 6928
rect 11756 6916 11762 6928
rect 11756 6888 12296 6916
rect 11756 6876 11762 6888
rect 8260 6820 9260 6848
rect 8260 6808 8266 6820
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 8022 6783 8080 6789
rect 8022 6749 8034 6783
rect 8068 6780 8080 6783
rect 8110 6780 8116 6792
rect 8068 6752 8116 6780
rect 8068 6749 8080 6752
rect 8022 6743 8080 6749
rect 5500 6684 6224 6712
rect 5500 6672 5506 6684
rect 6822 6672 6828 6724
rect 6880 6672 6886 6724
rect 5534 6644 5540 6656
rect 4540 6616 5540 6644
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 5718 6604 5724 6656
rect 5776 6644 5782 6656
rect 8036 6644 8064 6743
rect 8110 6740 8116 6752
rect 8168 6740 8174 6792
rect 8294 6740 8300 6792
rect 8352 6740 8358 6792
rect 8404 6789 8432 6820
rect 9950 6808 9956 6860
rect 10008 6808 10014 6860
rect 10042 6808 10048 6860
rect 10100 6848 10106 6860
rect 10229 6851 10287 6857
rect 10229 6848 10241 6851
rect 10100 6820 10241 6848
rect 10100 6808 10106 6820
rect 10229 6817 10241 6820
rect 10275 6817 10287 6851
rect 10229 6811 10287 6817
rect 10318 6808 10324 6860
rect 10376 6808 10382 6860
rect 10413 6851 10471 6857
rect 10413 6817 10425 6851
rect 10459 6848 10471 6851
rect 12158 6848 12164 6860
rect 10459 6820 12164 6848
rect 10459 6817 10471 6820
rect 10413 6811 10471 6817
rect 12158 6808 12164 6820
rect 12216 6808 12222 6860
rect 12268 6848 12296 6888
rect 12986 6876 12992 6928
rect 13044 6916 13050 6928
rect 13633 6919 13691 6925
rect 13633 6916 13645 6919
rect 13044 6888 13645 6916
rect 13044 6876 13050 6888
rect 13633 6885 13645 6888
rect 13679 6916 13691 6919
rect 13722 6916 13728 6928
rect 13679 6888 13728 6916
rect 13679 6885 13691 6888
rect 13633 6879 13691 6885
rect 13722 6876 13728 6888
rect 13780 6876 13786 6928
rect 12268 6820 13768 6848
rect 8394 6783 8452 6789
rect 8394 6749 8406 6783
rect 8440 6749 8452 6783
rect 10134 6780 10140 6792
rect 8394 6743 8452 6749
rect 9324 6752 10140 6780
rect 8205 6715 8263 6721
rect 8205 6681 8217 6715
rect 8251 6712 8263 6715
rect 9324 6712 9352 6752
rect 10134 6740 10140 6752
rect 10192 6780 10198 6792
rect 10870 6780 10876 6792
rect 10192 6752 10876 6780
rect 10192 6740 10198 6752
rect 10870 6740 10876 6752
rect 10928 6740 10934 6792
rect 10962 6740 10968 6792
rect 11020 6780 11026 6792
rect 11609 6783 11667 6789
rect 11609 6780 11621 6783
rect 11020 6752 11621 6780
rect 11020 6740 11026 6752
rect 11609 6749 11621 6752
rect 11655 6749 11667 6783
rect 11609 6743 11667 6749
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6780 11943 6783
rect 12066 6780 12072 6792
rect 11931 6752 12072 6780
rect 11931 6749 11943 6752
rect 11885 6743 11943 6749
rect 11900 6712 11928 6743
rect 12066 6740 12072 6752
rect 12124 6740 12130 6792
rect 13446 6740 13452 6792
rect 13504 6740 13510 6792
rect 13740 6789 13768 6820
rect 13906 6808 13912 6860
rect 13964 6848 13970 6860
rect 13964 6820 15332 6848
rect 13964 6808 13970 6820
rect 13725 6783 13783 6789
rect 13725 6749 13737 6783
rect 13771 6780 13783 6783
rect 14090 6780 14096 6792
rect 13771 6752 14096 6780
rect 13771 6749 13783 6752
rect 13725 6743 13783 6749
rect 14090 6740 14096 6752
rect 14148 6740 14154 6792
rect 14274 6740 14280 6792
rect 14332 6780 14338 6792
rect 15304 6789 15332 6820
rect 17034 6808 17040 6860
rect 17092 6848 17098 6860
rect 17313 6851 17371 6857
rect 17313 6848 17325 6851
rect 17092 6820 17325 6848
rect 17092 6808 17098 6820
rect 17313 6817 17325 6820
rect 17359 6817 17371 6851
rect 17313 6811 17371 6817
rect 17773 6851 17831 6857
rect 17773 6817 17785 6851
rect 17819 6848 17831 6851
rect 18322 6848 18328 6860
rect 17819 6820 18328 6848
rect 17819 6817 17831 6820
rect 17773 6811 17831 6817
rect 18322 6808 18328 6820
rect 18380 6808 18386 6860
rect 18966 6808 18972 6860
rect 19024 6848 19030 6860
rect 19889 6851 19947 6857
rect 19889 6848 19901 6851
rect 19024 6820 19901 6848
rect 19024 6808 19030 6820
rect 19889 6817 19901 6820
rect 19935 6817 19947 6851
rect 19889 6811 19947 6817
rect 21729 6851 21787 6857
rect 21729 6817 21741 6851
rect 21775 6848 21787 6851
rect 21775 6820 22094 6848
rect 21775 6817 21787 6820
rect 21729 6811 21787 6817
rect 15105 6783 15163 6789
rect 15105 6780 15117 6783
rect 14332 6752 15117 6780
rect 14332 6740 14338 6752
rect 15105 6749 15117 6752
rect 15151 6749 15163 6783
rect 15105 6743 15163 6749
rect 15289 6783 15347 6789
rect 15289 6749 15301 6783
rect 15335 6780 15347 6783
rect 16114 6780 16120 6792
rect 15335 6752 16120 6780
rect 15335 6749 15347 6752
rect 15289 6743 15347 6749
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 17497 6783 17555 6789
rect 17497 6749 17509 6783
rect 17543 6780 17555 6783
rect 18877 6783 18935 6789
rect 18877 6780 18889 6783
rect 17543 6752 18889 6780
rect 17543 6749 17555 6752
rect 17497 6743 17555 6749
rect 18877 6749 18889 6752
rect 18923 6780 18935 6783
rect 19058 6780 19064 6792
rect 18923 6752 19064 6780
rect 18923 6749 18935 6752
rect 18877 6743 18935 6749
rect 19058 6740 19064 6752
rect 19116 6740 19122 6792
rect 19334 6780 19340 6792
rect 19168 6752 19340 6780
rect 8251 6684 9352 6712
rect 9416 6684 11928 6712
rect 18325 6715 18383 6721
rect 8251 6681 8263 6684
rect 8205 6675 8263 6681
rect 9416 6644 9444 6684
rect 18325 6681 18337 6715
rect 18371 6712 18383 6715
rect 19168 6712 19196 6752
rect 19334 6740 19340 6752
rect 19392 6740 19398 6792
rect 19426 6740 19432 6792
rect 19484 6740 19490 6792
rect 19610 6740 19616 6792
rect 19668 6740 19674 6792
rect 19981 6783 20039 6789
rect 19981 6749 19993 6783
rect 20027 6749 20039 6783
rect 19981 6743 20039 6749
rect 18371 6684 19196 6712
rect 18371 6681 18383 6684
rect 18325 6675 18383 6681
rect 19242 6672 19248 6724
rect 19300 6712 19306 6724
rect 19996 6712 20024 6743
rect 20622 6740 20628 6792
rect 20680 6780 20686 6792
rect 21085 6783 21143 6789
rect 21085 6780 21097 6783
rect 20680 6752 21097 6780
rect 20680 6740 20686 6752
rect 21085 6749 21097 6752
rect 21131 6749 21143 6783
rect 21085 6743 21143 6749
rect 21266 6740 21272 6792
rect 21324 6740 21330 6792
rect 21361 6783 21419 6789
rect 21361 6749 21373 6783
rect 21407 6749 21419 6783
rect 21361 6743 21419 6749
rect 21453 6783 21511 6789
rect 21453 6749 21465 6783
rect 21499 6780 21511 6783
rect 21542 6780 21548 6792
rect 21499 6752 21548 6780
rect 21499 6749 21511 6752
rect 21453 6743 21511 6749
rect 19300 6684 20024 6712
rect 19300 6672 19306 6684
rect 5776 6616 9444 6644
rect 9493 6647 9551 6653
rect 5776 6604 5782 6616
rect 9493 6613 9505 6647
rect 9539 6644 9551 6647
rect 9674 6644 9680 6656
rect 9539 6616 9680 6644
rect 9539 6613 9551 6616
rect 9493 6607 9551 6613
rect 9674 6604 9680 6616
rect 9732 6644 9738 6656
rect 10318 6644 10324 6656
rect 9732 6616 10324 6644
rect 9732 6604 9738 6616
rect 10318 6604 10324 6616
rect 10376 6604 10382 6656
rect 10594 6604 10600 6656
rect 10652 6644 10658 6656
rect 11425 6647 11483 6653
rect 11425 6644 11437 6647
rect 10652 6616 11437 6644
rect 10652 6604 10658 6616
rect 11425 6613 11437 6616
rect 11471 6613 11483 6647
rect 11425 6607 11483 6613
rect 11606 6604 11612 6656
rect 11664 6644 11670 6656
rect 11793 6647 11851 6653
rect 11793 6644 11805 6647
rect 11664 6616 11805 6644
rect 11664 6604 11670 6616
rect 11793 6613 11805 6616
rect 11839 6613 11851 6647
rect 11793 6607 11851 6613
rect 12250 6604 12256 6656
rect 12308 6644 12314 6656
rect 13170 6644 13176 6656
rect 12308 6616 13176 6644
rect 12308 6604 12314 6616
rect 13170 6604 13176 6616
rect 13228 6604 13234 6656
rect 15197 6647 15255 6653
rect 15197 6613 15209 6647
rect 15243 6644 15255 6647
rect 15562 6644 15568 6656
rect 15243 6616 15568 6644
rect 15243 6613 15255 6616
rect 15197 6607 15255 6613
rect 15562 6604 15568 6616
rect 15620 6604 15626 6656
rect 18874 6604 18880 6656
rect 18932 6644 18938 6656
rect 20349 6647 20407 6653
rect 20349 6644 20361 6647
rect 18932 6616 20361 6644
rect 18932 6604 18938 6616
rect 20349 6613 20361 6616
rect 20395 6613 20407 6647
rect 20349 6607 20407 6613
rect 20530 6604 20536 6656
rect 20588 6644 20594 6656
rect 21376 6644 21404 6743
rect 21542 6740 21548 6752
rect 21600 6740 21606 6792
rect 22066 6780 22094 6820
rect 22186 6808 22192 6860
rect 22244 6808 22250 6860
rect 22646 6808 22652 6860
rect 22704 6808 22710 6860
rect 22373 6783 22431 6789
rect 22373 6780 22385 6783
rect 22066 6752 22385 6780
rect 22373 6749 22385 6752
rect 22419 6749 22431 6783
rect 22373 6743 22431 6749
rect 22465 6783 22523 6789
rect 22465 6749 22477 6783
rect 22511 6749 22523 6783
rect 22465 6743 22523 6749
rect 21634 6672 21640 6724
rect 21692 6712 21698 6724
rect 22480 6712 22508 6743
rect 22738 6740 22744 6792
rect 22796 6740 22802 6792
rect 21692 6684 22508 6712
rect 21692 6672 21698 6684
rect 22094 6644 22100 6656
rect 20588 6616 22100 6644
rect 20588 6604 20594 6616
rect 22094 6604 22100 6616
rect 22152 6604 22158 6656
rect 1104 6554 23987 6576
rect 1104 6502 6630 6554
rect 6682 6502 6694 6554
rect 6746 6502 6758 6554
rect 6810 6502 6822 6554
rect 6874 6502 6886 6554
rect 6938 6502 12311 6554
rect 12363 6502 12375 6554
rect 12427 6502 12439 6554
rect 12491 6502 12503 6554
rect 12555 6502 12567 6554
rect 12619 6502 17992 6554
rect 18044 6502 18056 6554
rect 18108 6502 18120 6554
rect 18172 6502 18184 6554
rect 18236 6502 18248 6554
rect 18300 6502 23673 6554
rect 23725 6502 23737 6554
rect 23789 6502 23801 6554
rect 23853 6502 23865 6554
rect 23917 6502 23929 6554
rect 23981 6502 23987 6554
rect 1104 6480 23987 6502
rect 3421 6443 3479 6449
rect 3421 6409 3433 6443
rect 3467 6440 3479 6443
rect 9674 6440 9680 6452
rect 3467 6412 9680 6440
rect 3467 6409 3479 6412
rect 3421 6403 3479 6409
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 10042 6400 10048 6452
rect 10100 6440 10106 6452
rect 10100 6412 12664 6440
rect 10100 6400 10106 6412
rect 4338 6332 4344 6384
rect 4396 6372 4402 6384
rect 4396 6344 8340 6372
rect 4396 6332 4402 6344
rect 2222 6264 2228 6316
rect 2280 6264 2286 6316
rect 2406 6264 2412 6316
rect 2464 6264 2470 6316
rect 2682 6264 2688 6316
rect 2740 6264 2746 6316
rect 2958 6264 2964 6316
rect 3016 6264 3022 6316
rect 3050 6264 3056 6316
rect 3108 6264 3114 6316
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6304 4215 6307
rect 4430 6304 4436 6316
rect 4203 6276 4436 6304
rect 4203 6273 4215 6276
rect 4157 6267 4215 6273
rect 4430 6264 4436 6276
rect 4488 6264 4494 6316
rect 4614 6264 4620 6316
rect 4672 6264 4678 6316
rect 4893 6307 4951 6313
rect 4893 6304 4905 6307
rect 4724 6276 4905 6304
rect 4724 6236 4752 6276
rect 4893 6273 4905 6276
rect 4939 6273 4951 6307
rect 4893 6267 4951 6273
rect 5353 6307 5411 6313
rect 5353 6273 5365 6307
rect 5399 6304 5411 6307
rect 5442 6304 5448 6316
rect 5399 6276 5448 6304
rect 5399 6273 5411 6276
rect 5353 6267 5411 6273
rect 5442 6264 5448 6276
rect 5500 6264 5506 6316
rect 5902 6264 5908 6316
rect 5960 6304 5966 6316
rect 6549 6307 6607 6313
rect 6549 6304 6561 6307
rect 5960 6276 6561 6304
rect 5960 6264 5966 6276
rect 6549 6273 6561 6276
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6638 6264 6644 6316
rect 6696 6304 6702 6316
rect 6733 6307 6791 6313
rect 6733 6304 6745 6307
rect 6696 6276 6745 6304
rect 6696 6264 6702 6276
rect 6733 6273 6745 6276
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 7374 6264 7380 6316
rect 7432 6264 7438 6316
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6304 7987 6307
rect 8202 6304 8208 6316
rect 7975 6276 8208 6304
rect 7975 6273 7987 6276
rect 7929 6267 7987 6273
rect 8202 6264 8208 6276
rect 8260 6264 8266 6316
rect 8312 6313 8340 6344
rect 12066 6332 12072 6384
rect 12124 6372 12130 6384
rect 12253 6375 12311 6381
rect 12253 6372 12265 6375
rect 12124 6344 12265 6372
rect 12124 6332 12130 6344
rect 12253 6341 12265 6344
rect 12299 6341 12311 6375
rect 12463 6375 12521 6381
rect 12463 6372 12475 6375
rect 12253 6335 12311 6341
rect 12452 6341 12475 6372
rect 12509 6341 12521 6375
rect 12452 6335 12521 6341
rect 8297 6307 8355 6313
rect 8297 6273 8309 6307
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6273 8447 6307
rect 8389 6267 8447 6273
rect 7392 6236 7420 6264
rect 2746 6208 4752 6236
rect 4908 6208 7420 6236
rect 2130 6128 2136 6180
rect 2188 6168 2194 6180
rect 2746 6168 2774 6208
rect 4908 6180 4936 6208
rect 7742 6196 7748 6248
rect 7800 6236 7806 6248
rect 8404 6236 8432 6267
rect 8938 6264 8944 6316
rect 8996 6264 9002 6316
rect 12161 6307 12219 6313
rect 12161 6304 12173 6307
rect 9140 6276 12173 6304
rect 9140 6245 9168 6276
rect 12161 6273 12173 6276
rect 12207 6273 12219 6307
rect 12161 6267 12219 6273
rect 12345 6307 12403 6313
rect 12345 6273 12357 6307
rect 12391 6273 12403 6307
rect 12345 6267 12403 6273
rect 7800 6208 8432 6236
rect 9125 6239 9183 6245
rect 7800 6196 7806 6208
rect 9125 6205 9137 6239
rect 9171 6205 9183 6239
rect 9125 6199 9183 6205
rect 11054 6196 11060 6248
rect 11112 6236 11118 6248
rect 12250 6236 12256 6248
rect 11112 6208 12256 6236
rect 11112 6196 11118 6208
rect 12250 6196 12256 6208
rect 12308 6236 12314 6248
rect 12360 6236 12388 6267
rect 12308 6208 12388 6236
rect 12452 6236 12480 6335
rect 12636 6313 12664 6412
rect 18322 6400 18328 6452
rect 18380 6440 18386 6452
rect 18782 6440 18788 6452
rect 18380 6412 18788 6440
rect 18380 6400 18386 6412
rect 18782 6400 18788 6412
rect 18840 6440 18846 6452
rect 18969 6443 19027 6449
rect 18969 6440 18981 6443
rect 18840 6412 18981 6440
rect 18840 6400 18846 6412
rect 18969 6409 18981 6412
rect 19015 6409 19027 6443
rect 18969 6403 19027 6409
rect 21453 6443 21511 6449
rect 21453 6409 21465 6443
rect 21499 6440 21511 6443
rect 22370 6440 22376 6452
rect 21499 6412 22376 6440
rect 21499 6409 21511 6412
rect 21453 6403 21511 6409
rect 22370 6400 22376 6412
rect 22428 6400 22434 6452
rect 23014 6400 23020 6452
rect 23072 6400 23078 6452
rect 13170 6332 13176 6384
rect 13228 6372 13234 6384
rect 16482 6372 16488 6384
rect 13228 6344 14780 6372
rect 13228 6332 13234 6344
rect 12621 6307 12679 6313
rect 12621 6273 12633 6307
rect 12667 6273 12679 6307
rect 12621 6267 12679 6273
rect 13446 6264 13452 6316
rect 13504 6304 13510 6316
rect 13817 6307 13875 6313
rect 13817 6304 13829 6307
rect 13504 6276 13829 6304
rect 13504 6264 13510 6276
rect 13817 6273 13829 6276
rect 13863 6273 13875 6307
rect 13817 6267 13875 6273
rect 13464 6236 13492 6264
rect 12452 6208 13492 6236
rect 12308 6196 12314 6208
rect 2188 6140 2774 6168
rect 2188 6128 2194 6140
rect 3050 6128 3056 6180
rect 3108 6168 3114 6180
rect 4154 6168 4160 6180
rect 3108 6140 4160 6168
rect 3108 6128 3114 6140
rect 4154 6128 4160 6140
rect 4212 6128 4218 6180
rect 4709 6171 4767 6177
rect 4709 6137 4721 6171
rect 4755 6168 4767 6171
rect 4890 6168 4896 6180
rect 4755 6140 4896 6168
rect 4755 6137 4767 6140
rect 4709 6131 4767 6137
rect 4890 6128 4896 6140
rect 4948 6128 4954 6180
rect 4982 6128 4988 6180
rect 5040 6168 5046 6180
rect 11977 6171 12035 6177
rect 11977 6168 11989 6171
rect 5040 6140 11989 6168
rect 5040 6128 5046 6140
rect 11977 6137 11989 6140
rect 12023 6137 12035 6171
rect 13832 6168 13860 6267
rect 14752 6248 14780 6344
rect 15488 6344 16488 6372
rect 15488 6313 15516 6344
rect 16482 6332 16488 6344
rect 16540 6332 16546 6384
rect 18049 6375 18107 6381
rect 18049 6341 18061 6375
rect 18095 6372 18107 6375
rect 19610 6372 19616 6384
rect 18095 6344 19616 6372
rect 18095 6341 18107 6344
rect 18049 6335 18107 6341
rect 19610 6332 19616 6344
rect 19668 6372 19674 6384
rect 19668 6344 19748 6372
rect 19668 6332 19674 6344
rect 15473 6307 15531 6313
rect 15473 6273 15485 6307
rect 15519 6273 15531 6307
rect 15473 6267 15531 6273
rect 15562 6264 15568 6316
rect 15620 6304 15626 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 15620 6276 16865 6304
rect 15620 6264 15626 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 17037 6307 17095 6313
rect 17037 6273 17049 6307
rect 17083 6304 17095 6307
rect 17126 6304 17132 6316
rect 17083 6276 17132 6304
rect 17083 6273 17095 6276
rect 17037 6267 17095 6273
rect 17126 6264 17132 6276
rect 17184 6264 17190 6316
rect 17402 6264 17408 6316
rect 17460 6264 17466 6316
rect 18509 6307 18567 6313
rect 18509 6273 18521 6307
rect 18555 6273 18567 6307
rect 18509 6267 18567 6273
rect 14090 6196 14096 6248
rect 14148 6236 14154 6248
rect 14550 6236 14556 6248
rect 14148 6208 14556 6236
rect 14148 6196 14154 6208
rect 14550 6196 14556 6208
rect 14608 6196 14614 6248
rect 14734 6196 14740 6248
rect 14792 6236 14798 6248
rect 15010 6236 15016 6248
rect 14792 6208 15016 6236
rect 14792 6196 14798 6208
rect 15010 6196 15016 6208
rect 15068 6236 15074 6248
rect 15381 6239 15439 6245
rect 15381 6236 15393 6239
rect 15068 6208 15393 6236
rect 15068 6196 15074 6208
rect 15381 6205 15393 6208
rect 15427 6236 15439 6239
rect 15427 6208 15700 6236
rect 15427 6205 15439 6208
rect 15381 6199 15439 6205
rect 15562 6168 15568 6180
rect 13832 6140 15568 6168
rect 11977 6131 12035 6137
rect 15562 6128 15568 6140
rect 15620 6128 15626 6180
rect 4065 6103 4123 6109
rect 4065 6069 4077 6103
rect 4111 6100 4123 6103
rect 4246 6100 4252 6112
rect 4111 6072 4252 6100
rect 4111 6069 4123 6072
rect 4065 6063 4123 6069
rect 4246 6060 4252 6072
rect 4304 6060 4310 6112
rect 4430 6060 4436 6112
rect 4488 6100 4494 6112
rect 5810 6100 5816 6112
rect 4488 6072 5816 6100
rect 4488 6060 4494 6072
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 5997 6103 6055 6109
rect 5997 6069 6009 6103
rect 6043 6100 6055 6103
rect 6362 6100 6368 6112
rect 6043 6072 6368 6100
rect 6043 6069 6055 6072
rect 5997 6063 6055 6069
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 6549 6103 6607 6109
rect 6549 6069 6561 6103
rect 6595 6100 6607 6103
rect 9306 6100 9312 6112
rect 6595 6072 9312 6100
rect 6595 6069 6607 6072
rect 6549 6063 6607 6069
rect 9306 6060 9312 6072
rect 9364 6060 9370 6112
rect 9398 6060 9404 6112
rect 9456 6100 9462 6112
rect 13538 6100 13544 6112
rect 9456 6072 13544 6100
rect 9456 6060 9462 6072
rect 13538 6060 13544 6072
rect 13596 6060 13602 6112
rect 13630 6060 13636 6112
rect 13688 6060 13694 6112
rect 13998 6060 14004 6112
rect 14056 6060 14062 6112
rect 15197 6103 15255 6109
rect 15197 6069 15209 6103
rect 15243 6100 15255 6103
rect 15470 6100 15476 6112
rect 15243 6072 15476 6100
rect 15243 6069 15255 6072
rect 15197 6063 15255 6069
rect 15470 6060 15476 6072
rect 15528 6060 15534 6112
rect 15672 6100 15700 6208
rect 15746 6196 15752 6248
rect 15804 6196 15810 6248
rect 15841 6239 15899 6245
rect 15841 6205 15853 6239
rect 15887 6236 15899 6239
rect 16758 6236 16764 6248
rect 15887 6208 16764 6236
rect 15887 6205 15899 6208
rect 15841 6199 15899 6205
rect 16758 6196 16764 6208
rect 16816 6196 16822 6248
rect 17313 6239 17371 6245
rect 17313 6205 17325 6239
rect 17359 6205 17371 6239
rect 17313 6199 17371 6205
rect 15930 6128 15936 6180
rect 15988 6168 15994 6180
rect 17328 6168 17356 6199
rect 18230 6196 18236 6248
rect 18288 6236 18294 6248
rect 18524 6236 18552 6267
rect 18782 6264 18788 6316
rect 18840 6264 18846 6316
rect 19720 6313 19748 6344
rect 20438 6332 20444 6384
rect 20496 6332 20502 6384
rect 22462 6372 22468 6384
rect 21100 6344 22468 6372
rect 19705 6307 19763 6313
rect 19705 6273 19717 6307
rect 19751 6273 19763 6307
rect 19705 6267 19763 6273
rect 19978 6264 19984 6316
rect 20036 6264 20042 6316
rect 21100 6313 21128 6344
rect 22462 6332 22468 6344
rect 22520 6372 22526 6384
rect 22925 6375 22983 6381
rect 22925 6372 22937 6375
rect 22520 6344 22937 6372
rect 22520 6332 22526 6344
rect 22925 6341 22937 6344
rect 22971 6341 22983 6375
rect 22925 6335 22983 6341
rect 21085 6307 21143 6313
rect 21085 6273 21097 6307
rect 21131 6273 21143 6307
rect 21085 6267 21143 6273
rect 21266 6264 21272 6316
rect 21324 6264 21330 6316
rect 22002 6264 22008 6316
rect 22060 6264 22066 6316
rect 22281 6307 22339 6313
rect 22281 6273 22293 6307
rect 22327 6304 22339 6307
rect 23198 6304 23204 6316
rect 22327 6276 23204 6304
rect 22327 6273 22339 6276
rect 22281 6267 22339 6273
rect 19150 6236 19156 6248
rect 18288 6208 19156 6236
rect 18288 6196 18294 6208
rect 19150 6196 19156 6208
rect 19208 6196 19214 6248
rect 19426 6196 19432 6248
rect 19484 6236 19490 6248
rect 19797 6239 19855 6245
rect 19797 6236 19809 6239
rect 19484 6208 19809 6236
rect 19484 6196 19490 6208
rect 19797 6205 19809 6208
rect 19843 6236 19855 6239
rect 20162 6236 20168 6248
rect 19843 6208 20168 6236
rect 19843 6205 19855 6208
rect 19797 6199 19855 6205
rect 20162 6196 20168 6208
rect 20220 6196 20226 6248
rect 20993 6239 21051 6245
rect 20993 6205 21005 6239
rect 21039 6205 21051 6239
rect 21284 6236 21312 6264
rect 22296 6236 22324 6267
rect 23198 6264 23204 6276
rect 23256 6264 23262 6316
rect 21284 6208 22324 6236
rect 20993 6199 21051 6205
rect 17494 6168 17500 6180
rect 15988 6140 17500 6168
rect 15988 6128 15994 6140
rect 17494 6128 17500 6140
rect 17552 6128 17558 6180
rect 18601 6171 18659 6177
rect 18601 6137 18613 6171
rect 18647 6168 18659 6171
rect 18966 6168 18972 6180
rect 18647 6140 18972 6168
rect 18647 6137 18659 6140
rect 18601 6131 18659 6137
rect 18966 6128 18972 6140
rect 19024 6128 19030 6180
rect 21008 6168 21036 6199
rect 23290 6196 23296 6248
rect 23348 6196 23354 6248
rect 21008 6140 22094 6168
rect 16666 6100 16672 6112
rect 15672 6072 16672 6100
rect 16666 6060 16672 6072
rect 16724 6060 16730 6112
rect 22066 6100 22094 6140
rect 22646 6100 22652 6112
rect 22066 6072 22652 6100
rect 22646 6060 22652 6072
rect 22704 6100 22710 6112
rect 22830 6100 22836 6112
rect 22704 6072 22836 6100
rect 22704 6060 22710 6072
rect 22830 6060 22836 6072
rect 22888 6100 22894 6112
rect 23109 6103 23167 6109
rect 23109 6100 23121 6103
rect 22888 6072 23121 6100
rect 22888 6060 22894 6072
rect 23109 6069 23121 6072
rect 23155 6069 23167 6103
rect 23109 6063 23167 6069
rect 1104 6010 23828 6032
rect 1104 5958 3790 6010
rect 3842 5958 3854 6010
rect 3906 5958 3918 6010
rect 3970 5958 3982 6010
rect 4034 5958 4046 6010
rect 4098 5958 9471 6010
rect 9523 5958 9535 6010
rect 9587 5958 9599 6010
rect 9651 5958 9663 6010
rect 9715 5958 9727 6010
rect 9779 5958 15152 6010
rect 15204 5958 15216 6010
rect 15268 5958 15280 6010
rect 15332 5958 15344 6010
rect 15396 5958 15408 6010
rect 15460 5958 20833 6010
rect 20885 5958 20897 6010
rect 20949 5958 20961 6010
rect 21013 5958 21025 6010
rect 21077 5958 21089 6010
rect 21141 5958 23828 6010
rect 1104 5936 23828 5958
rect 2130 5856 2136 5908
rect 2188 5856 2194 5908
rect 2222 5856 2228 5908
rect 2280 5896 2286 5908
rect 3973 5899 4031 5905
rect 3973 5896 3985 5899
rect 2280 5868 3985 5896
rect 2280 5856 2286 5868
rect 3973 5865 3985 5868
rect 4019 5865 4031 5899
rect 3973 5859 4031 5865
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 5592 5868 8156 5896
rect 5592 5856 5598 5868
rect 2682 5788 2688 5840
rect 2740 5828 2746 5840
rect 3050 5828 3056 5840
rect 2740 5800 3056 5828
rect 2740 5788 2746 5800
rect 3050 5788 3056 5800
rect 3108 5788 3114 5840
rect 3329 5831 3387 5837
rect 3329 5797 3341 5831
rect 3375 5828 3387 5831
rect 4338 5828 4344 5840
rect 3375 5800 4344 5828
rect 3375 5797 3387 5800
rect 3329 5791 3387 5797
rect 4338 5788 4344 5800
rect 4396 5788 4402 5840
rect 6362 5788 6368 5840
rect 6420 5828 6426 5840
rect 6420 5800 7236 5828
rect 6420 5788 6426 5800
rect 6092 5772 6144 5778
rect 2317 5763 2375 5769
rect 2317 5729 2329 5763
rect 2363 5760 2375 5763
rect 2363 5732 5028 5760
rect 2363 5729 2375 5732
rect 2317 5723 2375 5729
rect 2409 5695 2467 5701
rect 2409 5661 2421 5695
rect 2455 5661 2467 5695
rect 2409 5655 2467 5661
rect 2133 5627 2191 5633
rect 2133 5593 2145 5627
rect 2179 5624 2191 5627
rect 2222 5624 2228 5636
rect 2179 5596 2228 5624
rect 2179 5593 2191 5596
rect 2133 5587 2191 5593
rect 2222 5584 2228 5596
rect 2280 5584 2286 5636
rect 2424 5624 2452 5655
rect 2498 5652 2504 5704
rect 2556 5692 2562 5704
rect 3050 5692 3056 5704
rect 2556 5664 3056 5692
rect 2556 5652 2562 5664
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 3252 5701 3280 5732
rect 5000 5704 5028 5732
rect 7208 5760 7236 5800
rect 7926 5788 7932 5840
rect 7984 5828 7990 5840
rect 8128 5828 8156 5868
rect 8386 5856 8392 5908
rect 8444 5896 8450 5908
rect 9214 5896 9220 5908
rect 8444 5868 9220 5896
rect 8444 5856 8450 5868
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 11701 5899 11759 5905
rect 11701 5865 11713 5899
rect 11747 5896 11759 5899
rect 11974 5896 11980 5908
rect 11747 5868 11980 5896
rect 11747 5865 11759 5868
rect 11701 5859 11759 5865
rect 11974 5856 11980 5868
rect 12032 5856 12038 5908
rect 12158 5856 12164 5908
rect 12216 5896 12222 5908
rect 13357 5899 13415 5905
rect 13357 5896 13369 5899
rect 12216 5868 13369 5896
rect 12216 5856 12222 5868
rect 13357 5865 13369 5868
rect 13403 5865 13415 5899
rect 13357 5859 13415 5865
rect 14829 5899 14887 5905
rect 14829 5865 14841 5899
rect 14875 5896 14887 5899
rect 15930 5896 15936 5908
rect 14875 5868 15936 5896
rect 14875 5865 14887 5868
rect 14829 5859 14887 5865
rect 15930 5856 15936 5868
rect 15988 5856 15994 5908
rect 16390 5856 16396 5908
rect 16448 5896 16454 5908
rect 18782 5896 18788 5908
rect 16448 5868 18788 5896
rect 16448 5856 16454 5868
rect 18782 5856 18788 5868
rect 18840 5856 18846 5908
rect 19886 5856 19892 5908
rect 19944 5896 19950 5908
rect 21266 5896 21272 5908
rect 19944 5868 21272 5896
rect 19944 5856 19950 5868
rect 21266 5856 21272 5868
rect 21324 5856 21330 5908
rect 21913 5899 21971 5905
rect 21913 5865 21925 5899
rect 21959 5896 21971 5899
rect 22462 5896 22468 5908
rect 21959 5868 22468 5896
rect 21959 5865 21971 5868
rect 21913 5859 21971 5865
rect 22462 5856 22468 5868
rect 22520 5856 22526 5908
rect 8294 5828 8300 5840
rect 7984 5800 8064 5828
rect 7984 5788 7990 5800
rect 8036 5769 8064 5800
rect 8128 5800 8300 5828
rect 8128 5769 8156 5800
rect 8294 5788 8300 5800
rect 8352 5788 8358 5840
rect 8478 5788 8484 5840
rect 8536 5828 8542 5840
rect 9582 5828 9588 5840
rect 8536 5800 9588 5828
rect 8536 5788 8542 5800
rect 9582 5788 9588 5800
rect 9640 5788 9646 5840
rect 11330 5788 11336 5840
rect 11388 5828 11394 5840
rect 11790 5828 11796 5840
rect 11388 5800 11796 5828
rect 11388 5788 11394 5800
rect 11790 5788 11796 5800
rect 11848 5788 11854 5840
rect 11882 5788 11888 5840
rect 11940 5828 11946 5840
rect 12345 5831 12403 5837
rect 12345 5828 12357 5831
rect 11940 5800 12357 5828
rect 11940 5788 11946 5800
rect 12345 5797 12357 5800
rect 12391 5797 12403 5831
rect 20070 5828 20076 5840
rect 12345 5791 12403 5797
rect 12728 5800 20076 5828
rect 8021 5763 8079 5769
rect 6144 5732 7144 5760
rect 7208 5732 7972 5760
rect 6092 5714 6144 5720
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5661 3295 5695
rect 3237 5655 3295 5661
rect 4154 5652 4160 5704
rect 4212 5652 4218 5704
rect 4430 5652 4436 5704
rect 4488 5692 4494 5704
rect 4706 5692 4712 5704
rect 4488 5664 4712 5692
rect 4488 5652 4494 5664
rect 4706 5652 4712 5664
rect 4764 5692 4770 5704
rect 4801 5695 4859 5701
rect 4801 5692 4813 5695
rect 4764 5664 4813 5692
rect 4764 5652 4770 5664
rect 4801 5661 4813 5664
rect 4847 5661 4859 5695
rect 4801 5655 4859 5661
rect 4982 5652 4988 5704
rect 5040 5692 5046 5704
rect 5169 5695 5227 5701
rect 5169 5692 5181 5695
rect 5040 5664 5181 5692
rect 5040 5652 5046 5664
rect 5169 5661 5181 5664
rect 5215 5661 5227 5695
rect 5169 5655 5227 5661
rect 5997 5695 6055 5701
rect 5997 5661 6009 5695
rect 6043 5661 6055 5695
rect 5997 5655 6055 5661
rect 2866 5624 2872 5636
rect 2424 5596 2872 5624
rect 2866 5584 2872 5596
rect 2924 5584 2930 5636
rect 3602 5584 3608 5636
rect 3660 5624 3666 5636
rect 4341 5627 4399 5633
rect 4341 5624 4353 5627
rect 3660 5596 4353 5624
rect 3660 5584 3666 5596
rect 4341 5593 4353 5596
rect 4387 5593 4399 5627
rect 4341 5587 4399 5593
rect 1673 5559 1731 5565
rect 1673 5525 1685 5559
rect 1719 5556 1731 5559
rect 2038 5556 2044 5568
rect 1719 5528 2044 5556
rect 1719 5525 1731 5528
rect 1673 5519 1731 5525
rect 2038 5516 2044 5528
rect 2096 5556 2102 5568
rect 2406 5556 2412 5568
rect 2096 5528 2412 5556
rect 2096 5516 2102 5528
rect 2406 5516 2412 5528
rect 2464 5516 2470 5568
rect 2593 5559 2651 5565
rect 2593 5525 2605 5559
rect 2639 5556 2651 5559
rect 3234 5556 3240 5568
rect 2639 5528 3240 5556
rect 2639 5525 2651 5528
rect 2593 5519 2651 5525
rect 3234 5516 3240 5528
rect 3292 5556 3298 5568
rect 4062 5556 4068 5568
rect 3292 5528 4068 5556
rect 3292 5516 3298 5528
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 4356 5556 4384 5587
rect 5534 5584 5540 5636
rect 5592 5624 5598 5636
rect 6012 5624 6040 5655
rect 6546 5652 6552 5704
rect 6604 5692 6610 5704
rect 7009 5695 7067 5701
rect 7009 5692 7021 5695
rect 6604 5664 7021 5692
rect 6604 5652 6610 5664
rect 7009 5661 7021 5664
rect 7055 5661 7067 5695
rect 7009 5655 7067 5661
rect 6638 5624 6644 5636
rect 5592 5596 6644 5624
rect 5592 5584 5598 5596
rect 6638 5584 6644 5596
rect 6696 5584 6702 5636
rect 5626 5556 5632 5568
rect 4356 5528 5632 5556
rect 5626 5516 5632 5528
rect 5684 5516 5690 5568
rect 5718 5516 5724 5568
rect 5776 5565 5782 5568
rect 5776 5559 5805 5565
rect 5793 5525 5805 5559
rect 5776 5519 5805 5525
rect 5776 5516 5782 5519
rect 6454 5516 6460 5568
rect 6512 5556 6518 5568
rect 6822 5556 6828 5568
rect 6512 5528 6828 5556
rect 6512 5516 6518 5528
rect 6822 5516 6828 5528
rect 6880 5516 6886 5568
rect 6917 5559 6975 5565
rect 6917 5525 6929 5559
rect 6963 5556 6975 5559
rect 7116 5556 7144 5732
rect 7944 5701 7972 5732
rect 8021 5729 8033 5763
rect 8067 5729 8079 5763
rect 8021 5723 8079 5729
rect 8113 5763 8171 5769
rect 8113 5729 8125 5763
rect 8159 5729 8171 5763
rect 8113 5723 8171 5729
rect 8202 5720 8208 5772
rect 8260 5720 8266 5772
rect 8389 5763 8447 5769
rect 8389 5729 8401 5763
rect 8435 5729 8447 5763
rect 8389 5723 8447 5729
rect 10137 5763 10195 5769
rect 10137 5729 10149 5763
rect 10183 5760 10195 5763
rect 10183 5732 11284 5760
rect 10183 5729 10195 5732
rect 10137 5723 10195 5729
rect 7929 5695 7987 5701
rect 7929 5661 7941 5695
rect 7975 5692 7987 5695
rect 8294 5692 8300 5704
rect 7975 5664 8300 5692
rect 7975 5661 7987 5664
rect 7929 5655 7987 5661
rect 8294 5652 8300 5664
rect 8352 5652 8358 5704
rect 8404 5692 8432 5723
rect 10321 5695 10379 5701
rect 10321 5692 10333 5695
rect 8404 5664 10333 5692
rect 10321 5661 10333 5664
rect 10367 5692 10379 5695
rect 10502 5692 10508 5704
rect 10367 5664 10508 5692
rect 10367 5661 10379 5664
rect 10321 5655 10379 5661
rect 10502 5652 10508 5664
rect 10560 5652 10566 5704
rect 10594 5652 10600 5704
rect 10652 5652 10658 5704
rect 11054 5652 11060 5704
rect 11112 5652 11118 5704
rect 11256 5701 11284 5732
rect 12250 5720 12256 5772
rect 12308 5760 12314 5772
rect 12728 5769 12756 5800
rect 20070 5788 20076 5800
rect 20128 5788 20134 5840
rect 20162 5788 20168 5840
rect 20220 5788 20226 5840
rect 12713 5763 12771 5769
rect 12713 5760 12725 5763
rect 12308 5732 12725 5760
rect 12308 5720 12314 5732
rect 12713 5729 12725 5732
rect 12759 5729 12771 5763
rect 12713 5723 12771 5729
rect 12805 5763 12863 5769
rect 12805 5729 12817 5763
rect 12851 5760 12863 5763
rect 13630 5760 13636 5772
rect 12851 5732 13636 5760
rect 12851 5729 12863 5732
rect 12805 5723 12863 5729
rect 13630 5720 13636 5732
rect 13688 5720 13694 5772
rect 17126 5760 17132 5772
rect 15120 5732 17132 5760
rect 15120 5704 15148 5732
rect 17126 5720 17132 5732
rect 17184 5760 17190 5772
rect 17184 5732 17264 5760
rect 17184 5720 17190 5732
rect 11241 5695 11299 5701
rect 11241 5661 11253 5695
rect 11287 5661 11299 5695
rect 11241 5655 11299 5661
rect 11330 5652 11336 5704
rect 11388 5652 11394 5704
rect 11422 5652 11428 5704
rect 11480 5652 11486 5704
rect 12529 5695 12587 5701
rect 12529 5661 12541 5695
rect 12575 5661 12587 5695
rect 12529 5655 12587 5661
rect 12621 5695 12679 5701
rect 12621 5661 12633 5695
rect 12667 5661 12679 5695
rect 12621 5655 12679 5661
rect 7193 5627 7251 5633
rect 7193 5593 7205 5627
rect 7239 5624 7251 5627
rect 11698 5624 11704 5636
rect 7239 5596 11704 5624
rect 7239 5593 7251 5596
rect 7193 5587 7251 5593
rect 11698 5584 11704 5596
rect 11756 5584 11762 5636
rect 6963 5528 7144 5556
rect 10505 5559 10563 5565
rect 6963 5525 6975 5528
rect 6917 5519 6975 5525
rect 10505 5525 10517 5559
rect 10551 5556 10563 5559
rect 11790 5556 11796 5568
rect 10551 5528 11796 5556
rect 10551 5525 10563 5528
rect 10505 5519 10563 5525
rect 11790 5516 11796 5528
rect 11848 5516 11854 5568
rect 12544 5556 12572 5655
rect 12636 5624 12664 5655
rect 13354 5652 13360 5704
rect 13412 5652 13418 5704
rect 13541 5695 13599 5701
rect 13541 5661 13553 5695
rect 13587 5692 13599 5695
rect 14734 5692 14740 5704
rect 13587 5664 14740 5692
rect 13587 5661 13599 5664
rect 13541 5655 13599 5661
rect 14734 5652 14740 5664
rect 14792 5652 14798 5704
rect 15102 5652 15108 5704
rect 15160 5652 15166 5704
rect 15565 5695 15623 5701
rect 15565 5661 15577 5695
rect 15611 5692 15623 5695
rect 16022 5692 16028 5704
rect 15611 5664 16028 5692
rect 15611 5661 15623 5664
rect 15565 5655 15623 5661
rect 16022 5652 16028 5664
rect 16080 5652 16086 5704
rect 16298 5652 16304 5704
rect 16356 5692 16362 5704
rect 16574 5692 16580 5704
rect 16356 5664 16580 5692
rect 16356 5652 16362 5664
rect 16574 5652 16580 5664
rect 16632 5652 16638 5704
rect 16942 5652 16948 5704
rect 17000 5692 17006 5704
rect 17236 5701 17264 5732
rect 17494 5720 17500 5772
rect 17552 5720 17558 5772
rect 18230 5720 18236 5772
rect 18288 5720 18294 5772
rect 19521 5763 19579 5769
rect 19521 5729 19533 5763
rect 19567 5760 19579 5763
rect 19794 5760 19800 5772
rect 19567 5732 19800 5760
rect 19567 5729 19579 5732
rect 19521 5723 19579 5729
rect 19794 5720 19800 5732
rect 19852 5760 19858 5772
rect 19852 5732 20392 5760
rect 19852 5720 19858 5732
rect 17037 5695 17095 5701
rect 17037 5692 17049 5695
rect 17000 5664 17049 5692
rect 17000 5652 17006 5664
rect 17037 5661 17049 5664
rect 17083 5661 17095 5695
rect 17037 5655 17095 5661
rect 17221 5695 17279 5701
rect 17221 5661 17233 5695
rect 17267 5661 17279 5695
rect 17221 5655 17279 5661
rect 17310 5652 17316 5704
rect 17368 5692 17374 5704
rect 17589 5695 17647 5701
rect 17589 5692 17601 5695
rect 17368 5664 17601 5692
rect 17368 5652 17374 5664
rect 17589 5661 17601 5664
rect 17635 5661 17647 5695
rect 17589 5655 17647 5661
rect 19610 5652 19616 5704
rect 19668 5692 19674 5704
rect 20364 5701 20392 5732
rect 20622 5720 20628 5772
rect 20680 5720 20686 5772
rect 22278 5720 22284 5772
rect 22336 5720 22342 5772
rect 22922 5720 22928 5772
rect 22980 5720 22986 5772
rect 20073 5695 20131 5701
rect 20073 5692 20085 5695
rect 19668 5664 20085 5692
rect 19668 5652 19674 5664
rect 20073 5661 20085 5664
rect 20119 5661 20131 5695
rect 20073 5655 20131 5661
rect 20349 5695 20407 5701
rect 20349 5661 20361 5695
rect 20395 5692 20407 5695
rect 20395 5664 20668 5692
rect 20395 5661 20407 5664
rect 20349 5655 20407 5661
rect 14918 5624 14924 5636
rect 12636 5596 14924 5624
rect 14918 5584 14924 5596
rect 14976 5584 14982 5636
rect 15013 5627 15071 5633
rect 15013 5593 15025 5627
rect 15059 5593 15071 5627
rect 15838 5624 15844 5636
rect 15013 5587 15071 5593
rect 15672 5596 15844 5624
rect 12710 5556 12716 5568
rect 12544 5528 12716 5556
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 15028 5556 15056 5587
rect 15672 5556 15700 5596
rect 15838 5584 15844 5596
rect 15896 5624 15902 5636
rect 17328 5624 17356 5652
rect 20640 5636 20668 5664
rect 22094 5652 22100 5704
rect 22152 5652 22158 5704
rect 22554 5652 22560 5704
rect 22612 5692 22618 5704
rect 22741 5695 22799 5701
rect 22741 5692 22753 5695
rect 22612 5664 22753 5692
rect 22612 5652 22618 5664
rect 22741 5661 22753 5664
rect 22787 5661 22799 5695
rect 22741 5655 22799 5661
rect 15896 5596 17356 5624
rect 15896 5584 15902 5596
rect 20622 5584 20628 5636
rect 20680 5584 20686 5636
rect 15028 5528 15700 5556
rect 1104 5466 23987 5488
rect 1104 5414 6630 5466
rect 6682 5414 6694 5466
rect 6746 5414 6758 5466
rect 6810 5414 6822 5466
rect 6874 5414 6886 5466
rect 6938 5414 12311 5466
rect 12363 5414 12375 5466
rect 12427 5414 12439 5466
rect 12491 5414 12503 5466
rect 12555 5414 12567 5466
rect 12619 5414 17992 5466
rect 18044 5414 18056 5466
rect 18108 5414 18120 5466
rect 18172 5414 18184 5466
rect 18236 5414 18248 5466
rect 18300 5414 23673 5466
rect 23725 5414 23737 5466
rect 23789 5414 23801 5466
rect 23853 5414 23865 5466
rect 23917 5414 23929 5466
rect 23981 5414 23987 5466
rect 1104 5392 23987 5414
rect 2593 5355 2651 5361
rect 2593 5321 2605 5355
rect 2639 5352 2651 5355
rect 4614 5352 4620 5364
rect 2639 5324 4620 5352
rect 2639 5321 2651 5324
rect 2593 5315 2651 5321
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 6362 5312 6368 5364
rect 6420 5352 6426 5364
rect 6420 5324 6776 5352
rect 6420 5312 6426 5324
rect 2498 5284 2504 5296
rect 2332 5256 2504 5284
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5185 2099 5219
rect 2041 5179 2099 5185
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5216 2191 5219
rect 2222 5216 2228 5228
rect 2179 5188 2228 5216
rect 2179 5185 2191 5188
rect 2133 5179 2191 5185
rect 2056 5148 2084 5179
rect 2222 5176 2228 5188
rect 2280 5176 2286 5228
rect 2332 5225 2360 5256
rect 2498 5244 2504 5256
rect 2556 5244 2562 5296
rect 3694 5284 3700 5296
rect 3068 5256 3700 5284
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5185 2375 5219
rect 2317 5179 2375 5185
rect 2409 5219 2467 5225
rect 2409 5185 2421 5219
rect 2455 5216 2467 5219
rect 3068 5216 3096 5256
rect 3694 5244 3700 5256
rect 3752 5244 3758 5296
rect 4062 5244 4068 5296
rect 4120 5284 4126 5296
rect 4120 5256 6592 5284
rect 4120 5244 4126 5256
rect 2455 5188 3096 5216
rect 2455 5185 2467 5188
rect 2409 5179 2467 5185
rect 3142 5176 3148 5228
rect 3200 5216 3206 5228
rect 3237 5219 3295 5225
rect 3237 5216 3249 5219
rect 3200 5188 3249 5216
rect 3200 5176 3206 5188
rect 3237 5185 3249 5188
rect 3283 5216 3295 5219
rect 4157 5219 4215 5225
rect 3283 5188 4108 5216
rect 3283 5185 3295 5188
rect 3237 5179 3295 5185
rect 2682 5148 2688 5160
rect 2056 5120 2688 5148
rect 2682 5108 2688 5120
rect 2740 5108 2746 5160
rect 2866 5108 2872 5160
rect 2924 5148 2930 5160
rect 3510 5148 3516 5160
rect 2924 5120 3516 5148
rect 2924 5108 2930 5120
rect 3510 5108 3516 5120
rect 3568 5108 3574 5160
rect 4080 5080 4108 5188
rect 4157 5185 4169 5219
rect 4203 5216 4215 5219
rect 4522 5216 4528 5228
rect 4203 5188 4528 5216
rect 4203 5185 4215 5188
rect 4157 5179 4215 5185
rect 4522 5176 4528 5188
rect 4580 5216 4586 5228
rect 5074 5216 5080 5228
rect 4580 5188 5080 5216
rect 4580 5176 4586 5188
rect 5074 5176 5080 5188
rect 5132 5176 5138 5228
rect 5537 5219 5595 5225
rect 5537 5185 5549 5219
rect 5583 5216 5595 5219
rect 5810 5216 5816 5228
rect 5583 5188 5816 5216
rect 5583 5185 5595 5188
rect 5537 5179 5595 5185
rect 5810 5176 5816 5188
rect 5868 5176 5874 5228
rect 6564 5225 6592 5256
rect 6748 5225 6776 5324
rect 11330 5312 11336 5364
rect 11388 5352 11394 5364
rect 12437 5355 12495 5361
rect 12437 5352 12449 5355
rect 11388 5324 12449 5352
rect 11388 5312 11394 5324
rect 12437 5321 12449 5324
rect 12483 5321 12495 5355
rect 12437 5315 12495 5321
rect 12710 5312 12716 5364
rect 12768 5312 12774 5364
rect 13262 5312 13268 5364
rect 13320 5352 13326 5364
rect 14369 5355 14427 5361
rect 14369 5352 14381 5355
rect 13320 5324 14381 5352
rect 13320 5312 13326 5324
rect 14369 5321 14381 5324
rect 14415 5352 14427 5355
rect 14734 5352 14740 5364
rect 14415 5324 14740 5352
rect 14415 5321 14427 5324
rect 14369 5315 14427 5321
rect 14734 5312 14740 5324
rect 14792 5312 14798 5364
rect 14918 5312 14924 5364
rect 14976 5352 14982 5364
rect 15013 5355 15071 5361
rect 15013 5352 15025 5355
rect 14976 5324 15025 5352
rect 14976 5312 14982 5324
rect 15013 5321 15025 5324
rect 15059 5321 15071 5355
rect 15013 5315 15071 5321
rect 15470 5312 15476 5364
rect 15528 5312 15534 5364
rect 16209 5355 16267 5361
rect 16209 5321 16221 5355
rect 16255 5352 16267 5355
rect 16298 5352 16304 5364
rect 16255 5324 16304 5352
rect 16255 5321 16267 5324
rect 16209 5315 16267 5321
rect 16298 5312 16304 5324
rect 16356 5312 16362 5364
rect 16850 5312 16856 5364
rect 16908 5352 16914 5364
rect 17129 5355 17187 5361
rect 17129 5352 17141 5355
rect 16908 5324 17141 5352
rect 16908 5312 16914 5324
rect 17129 5321 17141 5324
rect 17175 5321 17187 5355
rect 17129 5315 17187 5321
rect 19242 5312 19248 5364
rect 19300 5312 19306 5364
rect 19978 5312 19984 5364
rect 20036 5352 20042 5364
rect 20441 5355 20499 5361
rect 20441 5352 20453 5355
rect 20036 5324 20453 5352
rect 20036 5312 20042 5324
rect 20441 5321 20453 5324
rect 20487 5321 20499 5355
rect 20441 5315 20499 5321
rect 7098 5244 7104 5296
rect 7156 5284 7162 5296
rect 7156 5256 8892 5284
rect 7156 5244 7162 5256
rect 8864 5228 8892 5256
rect 9214 5244 9220 5296
rect 9272 5284 9278 5296
rect 10965 5287 11023 5293
rect 9272 5256 10456 5284
rect 9272 5244 9278 5256
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 6733 5219 6791 5225
rect 6733 5185 6745 5219
rect 6779 5185 6791 5219
rect 6733 5179 6791 5185
rect 7006 5176 7012 5228
rect 7064 5216 7070 5228
rect 8021 5219 8079 5225
rect 8021 5216 8033 5219
rect 7064 5188 8033 5216
rect 7064 5176 7070 5188
rect 8021 5185 8033 5188
rect 8067 5185 8079 5219
rect 8021 5179 8079 5185
rect 8294 5176 8300 5228
rect 8352 5216 8358 5228
rect 8665 5219 8723 5225
rect 8665 5216 8677 5219
rect 8352 5188 8677 5216
rect 8352 5176 8358 5188
rect 8665 5185 8677 5188
rect 8711 5185 8723 5219
rect 8665 5179 8723 5185
rect 8846 5176 8852 5228
rect 8904 5216 8910 5228
rect 9401 5219 9459 5225
rect 9401 5216 9413 5219
rect 8904 5188 9413 5216
rect 8904 5176 8910 5188
rect 9401 5185 9413 5188
rect 9447 5185 9459 5219
rect 9677 5219 9735 5225
rect 9677 5216 9689 5219
rect 9401 5179 9459 5185
rect 9508 5188 9689 5216
rect 4982 5108 4988 5160
rect 5040 5108 5046 5160
rect 5718 5108 5724 5160
rect 5776 5108 5782 5160
rect 6086 5108 6092 5160
rect 6144 5148 6150 5160
rect 7745 5151 7803 5157
rect 7745 5148 7757 5151
rect 6144 5120 7757 5148
rect 6144 5108 6150 5120
rect 7745 5117 7757 5120
rect 7791 5117 7803 5151
rect 7745 5111 7803 5117
rect 6914 5080 6920 5092
rect 4080 5052 6920 5080
rect 6914 5040 6920 5052
rect 6972 5040 6978 5092
rect 6638 4972 6644 5024
rect 6696 4972 6702 5024
rect 7760 5012 7788 5111
rect 8570 5108 8576 5160
rect 8628 5148 8634 5160
rect 9508 5148 9536 5188
rect 9677 5185 9689 5188
rect 9723 5185 9735 5219
rect 9677 5179 9735 5185
rect 9769 5219 9827 5225
rect 9769 5185 9781 5219
rect 9815 5216 9827 5219
rect 9858 5216 9864 5228
rect 9815 5188 9864 5216
rect 9815 5185 9827 5188
rect 9769 5179 9827 5185
rect 9858 5176 9864 5188
rect 9916 5176 9922 5228
rect 10428 5225 10456 5256
rect 10965 5253 10977 5287
rect 11011 5284 11023 5287
rect 12728 5284 12756 5312
rect 11011 5256 12756 5284
rect 11011 5253 11023 5256
rect 10965 5247 11023 5253
rect 15286 5244 15292 5296
rect 15344 5244 15350 5296
rect 15381 5287 15439 5293
rect 15381 5253 15393 5287
rect 15427 5284 15439 5287
rect 15488 5284 15516 5312
rect 15427 5256 15516 5284
rect 15427 5253 15439 5256
rect 15381 5247 15439 5253
rect 16942 5244 16948 5296
rect 17000 5284 17006 5296
rect 17281 5287 17339 5293
rect 17281 5284 17293 5287
rect 17000 5256 17293 5284
rect 17000 5244 17006 5256
rect 17281 5253 17293 5256
rect 17327 5253 17339 5287
rect 17281 5247 17339 5253
rect 17494 5244 17500 5296
rect 17552 5244 17558 5296
rect 20456 5284 20484 5315
rect 21174 5312 21180 5364
rect 21232 5312 21238 5364
rect 22281 5355 22339 5361
rect 22281 5321 22293 5355
rect 22327 5352 22339 5355
rect 22830 5352 22836 5364
rect 22327 5324 22836 5352
rect 22327 5321 22339 5324
rect 22281 5315 22339 5321
rect 22830 5312 22836 5324
rect 22888 5312 22894 5364
rect 20456 5256 21128 5284
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5185 10011 5219
rect 9953 5179 10011 5185
rect 10413 5219 10471 5225
rect 10413 5185 10425 5219
rect 10459 5185 10471 5219
rect 10413 5179 10471 5185
rect 8628 5120 9536 5148
rect 8628 5108 8634 5120
rect 9582 5108 9588 5160
rect 9640 5108 9646 5160
rect 8018 5040 8024 5092
rect 8076 5080 8082 5092
rect 8481 5083 8539 5089
rect 8481 5080 8493 5083
rect 8076 5052 8493 5080
rect 8076 5040 8082 5052
rect 8481 5049 8493 5052
rect 8527 5049 8539 5083
rect 9968 5080 9996 5179
rect 10502 5176 10508 5228
rect 10560 5176 10566 5228
rect 10686 5176 10692 5228
rect 10744 5176 10750 5228
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5216 10839 5219
rect 10870 5216 10876 5228
rect 10827 5188 10876 5216
rect 10827 5185 10839 5188
rect 10781 5179 10839 5185
rect 10870 5176 10876 5188
rect 10928 5176 10934 5228
rect 11790 5176 11796 5228
rect 11848 5216 11854 5228
rect 11974 5216 11980 5228
rect 11848 5188 11980 5216
rect 11848 5176 11854 5188
rect 11974 5176 11980 5188
rect 12032 5216 12038 5228
rect 12621 5219 12679 5225
rect 12621 5216 12633 5219
rect 12032 5188 12633 5216
rect 12032 5176 12038 5188
rect 12621 5185 12633 5188
rect 12667 5185 12679 5219
rect 12621 5179 12679 5185
rect 12710 5176 12716 5228
rect 12768 5176 12774 5228
rect 12802 5176 12808 5228
rect 12860 5176 12866 5228
rect 12894 5176 12900 5228
rect 12952 5216 12958 5228
rect 12989 5219 13047 5225
rect 12989 5216 13001 5219
rect 12952 5188 13001 5216
rect 12952 5176 12958 5188
rect 12989 5185 13001 5188
rect 13035 5185 13047 5219
rect 12989 5179 13047 5185
rect 13998 5176 14004 5228
rect 14056 5216 14062 5228
rect 14642 5216 14648 5228
rect 14056 5188 14648 5216
rect 14056 5176 14062 5188
rect 14642 5176 14648 5188
rect 14700 5216 14706 5228
rect 15151 5219 15209 5225
rect 15151 5216 15163 5219
rect 14700 5188 15163 5216
rect 14700 5176 14706 5188
rect 15151 5185 15163 5188
rect 15197 5185 15209 5219
rect 15151 5179 15209 5185
rect 15470 5176 15476 5228
rect 15528 5216 15534 5228
rect 15564 5219 15622 5225
rect 15564 5216 15576 5219
rect 15528 5188 15576 5216
rect 15528 5176 15534 5188
rect 15564 5185 15576 5188
rect 15610 5185 15622 5219
rect 15564 5179 15622 5185
rect 15657 5219 15715 5225
rect 15657 5185 15669 5219
rect 15703 5216 15715 5219
rect 15838 5216 15844 5228
rect 15703 5188 15844 5216
rect 15703 5185 15715 5188
rect 15657 5179 15715 5185
rect 15838 5176 15844 5188
rect 15896 5176 15902 5228
rect 18138 5176 18144 5228
rect 18196 5176 18202 5228
rect 18233 5219 18291 5225
rect 18233 5185 18245 5219
rect 18279 5216 18291 5219
rect 18322 5216 18328 5228
rect 18279 5188 18328 5216
rect 18279 5185 18291 5188
rect 18233 5179 18291 5185
rect 18322 5176 18328 5188
rect 18380 5176 18386 5228
rect 18414 5176 18420 5228
rect 18472 5176 18478 5228
rect 19613 5219 19671 5225
rect 19613 5185 19625 5219
rect 19659 5216 19671 5219
rect 20254 5216 20260 5228
rect 19659 5188 20260 5216
rect 19659 5185 19671 5188
rect 19613 5179 19671 5185
rect 20254 5176 20260 5188
rect 20312 5176 20318 5228
rect 20533 5219 20591 5225
rect 20533 5185 20545 5219
rect 20579 5216 20591 5219
rect 20622 5216 20628 5228
rect 20579 5188 20628 5216
rect 20579 5185 20591 5188
rect 20533 5179 20591 5185
rect 20622 5176 20628 5188
rect 20680 5176 20686 5228
rect 21100 5225 21128 5256
rect 22094 5244 22100 5296
rect 22152 5284 22158 5296
rect 22922 5284 22928 5296
rect 22152 5256 22928 5284
rect 22152 5244 22158 5256
rect 22922 5244 22928 5256
rect 22980 5284 22986 5296
rect 23017 5287 23075 5293
rect 23017 5284 23029 5287
rect 22980 5256 23029 5284
rect 22980 5244 22986 5256
rect 23017 5253 23029 5256
rect 23063 5253 23075 5287
rect 23017 5247 23075 5253
rect 21085 5219 21143 5225
rect 21085 5185 21097 5219
rect 21131 5185 21143 5219
rect 21085 5179 21143 5185
rect 21266 5176 21272 5228
rect 21324 5176 21330 5228
rect 22741 5219 22799 5225
rect 22741 5185 22753 5219
rect 22787 5216 22799 5219
rect 22830 5216 22836 5228
rect 22787 5188 22836 5216
rect 22787 5185 22799 5188
rect 22741 5179 22799 5185
rect 22830 5176 22836 5188
rect 22888 5176 22894 5228
rect 19705 5151 19763 5157
rect 19705 5117 19717 5151
rect 19751 5148 19763 5151
rect 20438 5148 20444 5160
rect 19751 5120 20444 5148
rect 19751 5117 19763 5120
rect 19705 5111 19763 5117
rect 20438 5108 20444 5120
rect 20496 5108 20502 5160
rect 8481 5043 8539 5049
rect 8680 5052 9996 5080
rect 8680 5012 8708 5052
rect 12894 5040 12900 5092
rect 12952 5080 12958 5092
rect 15470 5080 15476 5092
rect 12952 5052 15476 5080
rect 12952 5040 12958 5052
rect 15470 5040 15476 5052
rect 15528 5040 15534 5092
rect 17494 5080 17500 5092
rect 15672 5052 17500 5080
rect 7760 4984 8708 5012
rect 8754 4972 8760 5024
rect 8812 5012 8818 5024
rect 9217 5015 9275 5021
rect 9217 5012 9229 5015
rect 8812 4984 9229 5012
rect 8812 4972 8818 4984
rect 9217 4981 9229 4984
rect 9263 4981 9275 5015
rect 9217 4975 9275 4981
rect 13354 4972 13360 5024
rect 13412 5012 13418 5024
rect 13541 5015 13599 5021
rect 13541 5012 13553 5015
rect 13412 4984 13553 5012
rect 13412 4972 13418 4984
rect 13541 4981 13553 4984
rect 13587 5012 13599 5015
rect 13630 5012 13636 5024
rect 13587 4984 13636 5012
rect 13587 4981 13599 4984
rect 13541 4975 13599 4981
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 13906 4972 13912 5024
rect 13964 5012 13970 5024
rect 15286 5012 15292 5024
rect 13964 4984 15292 5012
rect 13964 4972 13970 4984
rect 15286 4972 15292 4984
rect 15344 5012 15350 5024
rect 15672 5012 15700 5052
rect 17494 5040 17500 5052
rect 17552 5040 17558 5092
rect 18601 5083 18659 5089
rect 18601 5049 18613 5083
rect 18647 5080 18659 5083
rect 19794 5080 19800 5092
rect 18647 5052 19800 5080
rect 18647 5049 18659 5052
rect 18601 5043 18659 5049
rect 19794 5040 19800 5052
rect 19852 5040 19858 5092
rect 15344 4984 15700 5012
rect 15344 4972 15350 4984
rect 17310 4972 17316 5024
rect 17368 4972 17374 5024
rect 1104 4922 23828 4944
rect 1104 4870 3790 4922
rect 3842 4870 3854 4922
rect 3906 4870 3918 4922
rect 3970 4870 3982 4922
rect 4034 4870 4046 4922
rect 4098 4870 9471 4922
rect 9523 4870 9535 4922
rect 9587 4870 9599 4922
rect 9651 4870 9663 4922
rect 9715 4870 9727 4922
rect 9779 4870 15152 4922
rect 15204 4870 15216 4922
rect 15268 4870 15280 4922
rect 15332 4870 15344 4922
rect 15396 4870 15408 4922
rect 15460 4870 20833 4922
rect 20885 4870 20897 4922
rect 20949 4870 20961 4922
rect 21013 4870 21025 4922
rect 21077 4870 21089 4922
rect 21141 4870 23828 4922
rect 1104 4848 23828 4870
rect 5721 4811 5779 4817
rect 5721 4777 5733 4811
rect 5767 4808 5779 4811
rect 7742 4808 7748 4820
rect 5767 4780 7748 4808
rect 5767 4777 5779 4780
rect 5721 4771 5779 4777
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 9122 4768 9128 4820
rect 9180 4808 9186 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 9180 4780 9413 4808
rect 9180 4768 9186 4780
rect 9401 4777 9413 4780
rect 9447 4777 9459 4811
rect 9401 4771 9459 4777
rect 11149 4811 11207 4817
rect 11149 4777 11161 4811
rect 11195 4808 11207 4811
rect 11514 4808 11520 4820
rect 11195 4780 11520 4808
rect 11195 4777 11207 4780
rect 11149 4771 11207 4777
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 12066 4768 12072 4820
rect 12124 4768 12130 4820
rect 12158 4768 12164 4820
rect 12216 4808 12222 4820
rect 12710 4808 12716 4820
rect 12216 4780 12716 4808
rect 12216 4768 12222 4780
rect 12710 4768 12716 4780
rect 12768 4808 12774 4820
rect 13906 4808 13912 4820
rect 12768 4780 13912 4808
rect 12768 4768 12774 4780
rect 13906 4768 13912 4780
rect 13964 4768 13970 4820
rect 15010 4768 15016 4820
rect 15068 4768 15074 4820
rect 15562 4768 15568 4820
rect 15620 4768 15626 4820
rect 15930 4768 15936 4820
rect 15988 4808 15994 4820
rect 16574 4808 16580 4820
rect 15988 4780 16580 4808
rect 15988 4768 15994 4780
rect 16574 4768 16580 4780
rect 16632 4768 16638 4820
rect 16758 4768 16764 4820
rect 16816 4808 16822 4820
rect 17313 4811 17371 4817
rect 17313 4808 17325 4811
rect 16816 4780 17325 4808
rect 16816 4768 16822 4780
rect 17313 4777 17325 4780
rect 17359 4777 17371 4811
rect 17313 4771 17371 4777
rect 18138 4768 18144 4820
rect 18196 4808 18202 4820
rect 19797 4811 19855 4817
rect 19797 4808 19809 4811
rect 18196 4780 19809 4808
rect 18196 4768 18202 4780
rect 19797 4777 19809 4780
rect 19843 4777 19855 4811
rect 19797 4771 19855 4777
rect 20254 4768 20260 4820
rect 20312 4768 20318 4820
rect 20622 4768 20628 4820
rect 20680 4808 20686 4820
rect 20809 4811 20867 4817
rect 20809 4808 20821 4811
rect 20680 4780 20821 4808
rect 20680 4768 20686 4780
rect 20809 4777 20821 4780
rect 20855 4777 20867 4811
rect 20809 4771 20867 4777
rect 5626 4700 5632 4752
rect 5684 4740 5690 4752
rect 7098 4740 7104 4752
rect 5684 4712 7104 4740
rect 5684 4700 5690 4712
rect 7098 4700 7104 4712
rect 7156 4700 7162 4752
rect 8202 4700 8208 4752
rect 8260 4740 8266 4752
rect 12894 4740 12900 4752
rect 8260 4712 12900 4740
rect 8260 4700 8266 4712
rect 12894 4700 12900 4712
rect 12952 4700 12958 4752
rect 13630 4700 13636 4752
rect 13688 4740 13694 4752
rect 16393 4743 16451 4749
rect 16393 4740 16405 4743
rect 13688 4712 16405 4740
rect 13688 4700 13694 4712
rect 4801 4675 4859 4681
rect 4801 4641 4813 4675
rect 4847 4672 4859 4675
rect 7190 4672 7196 4684
rect 4847 4644 7196 4672
rect 4847 4641 4859 4644
rect 4801 4635 4859 4641
rect 7190 4632 7196 4644
rect 7248 4632 7254 4684
rect 7374 4672 7380 4684
rect 7300 4644 7380 4672
rect 1670 4564 1676 4616
rect 1728 4604 1734 4616
rect 2409 4607 2467 4613
rect 2409 4604 2421 4607
rect 1728 4576 2421 4604
rect 1728 4564 1734 4576
rect 2409 4573 2421 4576
rect 2455 4573 2467 4607
rect 2409 4567 2467 4573
rect 3329 4607 3387 4613
rect 3329 4573 3341 4607
rect 3375 4604 3387 4607
rect 3694 4604 3700 4616
rect 3375 4576 3700 4604
rect 3375 4573 3387 4576
rect 3329 4567 3387 4573
rect 3694 4564 3700 4576
rect 3752 4564 3758 4616
rect 4246 4564 4252 4616
rect 4304 4564 4310 4616
rect 4338 4564 4344 4616
rect 4396 4564 4402 4616
rect 4614 4564 4620 4616
rect 4672 4604 4678 4616
rect 5353 4607 5411 4613
rect 5353 4604 5365 4607
rect 4672 4576 5365 4604
rect 4672 4564 4678 4576
rect 5353 4573 5365 4576
rect 5399 4573 5411 4607
rect 5353 4567 5411 4573
rect 5534 4564 5540 4616
rect 5592 4564 5598 4616
rect 6914 4564 6920 4616
rect 6972 4564 6978 4616
rect 7300 4613 7328 4644
rect 7374 4632 7380 4644
rect 7432 4672 7438 4684
rect 8478 4672 8484 4684
rect 7432 4644 8484 4672
rect 7432 4632 7438 4644
rect 8478 4632 8484 4644
rect 8536 4632 8542 4684
rect 9306 4632 9312 4684
rect 9364 4672 9370 4684
rect 9585 4675 9643 4681
rect 9585 4672 9597 4675
rect 9364 4644 9597 4672
rect 9364 4632 9370 4644
rect 9585 4641 9597 4644
rect 9631 4641 9643 4675
rect 9585 4635 9643 4641
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 10134 4672 10140 4684
rect 10091 4644 10140 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 10134 4632 10140 4644
rect 10192 4632 10198 4684
rect 7009 4607 7067 4613
rect 7009 4573 7021 4607
rect 7055 4604 7067 4607
rect 7285 4607 7343 4613
rect 7055 4576 7144 4604
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 2130 4496 2136 4548
rect 2188 4496 2194 4548
rect 2774 4496 2780 4548
rect 2832 4536 2838 4548
rect 3053 4539 3111 4545
rect 3053 4536 3065 4539
rect 2832 4508 3065 4536
rect 2832 4496 2838 4508
rect 3053 4505 3065 4508
rect 3099 4505 3111 4539
rect 3053 4499 3111 4505
rect 3510 4496 3516 4548
rect 3568 4536 3574 4548
rect 4062 4536 4068 4548
rect 3568 4508 4068 4536
rect 3568 4496 3574 4508
rect 4062 4496 4068 4508
rect 4120 4496 4126 4548
rect 4430 4496 4436 4548
rect 4488 4496 4494 4548
rect 5258 4496 5264 4548
rect 5316 4496 5322 4548
rect 6270 4496 6276 4548
rect 6328 4496 6334 4548
rect 4522 4428 4528 4480
rect 4580 4468 4586 4480
rect 4982 4468 4988 4480
rect 4580 4440 4988 4468
rect 4580 4428 4586 4440
rect 4982 4428 4988 4440
rect 5040 4468 5046 4480
rect 7116 4468 7144 4576
rect 7285 4573 7297 4607
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 7466 4564 7472 4616
rect 7524 4564 7530 4616
rect 7929 4607 7987 4613
rect 7929 4573 7941 4607
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 7944 4536 7972 4567
rect 8110 4564 8116 4616
rect 8168 4564 8174 4616
rect 9677 4607 9735 4613
rect 9677 4573 9689 4607
rect 9723 4604 9735 4607
rect 10226 4604 10232 4616
rect 9723 4576 10232 4604
rect 9723 4573 9735 4576
rect 9677 4567 9735 4573
rect 10226 4564 10232 4576
rect 10284 4564 10290 4616
rect 12250 4564 12256 4616
rect 12308 4564 12314 4616
rect 12529 4607 12587 4613
rect 12529 4573 12541 4607
rect 12575 4604 12587 4607
rect 12710 4604 12716 4616
rect 12575 4576 12716 4604
rect 12575 4573 12587 4576
rect 12529 4567 12587 4573
rect 12710 4564 12716 4576
rect 12768 4564 12774 4616
rect 14550 4564 14556 4616
rect 14608 4564 14614 4616
rect 14734 4564 14740 4616
rect 14792 4604 14798 4616
rect 15764 4613 15792 4712
rect 16393 4709 16405 4712
rect 16439 4740 16451 4743
rect 18414 4740 18420 4752
rect 16439 4712 18420 4740
rect 16439 4709 16451 4712
rect 16393 4703 16451 4709
rect 18414 4700 18420 4712
rect 18472 4700 18478 4752
rect 16482 4672 16488 4684
rect 15856 4644 16488 4672
rect 14829 4607 14887 4613
rect 14829 4604 14841 4607
rect 14792 4576 14841 4604
rect 14792 4564 14798 4576
rect 14829 4573 14841 4576
rect 14875 4573 14887 4607
rect 14829 4567 14887 4573
rect 15749 4607 15807 4613
rect 15749 4573 15761 4607
rect 15795 4573 15807 4607
rect 15749 4567 15807 4573
rect 7944 4508 9168 4536
rect 5040 4440 7144 4468
rect 5040 4428 5046 4440
rect 7190 4428 7196 4480
rect 7248 4468 7254 4480
rect 7944 4468 7972 4508
rect 7248 4440 7972 4468
rect 8021 4471 8079 4477
rect 7248 4428 7254 4440
rect 8021 4437 8033 4471
rect 8067 4468 8079 4471
rect 9030 4468 9036 4480
rect 8067 4440 9036 4468
rect 8067 4437 8079 4440
rect 8021 4431 8079 4437
rect 9030 4428 9036 4440
rect 9088 4428 9094 4480
rect 9140 4468 9168 4508
rect 9950 4496 9956 4548
rect 10008 4496 10014 4548
rect 11330 4496 11336 4548
rect 11388 4536 11394 4548
rect 12437 4539 12495 4545
rect 12437 4536 12449 4539
rect 11388 4508 12449 4536
rect 11388 4496 11394 4508
rect 12437 4505 12449 4508
rect 12483 4536 12495 4539
rect 15856 4536 15884 4644
rect 16482 4632 16488 4644
rect 16540 4632 16546 4684
rect 16574 4632 16580 4684
rect 16632 4672 16638 4684
rect 18877 4675 18935 4681
rect 18877 4672 18889 4675
rect 16632 4644 18889 4672
rect 16632 4632 16638 4644
rect 18877 4641 18889 4644
rect 18923 4672 18935 4675
rect 18923 4644 19656 4672
rect 18923 4641 18935 4644
rect 18877 4635 18935 4641
rect 15930 4564 15936 4616
rect 15988 4564 15994 4616
rect 16022 4564 16028 4616
rect 16080 4604 16086 4616
rect 17497 4607 17555 4613
rect 17497 4604 17509 4607
rect 16080 4576 17509 4604
rect 16080 4564 16086 4576
rect 17497 4573 17509 4576
rect 17543 4573 17555 4607
rect 17497 4567 17555 4573
rect 17862 4564 17868 4616
rect 17920 4564 17926 4616
rect 19628 4613 19656 4644
rect 21450 4632 21456 4684
rect 21508 4672 21514 4684
rect 22649 4675 22707 4681
rect 22649 4672 22661 4675
rect 21508 4644 22661 4672
rect 21508 4632 21514 4644
rect 22649 4641 22661 4644
rect 22695 4641 22707 4675
rect 22649 4635 22707 4641
rect 19613 4607 19671 4613
rect 19613 4573 19625 4607
rect 19659 4573 19671 4607
rect 19613 4567 19671 4573
rect 22278 4564 22284 4616
rect 22336 4604 22342 4616
rect 22738 4604 22744 4616
rect 22336 4576 22744 4604
rect 22336 4564 22342 4576
rect 22738 4564 22744 4576
rect 22796 4564 22802 4616
rect 22922 4564 22928 4616
rect 22980 4564 22986 4616
rect 12483 4508 15884 4536
rect 12483 4505 12495 4508
rect 12437 4499 12495 4505
rect 16114 4496 16120 4548
rect 16172 4536 16178 4548
rect 17589 4539 17647 4545
rect 17589 4536 17601 4539
rect 16172 4508 17601 4536
rect 16172 4496 16178 4508
rect 17589 4505 17601 4508
rect 17635 4505 17647 4539
rect 17589 4499 17647 4505
rect 17681 4539 17739 4545
rect 17681 4505 17693 4539
rect 17727 4536 17739 4539
rect 19429 4539 19487 4545
rect 19429 4536 19441 4539
rect 17727 4508 19441 4536
rect 17727 4505 17739 4508
rect 17681 4499 17739 4505
rect 19429 4505 19441 4508
rect 19475 4505 19487 4539
rect 19429 4499 19487 4505
rect 10042 4468 10048 4480
rect 9140 4440 10048 4468
rect 10042 4428 10048 4440
rect 10100 4428 10106 4480
rect 10597 4471 10655 4477
rect 10597 4437 10609 4471
rect 10643 4468 10655 4471
rect 10778 4468 10784 4480
rect 10643 4440 10784 4468
rect 10643 4437 10655 4440
rect 10597 4431 10655 4437
rect 10778 4428 10784 4440
rect 10836 4428 10842 4480
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 12158 4468 12164 4480
rect 11112 4440 12164 4468
rect 11112 4428 11118 4440
rect 12158 4428 12164 4440
rect 12216 4428 12222 4480
rect 14550 4428 14556 4480
rect 14608 4468 14614 4480
rect 14645 4471 14703 4477
rect 14645 4468 14657 4471
rect 14608 4440 14657 4468
rect 14608 4428 14614 4440
rect 14645 4437 14657 4440
rect 14691 4437 14703 4471
rect 14645 4431 14703 4437
rect 16482 4428 16488 4480
rect 16540 4468 16546 4480
rect 17218 4468 17224 4480
rect 16540 4440 17224 4468
rect 16540 4428 16546 4440
rect 17218 4428 17224 4440
rect 17276 4468 17282 4480
rect 17696 4468 17724 4499
rect 17276 4440 17724 4468
rect 17276 4428 17282 4440
rect 1104 4378 23987 4400
rect 1104 4326 6630 4378
rect 6682 4326 6694 4378
rect 6746 4326 6758 4378
rect 6810 4326 6822 4378
rect 6874 4326 6886 4378
rect 6938 4326 12311 4378
rect 12363 4326 12375 4378
rect 12427 4326 12439 4378
rect 12491 4326 12503 4378
rect 12555 4326 12567 4378
rect 12619 4326 17992 4378
rect 18044 4326 18056 4378
rect 18108 4326 18120 4378
rect 18172 4326 18184 4378
rect 18236 4326 18248 4378
rect 18300 4326 23673 4378
rect 23725 4326 23737 4378
rect 23789 4326 23801 4378
rect 23853 4326 23865 4378
rect 23917 4326 23929 4378
rect 23981 4326 23987 4378
rect 1104 4304 23987 4326
rect 2222 4224 2228 4276
rect 2280 4264 2286 4276
rect 3050 4264 3056 4276
rect 2280 4236 3056 4264
rect 2280 4224 2286 4236
rect 3050 4224 3056 4236
rect 3108 4224 3114 4276
rect 4246 4224 4252 4276
rect 4304 4264 4310 4276
rect 5258 4264 5264 4276
rect 4304 4236 5264 4264
rect 4304 4224 4310 4236
rect 5258 4224 5264 4236
rect 5316 4264 5322 4276
rect 6086 4264 6092 4276
rect 5316 4236 6092 4264
rect 5316 4224 5322 4236
rect 6086 4224 6092 4236
rect 6144 4264 6150 4276
rect 6733 4267 6791 4273
rect 6733 4264 6745 4267
rect 6144 4236 6745 4264
rect 6144 4224 6150 4236
rect 6733 4233 6745 4236
rect 6779 4233 6791 4267
rect 6733 4227 6791 4233
rect 6825 4267 6883 4273
rect 6825 4233 6837 4267
rect 6871 4264 6883 4267
rect 7098 4264 7104 4276
rect 6871 4236 7104 4264
rect 6871 4233 6883 4236
rect 6825 4227 6883 4233
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 8110 4224 8116 4276
rect 8168 4264 8174 4276
rect 13446 4264 13452 4276
rect 8168 4236 13452 4264
rect 8168 4224 8174 4236
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 13538 4224 13544 4276
rect 13596 4264 13602 4276
rect 13633 4267 13691 4273
rect 13633 4264 13645 4267
rect 13596 4236 13645 4264
rect 13596 4224 13602 4236
rect 13633 4233 13645 4236
rect 13679 4233 13691 4267
rect 17954 4264 17960 4276
rect 13633 4227 13691 4233
rect 15212 4236 17960 4264
rect 3694 4156 3700 4208
rect 3752 4156 3758 4208
rect 4062 4156 4068 4208
rect 4120 4196 4126 4208
rect 5534 4196 5540 4208
rect 4120 4168 5540 4196
rect 4120 4156 4126 4168
rect 1946 4088 1952 4140
rect 2004 4088 2010 4140
rect 2038 4088 2044 4140
rect 2096 4088 2102 4140
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4128 2191 4131
rect 2498 4128 2504 4140
rect 2179 4100 2504 4128
rect 2179 4097 2191 4100
rect 2133 4091 2191 4097
rect 2498 4088 2504 4100
rect 2556 4128 2562 4140
rect 2777 4131 2835 4137
rect 2777 4128 2789 4131
rect 2556 4100 2789 4128
rect 2556 4088 2562 4100
rect 2777 4097 2789 4100
rect 2823 4097 2835 4131
rect 2777 4091 2835 4097
rect 1964 4060 1992 4088
rect 2590 4060 2596 4072
rect 1964 4032 2596 4060
rect 2590 4020 2596 4032
rect 2648 4060 2654 4072
rect 2685 4063 2743 4069
rect 2685 4060 2697 4063
rect 2648 4032 2697 4060
rect 2648 4020 2654 4032
rect 2685 4029 2697 4032
rect 2731 4029 2743 4063
rect 2792 4060 2820 4091
rect 3878 4088 3884 4140
rect 3936 4088 3942 4140
rect 4433 4131 4491 4137
rect 4433 4128 4445 4131
rect 3988 4100 4445 4128
rect 3694 4060 3700 4072
rect 2792 4032 3700 4060
rect 2685 4023 2743 4029
rect 3694 4020 3700 4032
rect 3752 4060 3758 4072
rect 3988 4060 4016 4100
rect 4433 4097 4445 4100
rect 4479 4128 4491 4131
rect 4522 4128 4528 4140
rect 4479 4100 4528 4128
rect 4479 4097 4491 4100
rect 4433 4091 4491 4097
rect 4522 4088 4528 4100
rect 4580 4088 4586 4140
rect 4632 4137 4660 4168
rect 5534 4156 5540 4168
rect 5592 4156 5598 4208
rect 6641 4199 6699 4205
rect 6641 4165 6653 4199
rect 6687 4196 6699 4199
rect 7006 4196 7012 4208
rect 6687 4168 7012 4196
rect 6687 4165 6699 4168
rect 6641 4159 6699 4165
rect 7006 4156 7012 4168
rect 7064 4196 7070 4208
rect 7064 4168 8340 4196
rect 7064 4156 7070 4168
rect 8312 4140 8340 4168
rect 14734 4156 14740 4208
rect 14792 4196 14798 4208
rect 15212 4196 15240 4236
rect 17954 4224 17960 4236
rect 18012 4224 18018 4276
rect 22646 4224 22652 4276
rect 22704 4224 22710 4276
rect 14792 4168 15240 4196
rect 14792 4156 14798 4168
rect 15378 4156 15384 4208
rect 15436 4196 15442 4208
rect 15436 4168 15976 4196
rect 15436 4156 15442 4168
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4097 4675 4131
rect 5258 4128 5264 4140
rect 4617 4091 4675 4097
rect 4724 4100 5264 4128
rect 3752 4032 4016 4060
rect 3752 4020 3758 4032
rect 4154 4020 4160 4072
rect 4212 4060 4218 4072
rect 4724 4060 4752 4100
rect 5258 4088 5264 4100
rect 5316 4128 5322 4140
rect 5445 4131 5503 4137
rect 5445 4128 5457 4131
rect 5316 4100 5457 4128
rect 5316 4088 5322 4100
rect 5445 4097 5457 4100
rect 5491 4097 5503 4131
rect 5445 4091 5503 4097
rect 5629 4131 5687 4137
rect 5629 4097 5641 4131
rect 5675 4097 5687 4131
rect 5629 4091 5687 4097
rect 5997 4131 6055 4137
rect 5997 4097 6009 4131
rect 6043 4128 6055 4131
rect 6454 4128 6460 4140
rect 6043 4100 6460 4128
rect 6043 4097 6055 4100
rect 5997 4091 6055 4097
rect 4212 4032 4752 4060
rect 4212 4020 4218 4032
rect 4890 4020 4896 4072
rect 4948 4020 4954 4072
rect 2038 3952 2044 4004
rect 2096 3992 2102 4004
rect 2866 3992 2872 4004
rect 2096 3964 2872 3992
rect 2096 3952 2102 3964
rect 2866 3952 2872 3964
rect 2924 3952 2930 4004
rect 3602 3952 3608 4004
rect 3660 3992 3666 4004
rect 3878 3992 3884 4004
rect 3660 3964 3884 3992
rect 3660 3952 3666 3964
rect 3878 3952 3884 3964
rect 3936 3992 3942 4004
rect 3936 3964 4384 3992
rect 3936 3952 3942 3964
rect 1765 3927 1823 3933
rect 1765 3893 1777 3927
rect 1811 3924 1823 3927
rect 2314 3924 2320 3936
rect 1811 3896 2320 3924
rect 1811 3893 1823 3896
rect 1765 3887 1823 3893
rect 2314 3884 2320 3896
rect 2372 3884 2378 3936
rect 2961 3927 3019 3933
rect 2961 3893 2973 3927
rect 3007 3924 3019 3927
rect 4246 3924 4252 3936
rect 3007 3896 4252 3924
rect 3007 3893 3019 3896
rect 2961 3887 3019 3893
rect 4246 3884 4252 3896
rect 4304 3884 4310 3936
rect 4356 3924 4384 3964
rect 4614 3952 4620 4004
rect 4672 3992 4678 4004
rect 5644 3992 5672 4091
rect 6454 4088 6460 4100
rect 6512 4128 6518 4140
rect 7377 4131 7435 4137
rect 7377 4128 7389 4131
rect 6512 4100 7389 4128
rect 6512 4088 6518 4100
rect 7377 4097 7389 4100
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 7834 4088 7840 4140
rect 7892 4128 7898 4140
rect 8113 4131 8171 4137
rect 8113 4128 8125 4131
rect 7892 4100 8125 4128
rect 7892 4088 7898 4100
rect 8113 4097 8125 4100
rect 8159 4097 8171 4131
rect 8113 4091 8171 4097
rect 8294 4088 8300 4140
rect 8352 4088 8358 4140
rect 8754 4088 8760 4140
rect 8812 4088 8818 4140
rect 9033 4131 9091 4137
rect 9033 4097 9045 4131
rect 9079 4097 9091 4131
rect 9033 4091 9091 4097
rect 7190 4020 7196 4072
rect 7248 4020 7254 4072
rect 7926 4020 7932 4072
rect 7984 4060 7990 4072
rect 9048 4060 9076 4091
rect 9214 4088 9220 4140
rect 9272 4088 9278 4140
rect 14277 4131 14335 4137
rect 14277 4097 14289 4131
rect 14323 4128 14335 4131
rect 14550 4128 14556 4140
rect 14323 4100 14556 4128
rect 14323 4097 14335 4100
rect 14277 4091 14335 4097
rect 14550 4088 14556 4100
rect 14608 4128 14614 4140
rect 15197 4131 15255 4137
rect 15197 4128 15209 4131
rect 14608 4100 15209 4128
rect 14608 4088 14614 4100
rect 15197 4097 15209 4100
rect 15243 4128 15255 4131
rect 15838 4128 15844 4140
rect 15243 4100 15844 4128
rect 15243 4097 15255 4100
rect 15197 4091 15255 4097
rect 15838 4088 15844 4100
rect 15896 4088 15902 4140
rect 15948 4137 15976 4168
rect 18690 4156 18696 4208
rect 18748 4196 18754 4208
rect 22922 4196 22928 4208
rect 18748 4168 19288 4196
rect 18748 4156 18754 4168
rect 15933 4131 15991 4137
rect 15933 4097 15945 4131
rect 15979 4097 15991 4131
rect 15933 4091 15991 4097
rect 16025 4131 16083 4137
rect 16025 4097 16037 4131
rect 16071 4097 16083 4131
rect 16025 4091 16083 4097
rect 16114 4091 16120 4143
rect 16172 4091 16178 4143
rect 19260 4140 19288 4168
rect 22572 4168 22928 4196
rect 7984 4032 9076 4060
rect 7984 4020 7990 4032
rect 9122 4020 9128 4072
rect 9180 4060 9186 4072
rect 11606 4060 11612 4072
rect 9180 4032 11612 4060
rect 9180 4020 9186 4032
rect 11606 4020 11612 4032
rect 11664 4020 11670 4072
rect 7466 3992 7472 4004
rect 4672 3964 7472 3992
rect 4672 3952 4678 3964
rect 7466 3952 7472 3964
rect 7524 3952 7530 4004
rect 8478 3952 8484 4004
rect 8536 3992 8542 4004
rect 12158 3992 12164 4004
rect 8536 3964 12164 3992
rect 8536 3952 8542 3964
rect 12158 3952 12164 3964
rect 12216 3952 12222 4004
rect 13722 3952 13728 4004
rect 13780 3992 13786 4004
rect 16040 3992 16068 4091
rect 16298 4088 16304 4140
rect 16356 4128 16362 4140
rect 16853 4131 16911 4137
rect 16853 4128 16865 4131
rect 16356 4100 16865 4128
rect 16356 4088 16362 4100
rect 16853 4097 16865 4100
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 17310 4088 17316 4140
rect 17368 4128 17374 4140
rect 18509 4131 18567 4137
rect 18509 4128 18521 4131
rect 17368 4100 18521 4128
rect 17368 4088 17374 4100
rect 18509 4097 18521 4100
rect 18555 4097 18567 4131
rect 18969 4131 19027 4137
rect 18969 4128 18981 4131
rect 18509 4091 18567 4097
rect 18600 4100 18981 4128
rect 17954 4020 17960 4072
rect 18012 4060 18018 4072
rect 18600 4060 18628 4100
rect 18969 4097 18981 4100
rect 19015 4097 19027 4131
rect 18969 4091 19027 4097
rect 19153 4131 19211 4137
rect 19153 4097 19165 4131
rect 19199 4097 19211 4131
rect 19153 4091 19211 4097
rect 18012 4032 18628 4060
rect 18012 4020 18018 4032
rect 18874 4020 18880 4072
rect 18932 4060 18938 4072
rect 19168 4060 19196 4091
rect 19242 4088 19248 4140
rect 19300 4128 19306 4140
rect 19337 4131 19395 4137
rect 19337 4128 19349 4131
rect 19300 4100 19349 4128
rect 19300 4088 19306 4100
rect 19337 4097 19349 4100
rect 19383 4097 19395 4131
rect 19337 4091 19395 4097
rect 19518 4088 19524 4140
rect 19576 4088 19582 4140
rect 19794 4088 19800 4140
rect 19852 4088 19858 4140
rect 22572 4137 22600 4168
rect 22922 4156 22928 4168
rect 22980 4156 22986 4208
rect 22557 4131 22615 4137
rect 22557 4097 22569 4131
rect 22603 4097 22615 4131
rect 22557 4091 22615 4097
rect 22738 4088 22744 4140
rect 22796 4088 22802 4140
rect 18932 4032 19196 4060
rect 18932 4020 18938 4032
rect 13780 3964 16068 3992
rect 13780 3952 13786 3964
rect 7098 3924 7104 3936
rect 4356 3896 7104 3924
rect 7098 3884 7104 3896
rect 7156 3884 7162 3936
rect 8113 3927 8171 3933
rect 8113 3893 8125 3927
rect 8159 3924 8171 3927
rect 8386 3924 8392 3936
rect 8159 3896 8392 3924
rect 8159 3893 8171 3896
rect 8113 3887 8171 3893
rect 8386 3884 8392 3896
rect 8444 3884 8450 3936
rect 8846 3884 8852 3936
rect 8904 3884 8910 3936
rect 9677 3927 9735 3933
rect 9677 3893 9689 3927
rect 9723 3924 9735 3927
rect 9858 3924 9864 3936
rect 9723 3896 9864 3924
rect 9723 3893 9735 3896
rect 9677 3887 9735 3893
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 10318 3884 10324 3936
rect 10376 3884 10382 3936
rect 10410 3884 10416 3936
rect 10468 3924 10474 3936
rect 10965 3927 11023 3933
rect 10965 3924 10977 3927
rect 10468 3896 10977 3924
rect 10468 3884 10474 3896
rect 10965 3893 10977 3896
rect 11011 3893 11023 3927
rect 10965 3887 11023 3893
rect 11698 3884 11704 3936
rect 11756 3884 11762 3936
rect 11790 3884 11796 3936
rect 11848 3924 11854 3936
rect 12253 3927 12311 3933
rect 12253 3924 12265 3927
rect 11848 3896 12265 3924
rect 11848 3884 11854 3896
rect 12253 3893 12265 3896
rect 12299 3893 12311 3927
rect 12253 3887 12311 3893
rect 15654 3884 15660 3936
rect 15712 3884 15718 3936
rect 16040 3924 16068 3964
rect 17310 3924 17316 3936
rect 16040 3896 17316 3924
rect 17310 3884 17316 3896
rect 17368 3884 17374 3936
rect 1104 3834 23828 3856
rect 1104 3782 3790 3834
rect 3842 3782 3854 3834
rect 3906 3782 3918 3834
rect 3970 3782 3982 3834
rect 4034 3782 4046 3834
rect 4098 3782 9471 3834
rect 9523 3782 9535 3834
rect 9587 3782 9599 3834
rect 9651 3782 9663 3834
rect 9715 3782 9727 3834
rect 9779 3782 15152 3834
rect 15204 3782 15216 3834
rect 15268 3782 15280 3834
rect 15332 3782 15344 3834
rect 15396 3782 15408 3834
rect 15460 3782 20833 3834
rect 20885 3782 20897 3834
rect 20949 3782 20961 3834
rect 21013 3782 21025 3834
rect 21077 3782 21089 3834
rect 21141 3782 23828 3834
rect 1104 3760 23828 3782
rect 2498 3680 2504 3732
rect 2556 3680 2562 3732
rect 4430 3720 4436 3732
rect 3160 3692 4436 3720
rect 2866 3652 2872 3664
rect 2332 3624 2872 3652
rect 2332 3525 2360 3624
rect 2866 3612 2872 3624
rect 2924 3612 2930 3664
rect 2958 3612 2964 3664
rect 3016 3652 3022 3664
rect 3053 3655 3111 3661
rect 3053 3652 3065 3655
rect 3016 3624 3065 3652
rect 3016 3612 3022 3624
rect 3053 3621 3065 3624
rect 3099 3621 3111 3655
rect 3053 3615 3111 3621
rect 2590 3544 2596 3596
rect 2648 3544 2654 3596
rect 3160 3584 3188 3692
rect 4430 3680 4436 3692
rect 4488 3720 4494 3732
rect 8570 3720 8576 3732
rect 4488 3692 8576 3720
rect 4488 3680 4494 3692
rect 8570 3680 8576 3692
rect 8628 3720 8634 3732
rect 10778 3720 10784 3732
rect 8628 3692 10784 3720
rect 8628 3680 8634 3692
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 12802 3680 12808 3732
rect 12860 3720 12866 3732
rect 13081 3723 13139 3729
rect 13081 3720 13093 3723
rect 12860 3692 13093 3720
rect 12860 3680 12866 3692
rect 13081 3689 13093 3692
rect 13127 3689 13139 3723
rect 13081 3683 13139 3689
rect 14826 3680 14832 3732
rect 14884 3720 14890 3732
rect 17586 3720 17592 3732
rect 14884 3692 17592 3720
rect 14884 3680 14890 3692
rect 17586 3680 17592 3692
rect 17644 3680 17650 3732
rect 17770 3680 17776 3732
rect 17828 3720 17834 3732
rect 17954 3720 17960 3732
rect 17828 3692 17960 3720
rect 17828 3680 17834 3692
rect 17954 3680 17960 3692
rect 18012 3680 18018 3732
rect 6089 3655 6147 3661
rect 6089 3621 6101 3655
rect 6135 3652 6147 3655
rect 8202 3652 8208 3664
rect 6135 3624 8208 3652
rect 6135 3621 6147 3624
rect 6089 3615 6147 3621
rect 8202 3612 8208 3624
rect 8260 3612 8266 3664
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 10873 3655 10931 3661
rect 10873 3652 10885 3655
rect 10008 3624 10885 3652
rect 10008 3612 10014 3624
rect 10873 3621 10885 3624
rect 10919 3621 10931 3655
rect 10873 3615 10931 3621
rect 11882 3612 11888 3664
rect 11940 3652 11946 3664
rect 17862 3652 17868 3664
rect 11940 3624 17868 3652
rect 11940 3612 11946 3624
rect 2700 3556 3188 3584
rect 2317 3519 2375 3525
rect 2317 3485 2329 3519
rect 2363 3485 2375 3519
rect 2317 3479 2375 3485
rect 2498 3476 2504 3528
rect 2556 3516 2562 3528
rect 2700 3516 2728 3556
rect 3510 3544 3516 3596
rect 3568 3544 3574 3596
rect 4706 3544 4712 3596
rect 4764 3584 4770 3596
rect 5718 3584 5724 3596
rect 4764 3556 5724 3584
rect 4764 3544 4770 3556
rect 2556 3488 2728 3516
rect 2556 3476 2562 3488
rect 3050 3476 3056 3528
rect 3108 3516 3114 3528
rect 3328 3519 3386 3525
rect 3328 3516 3340 3519
rect 3108 3488 3340 3516
rect 3108 3476 3114 3488
rect 3328 3485 3340 3488
rect 3374 3485 3386 3519
rect 3328 3479 3386 3485
rect 3414 3519 3472 3525
rect 3414 3485 3426 3519
rect 3460 3516 3472 3519
rect 3528 3516 3556 3544
rect 3460 3488 3556 3516
rect 4433 3519 4491 3525
rect 3460 3485 3472 3488
rect 3414 3479 3472 3485
rect 4433 3485 4445 3519
rect 4479 3516 4491 3519
rect 4798 3516 4804 3528
rect 4479 3488 4804 3516
rect 4479 3485 4491 3488
rect 4433 3479 4491 3485
rect 1673 3451 1731 3457
rect 1673 3417 1685 3451
rect 1719 3448 1731 3451
rect 3234 3448 3240 3460
rect 1719 3420 3240 3448
rect 1719 3417 1731 3420
rect 1673 3411 1731 3417
rect 3234 3408 3240 3420
rect 3292 3408 3298 3460
rect 2133 3383 2191 3389
rect 2133 3349 2145 3383
rect 2179 3380 2191 3383
rect 2222 3380 2228 3392
rect 2179 3352 2228 3380
rect 2179 3349 2191 3352
rect 2133 3343 2191 3349
rect 2222 3340 2228 3352
rect 2280 3340 2286 3392
rect 3344 3380 3372 3479
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 5184 3525 5212 3556
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 5810 3544 5816 3596
rect 5868 3584 5874 3596
rect 6733 3587 6791 3593
rect 6733 3584 6745 3587
rect 5868 3556 6745 3584
rect 5868 3544 5874 3556
rect 6733 3553 6745 3556
rect 6779 3553 6791 3587
rect 6733 3547 6791 3553
rect 7929 3587 7987 3593
rect 7929 3553 7941 3587
rect 7975 3584 7987 3587
rect 10413 3587 10471 3593
rect 10413 3584 10425 3587
rect 7975 3556 10425 3584
rect 7975 3553 7987 3556
rect 7929 3547 7987 3553
rect 10413 3553 10425 3556
rect 10459 3584 10471 3587
rect 10502 3584 10508 3596
rect 10459 3556 10508 3584
rect 10459 3553 10471 3556
rect 10413 3547 10471 3553
rect 10502 3544 10508 3556
rect 10560 3544 10566 3596
rect 11149 3587 11207 3593
rect 11149 3553 11161 3587
rect 11195 3584 11207 3587
rect 11900 3584 11928 3612
rect 11195 3556 11928 3584
rect 11195 3553 11207 3556
rect 11149 3547 11207 3553
rect 12710 3544 12716 3596
rect 12768 3584 12774 3596
rect 12805 3587 12863 3593
rect 12805 3584 12817 3587
rect 12768 3556 12817 3584
rect 12768 3544 12774 3556
rect 12805 3553 12817 3556
rect 12851 3553 12863 3587
rect 12805 3547 12863 3553
rect 4893 3519 4951 3525
rect 4893 3485 4905 3519
rect 4939 3516 4951 3519
rect 5169 3519 5227 3525
rect 4939 3488 5028 3516
rect 4939 3485 4951 3488
rect 4893 3479 4951 3485
rect 4062 3408 4068 3460
rect 4120 3448 4126 3460
rect 4157 3451 4215 3457
rect 4157 3448 4169 3451
rect 4120 3420 4169 3448
rect 4120 3408 4126 3420
rect 4157 3417 4169 3420
rect 4203 3417 4215 3451
rect 4157 3411 4215 3417
rect 4246 3408 4252 3460
rect 4304 3448 4310 3460
rect 5000 3448 5028 3488
rect 5169 3485 5181 3519
rect 5215 3485 5227 3519
rect 5169 3479 5227 3485
rect 5258 3476 5264 3528
rect 5316 3476 5322 3528
rect 5629 3519 5687 3525
rect 5629 3485 5641 3519
rect 5675 3516 5687 3519
rect 6270 3516 6276 3528
rect 5675 3488 6276 3516
rect 5675 3485 5687 3488
rect 5629 3479 5687 3485
rect 6270 3476 6276 3488
rect 6328 3476 6334 3528
rect 6546 3476 6552 3528
rect 6604 3476 6610 3528
rect 7834 3476 7840 3528
rect 7892 3476 7898 3528
rect 8021 3519 8079 3525
rect 8021 3485 8033 3519
rect 8067 3516 8079 3519
rect 8110 3516 8116 3528
rect 8067 3488 8116 3516
rect 8067 3485 8079 3488
rect 8021 3479 8079 3485
rect 8110 3476 8116 3488
rect 8168 3476 8174 3528
rect 9214 3476 9220 3528
rect 9272 3516 9278 3528
rect 9309 3519 9367 3525
rect 9309 3516 9321 3519
rect 9272 3488 9321 3516
rect 9272 3476 9278 3488
rect 9309 3485 9321 3488
rect 9355 3485 9367 3519
rect 9309 3479 9367 3485
rect 9950 3476 9956 3528
rect 10008 3476 10014 3528
rect 10226 3476 10232 3528
rect 10284 3476 10290 3528
rect 11054 3476 11060 3528
rect 11112 3476 11118 3528
rect 11517 3519 11575 3525
rect 11517 3485 11529 3519
rect 11563 3516 11575 3519
rect 11563 3488 12434 3516
rect 11563 3485 11575 3488
rect 11517 3479 11575 3485
rect 4304 3420 5028 3448
rect 4304 3408 4310 3420
rect 4614 3380 4620 3392
rect 3344 3352 4620 3380
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 5000 3380 5028 3420
rect 5074 3408 5080 3460
rect 5132 3448 5138 3460
rect 5132 3420 5764 3448
rect 5132 3408 5138 3420
rect 5626 3380 5632 3392
rect 5000 3352 5632 3380
rect 5626 3340 5632 3352
rect 5684 3340 5690 3392
rect 5736 3380 5764 3420
rect 6178 3408 6184 3460
rect 6236 3448 6242 3460
rect 7852 3448 7880 3476
rect 6236 3420 7880 3448
rect 6236 3408 6242 3420
rect 8294 3408 8300 3460
rect 8352 3448 8358 3460
rect 11146 3448 11152 3460
rect 8352 3420 11152 3448
rect 8352 3408 8358 3420
rect 11146 3408 11152 3420
rect 11204 3408 11210 3460
rect 11422 3408 11428 3460
rect 11480 3408 11486 3460
rect 12406 3448 12434 3488
rect 12894 3476 12900 3528
rect 12952 3476 12958 3528
rect 13556 3525 13584 3624
rect 17862 3612 17868 3624
rect 17920 3612 17926 3664
rect 14366 3544 14372 3596
rect 14424 3584 14430 3596
rect 14921 3587 14979 3593
rect 14921 3584 14933 3587
rect 14424 3556 14933 3584
rect 14424 3544 14430 3556
rect 14921 3553 14933 3556
rect 14967 3553 14979 3587
rect 14921 3547 14979 3553
rect 20070 3544 20076 3596
rect 20128 3544 20134 3596
rect 22373 3587 22431 3593
rect 22373 3553 22385 3587
rect 22419 3584 22431 3587
rect 23382 3584 23388 3596
rect 22419 3556 23388 3584
rect 22419 3553 22431 3556
rect 22373 3547 22431 3553
rect 23382 3544 23388 3556
rect 23440 3544 23446 3596
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3485 13599 3519
rect 13541 3479 13599 3485
rect 13725 3519 13783 3525
rect 13725 3485 13737 3519
rect 13771 3485 13783 3519
rect 13725 3479 13783 3485
rect 13740 3448 13768 3479
rect 14274 3476 14280 3528
rect 14332 3476 14338 3528
rect 14461 3519 14519 3525
rect 14461 3485 14473 3519
rect 14507 3485 14519 3519
rect 14461 3479 14519 3485
rect 14369 3451 14427 3457
rect 14369 3448 14381 3451
rect 12406 3420 14381 3448
rect 14369 3417 14381 3420
rect 14415 3417 14427 3451
rect 14476 3448 14504 3479
rect 15010 3476 15016 3528
rect 15068 3516 15074 3528
rect 15565 3519 15623 3525
rect 15565 3516 15577 3519
rect 15068 3488 15577 3516
rect 15068 3476 15074 3488
rect 15565 3485 15577 3488
rect 15611 3485 15623 3519
rect 15565 3479 15623 3485
rect 15654 3476 15660 3528
rect 15712 3516 15718 3528
rect 16209 3519 16267 3525
rect 16209 3516 16221 3519
rect 15712 3488 16221 3516
rect 15712 3476 15718 3488
rect 16209 3485 16221 3488
rect 16255 3485 16267 3519
rect 16209 3479 16267 3485
rect 18414 3476 18420 3528
rect 18472 3516 18478 3528
rect 18877 3519 18935 3525
rect 18877 3516 18889 3519
rect 18472 3488 18889 3516
rect 18472 3476 18478 3488
rect 18877 3485 18889 3488
rect 18923 3516 18935 3519
rect 19797 3519 19855 3525
rect 19797 3516 19809 3519
rect 18923 3488 19809 3516
rect 18923 3485 18935 3488
rect 18877 3479 18935 3485
rect 19797 3485 19809 3488
rect 19843 3485 19855 3519
rect 19797 3479 19855 3485
rect 22738 3476 22744 3528
rect 22796 3516 22802 3528
rect 22833 3519 22891 3525
rect 22833 3516 22845 3519
rect 22796 3488 22845 3516
rect 22796 3476 22802 3488
rect 22833 3485 22845 3488
rect 22879 3485 22891 3519
rect 22833 3479 22891 3485
rect 15194 3448 15200 3460
rect 14476 3420 15200 3448
rect 14369 3411 14427 3417
rect 15194 3408 15200 3420
rect 15252 3448 15258 3460
rect 16022 3448 16028 3460
rect 15252 3420 16028 3448
rect 15252 3408 15258 3420
rect 16022 3408 16028 3420
rect 16080 3408 16086 3460
rect 8110 3380 8116 3392
rect 5736 3352 8116 3380
rect 8110 3340 8116 3352
rect 8168 3340 8174 3392
rect 8938 3340 8944 3392
rect 8996 3380 9002 3392
rect 10045 3383 10103 3389
rect 10045 3380 10057 3383
rect 8996 3352 10057 3380
rect 8996 3340 9002 3352
rect 10045 3349 10057 3352
rect 10091 3380 10103 3383
rect 10134 3380 10140 3392
rect 10091 3352 10140 3380
rect 10091 3349 10103 3352
rect 10045 3343 10103 3349
rect 10134 3340 10140 3352
rect 10192 3380 10198 3392
rect 11238 3380 11244 3392
rect 10192 3352 11244 3380
rect 10192 3340 10198 3352
rect 11238 3340 11244 3352
rect 11296 3340 11302 3392
rect 11330 3340 11336 3392
rect 11388 3340 11394 3392
rect 11514 3340 11520 3392
rect 11572 3380 11578 3392
rect 12437 3383 12495 3389
rect 12437 3380 12449 3383
rect 11572 3352 12449 3380
rect 11572 3340 11578 3352
rect 12437 3349 12449 3352
rect 12483 3349 12495 3383
rect 12437 3343 12495 3349
rect 13262 3340 13268 3392
rect 13320 3380 13326 3392
rect 13633 3383 13691 3389
rect 13633 3380 13645 3383
rect 13320 3352 13645 3380
rect 13320 3340 13326 3352
rect 13633 3349 13645 3352
rect 13679 3380 13691 3383
rect 15470 3380 15476 3392
rect 13679 3352 15476 3380
rect 13679 3349 13691 3352
rect 13633 3343 13691 3349
rect 15470 3340 15476 3352
rect 15528 3340 15534 3392
rect 15562 3340 15568 3392
rect 15620 3380 15626 3392
rect 15838 3380 15844 3392
rect 15620 3352 15844 3380
rect 15620 3340 15626 3352
rect 15838 3340 15844 3352
rect 15896 3340 15902 3392
rect 16758 3340 16764 3392
rect 16816 3380 16822 3392
rect 16853 3383 16911 3389
rect 16853 3380 16865 3383
rect 16816 3352 16865 3380
rect 16816 3340 16822 3352
rect 16853 3349 16865 3352
rect 16899 3349 16911 3383
rect 16853 3343 16911 3349
rect 17402 3340 17408 3392
rect 17460 3340 17466 3392
rect 18874 3340 18880 3392
rect 18932 3380 18938 3392
rect 19503 3383 19561 3389
rect 19503 3380 19515 3383
rect 18932 3352 19515 3380
rect 18932 3340 18938 3352
rect 19503 3349 19515 3352
rect 19549 3349 19561 3383
rect 19503 3343 19561 3349
rect 19978 3340 19984 3392
rect 20036 3340 20042 3392
rect 20622 3340 20628 3392
rect 20680 3340 20686 3392
rect 1104 3290 23987 3312
rect 1104 3238 6630 3290
rect 6682 3238 6694 3290
rect 6746 3238 6758 3290
rect 6810 3238 6822 3290
rect 6874 3238 6886 3290
rect 6938 3238 12311 3290
rect 12363 3238 12375 3290
rect 12427 3238 12439 3290
rect 12491 3238 12503 3290
rect 12555 3238 12567 3290
rect 12619 3238 17992 3290
rect 18044 3238 18056 3290
rect 18108 3238 18120 3290
rect 18172 3238 18184 3290
rect 18236 3238 18248 3290
rect 18300 3238 23673 3290
rect 23725 3238 23737 3290
rect 23789 3238 23801 3290
rect 23853 3238 23865 3290
rect 23917 3238 23929 3290
rect 23981 3238 23987 3290
rect 1104 3216 23987 3238
rect 2958 3176 2964 3188
rect 2516 3148 2964 3176
rect 2222 3000 2228 3052
rect 2280 3000 2286 3052
rect 2314 3000 2320 3052
rect 2372 3040 2378 3052
rect 2516 3049 2544 3148
rect 2958 3136 2964 3148
rect 3016 3136 3022 3188
rect 5442 3136 5448 3188
rect 5500 3136 5506 3188
rect 5718 3136 5724 3188
rect 5776 3176 5782 3188
rect 6546 3176 6552 3188
rect 5776 3148 6552 3176
rect 5776 3136 5782 3148
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 9122 3176 9128 3188
rect 8168 3148 9128 3176
rect 8168 3136 8174 3148
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 9585 3179 9643 3185
rect 9585 3145 9597 3179
rect 9631 3176 9643 3179
rect 11514 3176 11520 3188
rect 9631 3148 11520 3176
rect 9631 3145 9643 3148
rect 9585 3139 9643 3145
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 11882 3136 11888 3188
rect 11940 3136 11946 3188
rect 12710 3136 12716 3188
rect 12768 3176 12774 3188
rect 13173 3179 13231 3185
rect 13173 3176 13185 3179
rect 12768 3148 13185 3176
rect 12768 3136 12774 3148
rect 13173 3145 13185 3148
rect 13219 3145 13231 3179
rect 13173 3139 13231 3145
rect 16114 3136 16120 3188
rect 16172 3176 16178 3188
rect 16853 3179 16911 3185
rect 16853 3176 16865 3179
rect 16172 3148 16865 3176
rect 16172 3136 16178 3148
rect 16853 3145 16865 3148
rect 16899 3145 16911 3179
rect 16853 3139 16911 3145
rect 17402 3136 17408 3188
rect 17460 3176 17466 3188
rect 17460 3148 19656 3176
rect 17460 3136 17466 3148
rect 2590 3068 2596 3120
rect 2648 3068 2654 3120
rect 2682 3068 2688 3120
rect 2740 3108 2746 3120
rect 2740 3080 2820 3108
rect 2740 3068 2746 3080
rect 2408 3043 2466 3049
rect 2408 3040 2420 3043
rect 2372 3012 2420 3040
rect 2372 3000 2378 3012
rect 2408 3009 2420 3012
rect 2454 3009 2466 3043
rect 2408 3003 2466 3009
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3009 2559 3043
rect 2608 3040 2636 3068
rect 2792 3049 2820 3080
rect 3694 3068 3700 3120
rect 3752 3108 3758 3120
rect 4433 3111 4491 3117
rect 3752 3080 4016 3108
rect 3752 3068 3758 3080
rect 3988 3049 4016 3080
rect 4433 3077 4445 3111
rect 4479 3108 4491 3111
rect 5902 3108 5908 3120
rect 4479 3080 5908 3108
rect 4479 3077 4491 3080
rect 4433 3071 4491 3077
rect 2777 3043 2835 3049
rect 2608 3012 2728 3040
rect 2501 3003 2559 3009
rect 2590 2932 2596 2984
rect 2648 2932 2654 2984
rect 2700 2972 2728 3012
rect 2777 3009 2789 3043
rect 2823 3009 2835 3043
rect 2777 3003 2835 3009
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3009 3847 3043
rect 3789 3003 3847 3009
rect 3973 3043 4031 3049
rect 3973 3009 3985 3043
rect 4019 3009 4031 3043
rect 3973 3003 4031 3009
rect 4065 3043 4123 3049
rect 4065 3009 4077 3043
rect 4111 3040 4123 3043
rect 4154 3040 4160 3052
rect 4111 3012 4160 3040
rect 4111 3009 4123 3012
rect 4065 3003 4123 3009
rect 3804 2972 3832 3003
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3040 4307 3043
rect 4614 3040 4620 3052
rect 4295 3012 4620 3040
rect 4295 3009 4307 3012
rect 4249 3003 4307 3009
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 5092 3049 5120 3080
rect 5902 3068 5908 3080
rect 5960 3068 5966 3120
rect 6270 3068 6276 3120
rect 6328 3108 6334 3120
rect 6328 3080 9352 3108
rect 6328 3068 6334 3080
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3009 5135 3043
rect 5077 3003 5135 3009
rect 5442 3000 5448 3052
rect 5500 3000 5506 3052
rect 5629 3043 5687 3049
rect 5629 3009 5641 3043
rect 5675 3040 5687 3043
rect 5718 3040 5724 3052
rect 5675 3012 5724 3040
rect 5675 3009 5687 3012
rect 5629 3003 5687 3009
rect 5718 3000 5724 3012
rect 5776 3040 5782 3052
rect 6178 3040 6184 3052
rect 5776 3012 6184 3040
rect 5776 3000 5782 3012
rect 6178 3000 6184 3012
rect 6236 3000 6242 3052
rect 6546 3000 6552 3052
rect 6604 3000 6610 3052
rect 7377 3043 7435 3049
rect 7377 3040 7389 3043
rect 6932 3012 7389 3040
rect 4706 2972 4712 2984
rect 2700 2944 4712 2972
rect 4706 2932 4712 2944
rect 4764 2932 4770 2984
rect 5169 2975 5227 2981
rect 5169 2941 5181 2975
rect 5215 2972 5227 2975
rect 5460 2972 5488 3000
rect 5215 2944 5488 2972
rect 5215 2941 5227 2944
rect 5169 2935 5227 2941
rect 1854 2864 1860 2916
rect 1912 2904 1918 2916
rect 2682 2904 2688 2916
rect 1912 2876 2688 2904
rect 1912 2864 1918 2876
rect 2682 2864 2688 2876
rect 2740 2864 2746 2916
rect 2958 2864 2964 2916
rect 3016 2864 3022 2916
rect 4157 2907 4215 2913
rect 4157 2873 4169 2907
rect 4203 2904 4215 2907
rect 4522 2904 4528 2916
rect 4203 2876 4528 2904
rect 4203 2873 4215 2876
rect 4157 2867 4215 2873
rect 4522 2864 4528 2876
rect 4580 2864 4586 2916
rect 6546 2904 6552 2916
rect 4632 2876 6552 2904
rect 1765 2839 1823 2845
rect 1765 2805 1777 2839
rect 1811 2836 1823 2839
rect 4632 2836 4660 2876
rect 6546 2864 6552 2876
rect 6604 2864 6610 2916
rect 1811 2808 4660 2836
rect 1811 2805 1823 2808
rect 1765 2799 1823 2805
rect 4890 2796 4896 2848
rect 4948 2836 4954 2848
rect 6932 2836 6960 3012
rect 7377 3009 7389 3012
rect 7423 3040 7435 3043
rect 7926 3040 7932 3052
rect 7423 3012 7932 3040
rect 7423 3009 7435 3012
rect 7377 3003 7435 3009
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 8389 3043 8447 3049
rect 8389 3009 8401 3043
rect 8435 3040 8447 3043
rect 8478 3040 8484 3052
rect 8435 3012 8484 3040
rect 8435 3009 8447 3012
rect 8389 3003 8447 3009
rect 8478 3000 8484 3012
rect 8536 3000 8542 3052
rect 8849 3043 8907 3049
rect 8849 3009 8861 3043
rect 8895 3040 8907 3043
rect 8938 3040 8944 3052
rect 8895 3012 8944 3040
rect 8895 3009 8907 3012
rect 8849 3003 8907 3009
rect 8938 3000 8944 3012
rect 8996 3000 9002 3052
rect 9030 3000 9036 3052
rect 9088 3000 9094 3052
rect 9324 3049 9352 3080
rect 10134 3068 10140 3120
rect 10192 3068 10198 3120
rect 10502 3068 10508 3120
rect 10560 3108 10566 3120
rect 15562 3108 15568 3120
rect 10560 3080 15568 3108
rect 10560 3068 10566 3080
rect 15562 3068 15568 3080
rect 15620 3068 15626 3120
rect 15930 3108 15936 3120
rect 15672 3080 15936 3108
rect 9309 3043 9367 3049
rect 9309 3009 9321 3043
rect 9355 3040 9367 3043
rect 11330 3040 11336 3052
rect 9355 3012 11336 3040
rect 9355 3009 9367 3012
rect 9309 3003 9367 3009
rect 11330 3000 11336 3012
rect 11388 3000 11394 3052
rect 11606 3000 11612 3052
rect 11664 3040 11670 3052
rect 12253 3043 12311 3049
rect 12253 3040 12265 3043
rect 11664 3012 12265 3040
rect 11664 3000 11670 3012
rect 12253 3009 12265 3012
rect 12299 3009 12311 3043
rect 12253 3003 12311 3009
rect 13262 3000 13268 3052
rect 13320 3000 13326 3052
rect 13446 3000 13452 3052
rect 13504 3000 13510 3052
rect 13722 3000 13728 3052
rect 13780 3040 13786 3052
rect 14185 3043 14243 3049
rect 14185 3040 14197 3043
rect 13780 3012 14197 3040
rect 13780 3000 13786 3012
rect 14185 3009 14197 3012
rect 14231 3009 14243 3043
rect 14185 3003 14243 3009
rect 7466 2932 7472 2984
rect 7524 2932 7530 2984
rect 8110 2932 8116 2984
rect 8168 2932 8174 2984
rect 11054 2972 11060 2984
rect 8312 2944 11060 2972
rect 7653 2907 7711 2913
rect 7653 2873 7665 2907
rect 7699 2904 7711 2907
rect 8312 2904 8340 2944
rect 11054 2932 11060 2944
rect 11112 2932 11118 2984
rect 11146 2932 11152 2984
rect 11204 2972 11210 2984
rect 11701 2975 11759 2981
rect 11701 2972 11713 2975
rect 11204 2944 11713 2972
rect 11204 2932 11210 2944
rect 11701 2941 11713 2944
rect 11747 2941 11759 2975
rect 11701 2935 11759 2941
rect 12158 2932 12164 2984
rect 12216 2932 12222 2984
rect 14200 2972 14228 3003
rect 14274 3000 14280 3052
rect 14332 3040 14338 3052
rect 14550 3040 14556 3052
rect 14332 3012 14556 3040
rect 14332 3000 14338 3012
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 14918 3000 14924 3052
rect 14976 3000 14982 3052
rect 15672 3049 15700 3080
rect 15930 3068 15936 3080
rect 15988 3068 15994 3120
rect 16025 3111 16083 3117
rect 16025 3077 16037 3111
rect 16071 3108 16083 3111
rect 19518 3108 19524 3120
rect 16071 3080 19524 3108
rect 16071 3077 16083 3080
rect 16025 3071 16083 3077
rect 15657 3043 15715 3049
rect 15657 3009 15669 3043
rect 15703 3009 15715 3043
rect 15657 3003 15715 3009
rect 15838 3000 15844 3052
rect 15896 3000 15902 3052
rect 17034 3000 17040 3052
rect 17092 3000 17098 3052
rect 17129 3043 17187 3049
rect 17129 3009 17141 3043
rect 17175 3009 17187 3043
rect 17129 3003 17187 3009
rect 15194 2972 15200 2984
rect 14200 2944 15200 2972
rect 15194 2932 15200 2944
rect 15252 2932 15258 2984
rect 15562 2932 15568 2984
rect 15620 2972 15626 2984
rect 17144 2972 17172 3003
rect 17218 3000 17224 3052
rect 17276 3000 17282 3052
rect 17310 3000 17316 3052
rect 17368 3049 17374 3052
rect 17368 3043 17397 3049
rect 17385 3009 17397 3043
rect 17368 3003 17397 3009
rect 17368 3000 17374 3003
rect 17494 3000 17500 3052
rect 17552 3000 17558 3052
rect 17586 3000 17592 3052
rect 17644 3040 17650 3052
rect 18417 3043 18475 3049
rect 18417 3040 18429 3043
rect 17644 3012 18429 3040
rect 17644 3000 17650 3012
rect 18417 3009 18429 3012
rect 18463 3009 18475 3043
rect 18417 3003 18475 3009
rect 18785 3043 18843 3049
rect 18785 3009 18797 3043
rect 18831 3040 18843 3043
rect 18874 3040 18880 3052
rect 18831 3012 18880 3040
rect 18831 3009 18843 3012
rect 18785 3003 18843 3009
rect 18874 3000 18880 3012
rect 18932 3000 18938 3052
rect 19242 3000 19248 3052
rect 19300 3000 19306 3052
rect 19352 3049 19380 3080
rect 19518 3068 19524 3080
rect 19576 3068 19582 3120
rect 19628 3108 19656 3148
rect 19978 3136 19984 3188
rect 20036 3176 20042 3188
rect 20809 3179 20867 3185
rect 20809 3176 20821 3179
rect 20036 3148 20821 3176
rect 20036 3136 20042 3148
rect 20809 3145 20821 3148
rect 20855 3145 20867 3179
rect 20809 3139 20867 3145
rect 20622 3108 20628 3120
rect 19628 3080 20628 3108
rect 20622 3068 20628 3080
rect 20680 3068 20686 3120
rect 19337 3043 19395 3049
rect 19337 3009 19349 3043
rect 19383 3009 19395 3043
rect 19337 3003 19395 3009
rect 19794 3000 19800 3052
rect 19852 3000 19858 3052
rect 20441 3043 20499 3049
rect 20441 3009 20453 3043
rect 20487 3009 20499 3043
rect 20441 3003 20499 3009
rect 15620 2944 17172 2972
rect 15620 2932 15626 2944
rect 17862 2932 17868 2984
rect 17920 2972 17926 2984
rect 20456 2972 20484 3003
rect 17920 2944 20484 2972
rect 17920 2932 17926 2944
rect 7699 2876 8340 2904
rect 7699 2873 7711 2876
rect 7653 2867 7711 2873
rect 8386 2864 8392 2916
rect 8444 2904 8450 2916
rect 9217 2907 9275 2913
rect 9217 2904 9229 2907
rect 8444 2876 9229 2904
rect 8444 2864 8450 2876
rect 9217 2873 9229 2876
rect 9263 2904 9275 2907
rect 12989 2907 13047 2913
rect 12989 2904 13001 2907
rect 9263 2876 13001 2904
rect 9263 2873 9275 2876
rect 9217 2867 9275 2873
rect 12989 2873 13001 2876
rect 13035 2873 13047 2907
rect 12989 2867 13047 2873
rect 17126 2864 17132 2916
rect 17184 2904 17190 2916
rect 17880 2904 17908 2932
rect 17184 2876 17908 2904
rect 18049 2907 18107 2913
rect 17184 2864 17190 2876
rect 18049 2873 18061 2907
rect 18095 2873 18107 2907
rect 18049 2867 18107 2873
rect 4948 2808 6960 2836
rect 4948 2796 4954 2808
rect 8110 2796 8116 2848
rect 8168 2836 8174 2848
rect 8205 2839 8263 2845
rect 8205 2836 8217 2839
rect 8168 2808 8217 2836
rect 8168 2796 8174 2808
rect 8205 2805 8217 2808
rect 8251 2805 8263 2839
rect 8205 2799 8263 2805
rect 8297 2839 8355 2845
rect 8297 2805 8309 2839
rect 8343 2836 8355 2839
rect 8570 2836 8576 2848
rect 8343 2808 8576 2836
rect 8343 2805 8355 2808
rect 8297 2799 8355 2805
rect 8570 2796 8576 2808
rect 8628 2796 8634 2848
rect 9125 2839 9183 2845
rect 9125 2805 9137 2839
rect 9171 2836 9183 2839
rect 9306 2836 9312 2848
rect 9171 2808 9312 2836
rect 9171 2805 9183 2808
rect 9125 2799 9183 2805
rect 9306 2796 9312 2808
rect 9364 2796 9370 2848
rect 10502 2796 10508 2848
rect 10560 2836 10566 2848
rect 10597 2839 10655 2845
rect 10597 2836 10609 2839
rect 10560 2808 10609 2836
rect 10560 2796 10566 2808
rect 10597 2805 10609 2808
rect 10643 2805 10655 2839
rect 10597 2799 10655 2805
rect 10778 2796 10784 2848
rect 10836 2836 10842 2848
rect 17402 2836 17408 2848
rect 10836 2808 17408 2836
rect 10836 2796 10842 2808
rect 17402 2796 17408 2808
rect 17460 2796 17466 2848
rect 17770 2796 17776 2848
rect 17828 2836 17834 2848
rect 18064 2836 18092 2867
rect 19518 2864 19524 2916
rect 19576 2904 19582 2916
rect 21269 2907 21327 2913
rect 21269 2904 21281 2907
rect 19576 2876 21281 2904
rect 19576 2864 19582 2876
rect 21269 2873 21281 2876
rect 21315 2873 21327 2907
rect 21269 2867 21327 2873
rect 17828 2808 18092 2836
rect 17828 2796 17834 2808
rect 21450 2796 21456 2848
rect 21508 2836 21514 2848
rect 22005 2839 22063 2845
rect 22005 2836 22017 2839
rect 21508 2808 22017 2836
rect 21508 2796 21514 2808
rect 22005 2805 22017 2808
rect 22051 2805 22063 2839
rect 22005 2799 22063 2805
rect 22094 2796 22100 2848
rect 22152 2836 22158 2848
rect 22649 2839 22707 2845
rect 22649 2836 22661 2839
rect 22152 2808 22661 2836
rect 22152 2796 22158 2808
rect 22649 2805 22661 2808
rect 22695 2805 22707 2839
rect 22649 2799 22707 2805
rect 1104 2746 23828 2768
rect 1104 2694 3790 2746
rect 3842 2694 3854 2746
rect 3906 2694 3918 2746
rect 3970 2694 3982 2746
rect 4034 2694 4046 2746
rect 4098 2694 9471 2746
rect 9523 2694 9535 2746
rect 9587 2694 9599 2746
rect 9651 2694 9663 2746
rect 9715 2694 9727 2746
rect 9779 2694 15152 2746
rect 15204 2694 15216 2746
rect 15268 2694 15280 2746
rect 15332 2694 15344 2746
rect 15396 2694 15408 2746
rect 15460 2694 20833 2746
rect 20885 2694 20897 2746
rect 20949 2694 20961 2746
rect 21013 2694 21025 2746
rect 21077 2694 21089 2746
rect 21141 2694 23828 2746
rect 1104 2672 23828 2694
rect 4893 2635 4951 2641
rect 4893 2601 4905 2635
rect 4939 2632 4951 2635
rect 5718 2632 5724 2644
rect 4939 2604 5724 2632
rect 4939 2601 4951 2604
rect 4893 2595 4951 2601
rect 5718 2592 5724 2604
rect 5776 2592 5782 2644
rect 8389 2635 8447 2641
rect 8389 2601 8401 2635
rect 8435 2632 8447 2635
rect 8846 2632 8852 2644
rect 8435 2604 8852 2632
rect 8435 2601 8447 2604
rect 8389 2595 8447 2601
rect 8846 2592 8852 2604
rect 8904 2592 8910 2644
rect 9122 2592 9128 2644
rect 9180 2592 9186 2644
rect 12069 2635 12127 2641
rect 12069 2601 12081 2635
rect 12115 2632 12127 2635
rect 12894 2632 12900 2644
rect 12115 2604 12900 2632
rect 12115 2601 12127 2604
rect 12069 2595 12127 2601
rect 12894 2592 12900 2604
rect 12952 2592 12958 2644
rect 15746 2592 15752 2644
rect 15804 2632 15810 2644
rect 15841 2635 15899 2641
rect 15841 2632 15853 2635
rect 15804 2604 15853 2632
rect 15804 2592 15810 2604
rect 15841 2601 15853 2604
rect 15887 2601 15899 2635
rect 15841 2595 15899 2601
rect 16945 2635 17003 2641
rect 16945 2601 16957 2635
rect 16991 2632 17003 2635
rect 17034 2632 17040 2644
rect 16991 2604 17040 2632
rect 16991 2601 17003 2604
rect 16945 2595 17003 2601
rect 17034 2592 17040 2604
rect 17092 2592 17098 2644
rect 4522 2524 4528 2576
rect 4580 2524 4586 2576
rect 4614 2524 4620 2576
rect 4672 2524 4678 2576
rect 15470 2524 15476 2576
rect 15528 2524 15534 2576
rect 3142 2496 3148 2508
rect 2516 2468 3148 2496
rect 2516 2437 2544 2468
rect 3142 2456 3148 2468
rect 3200 2456 3206 2508
rect 4540 2496 4568 2524
rect 5258 2496 5264 2508
rect 4540 2468 5264 2496
rect 5258 2456 5264 2468
rect 5316 2456 5322 2508
rect 7745 2499 7803 2505
rect 7745 2465 7757 2499
rect 7791 2496 7803 2499
rect 8018 2496 8024 2508
rect 7791 2468 8024 2496
rect 7791 2465 7803 2468
rect 7745 2459 7803 2465
rect 8018 2456 8024 2468
rect 8076 2456 8082 2508
rect 8110 2456 8116 2508
rect 8168 2456 8174 2508
rect 8205 2499 8263 2505
rect 8205 2465 8217 2499
rect 8251 2496 8263 2499
rect 10686 2496 10692 2508
rect 8251 2468 10692 2496
rect 8251 2465 8263 2468
rect 8205 2459 8263 2465
rect 10686 2456 10692 2468
rect 10744 2456 10750 2508
rect 11149 2499 11207 2505
rect 11149 2465 11161 2499
rect 11195 2496 11207 2499
rect 11790 2496 11796 2508
rect 11195 2468 11796 2496
rect 11195 2465 11207 2468
rect 11149 2459 11207 2465
rect 11790 2456 11796 2468
rect 11848 2456 11854 2508
rect 14642 2456 14648 2508
rect 14700 2496 14706 2508
rect 15381 2499 15439 2505
rect 15381 2496 15393 2499
rect 14700 2468 15393 2496
rect 14700 2456 14706 2468
rect 15381 2465 15393 2468
rect 15427 2465 15439 2499
rect 15381 2459 15439 2465
rect 16574 2456 16580 2508
rect 16632 2496 16638 2508
rect 17865 2499 17923 2505
rect 17865 2496 17877 2499
rect 16632 2468 17877 2496
rect 16632 2456 16638 2468
rect 17865 2465 17877 2468
rect 17911 2465 17923 2499
rect 17865 2459 17923 2465
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 3418 2388 3424 2440
rect 3476 2388 3482 2440
rect 3694 2388 3700 2440
rect 3752 2428 3758 2440
rect 4433 2431 4491 2437
rect 4433 2428 4445 2431
rect 3752 2400 4445 2428
rect 3752 2388 3758 2400
rect 4433 2397 4445 2400
rect 4479 2397 4491 2431
rect 4433 2391 4491 2397
rect 4706 2388 4712 2440
rect 4764 2388 4770 2440
rect 5902 2388 5908 2440
rect 5960 2388 5966 2440
rect 7009 2431 7067 2437
rect 7009 2397 7021 2431
rect 7055 2428 7067 2431
rect 7098 2428 7104 2440
rect 7055 2400 7104 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 9858 2388 9864 2440
rect 9916 2388 9922 2440
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2428 10563 2431
rect 10962 2428 10968 2440
rect 10551 2400 10968 2428
rect 10551 2397 10563 2400
rect 10505 2391 10563 2397
rect 10962 2388 10968 2400
rect 11020 2388 11026 2440
rect 11422 2388 11428 2440
rect 11480 2428 11486 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11480 2400 11713 2428
rect 11480 2388 11486 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2428 11943 2431
rect 11974 2428 11980 2440
rect 11931 2400 11980 2428
rect 11931 2397 11943 2400
rect 11885 2391 11943 2397
rect 11974 2388 11980 2400
rect 12032 2388 12038 2440
rect 12529 2431 12587 2437
rect 12529 2397 12541 2431
rect 12575 2428 12587 2431
rect 12710 2428 12716 2440
rect 12575 2400 12716 2428
rect 12575 2397 12587 2400
rect 12529 2391 12587 2397
rect 12710 2388 12716 2400
rect 12768 2388 12774 2440
rect 13078 2388 13084 2440
rect 13136 2428 13142 2440
rect 13173 2431 13231 2437
rect 13173 2428 13185 2431
rect 13136 2400 13185 2428
rect 13136 2388 13142 2400
rect 13173 2397 13185 2400
rect 13219 2397 13231 2431
rect 13173 2391 13231 2397
rect 13814 2388 13820 2440
rect 13872 2428 13878 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 13872 2400 14289 2428
rect 13872 2388 13878 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 15562 2388 15568 2440
rect 15620 2428 15626 2440
rect 15657 2431 15715 2437
rect 15657 2428 15669 2431
rect 15620 2400 15669 2428
rect 15620 2388 15626 2400
rect 15657 2397 15669 2400
rect 15703 2397 15715 2431
rect 15657 2391 15715 2397
rect 17126 2388 17132 2440
rect 17184 2388 17190 2440
rect 17402 2388 17408 2440
rect 17460 2388 17466 2440
rect 18506 2388 18512 2440
rect 18564 2388 18570 2440
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 20070 2388 20076 2440
rect 20128 2388 20134 2440
rect 20714 2388 20720 2440
rect 20772 2388 20778 2440
rect 22002 2388 22008 2440
rect 22060 2388 22066 2440
rect 22646 2388 22652 2440
rect 22704 2388 22710 2440
rect 2225 2363 2283 2369
rect 2225 2329 2237 2363
rect 2271 2329 2283 2363
rect 2225 2323 2283 2329
rect 2240 2292 2268 2323
rect 3142 2320 3148 2372
rect 3200 2320 3206 2372
rect 5534 2320 5540 2372
rect 5592 2360 5598 2372
rect 5629 2363 5687 2369
rect 5629 2360 5641 2363
rect 5592 2332 5641 2360
rect 5592 2320 5598 2332
rect 5629 2329 5641 2332
rect 5675 2329 5687 2363
rect 5629 2323 5687 2329
rect 5994 2320 6000 2372
rect 6052 2360 6058 2372
rect 6733 2363 6791 2369
rect 6733 2360 6745 2363
rect 6052 2332 6745 2360
rect 6052 2320 6058 2332
rect 6733 2329 6745 2332
rect 6779 2329 6791 2363
rect 6733 2323 6791 2329
rect 16758 2320 16764 2372
rect 16816 2360 16822 2372
rect 17313 2363 17371 2369
rect 17313 2360 17325 2363
rect 16816 2332 17325 2360
rect 16816 2320 16822 2332
rect 17313 2329 17325 2332
rect 17359 2329 17371 2363
rect 17313 2323 17371 2329
rect 3418 2292 3424 2304
rect 2240 2264 3424 2292
rect 3418 2252 3424 2264
rect 3476 2252 3482 2304
rect 1104 2202 23987 2224
rect 1104 2150 6630 2202
rect 6682 2150 6694 2202
rect 6746 2150 6758 2202
rect 6810 2150 6822 2202
rect 6874 2150 6886 2202
rect 6938 2150 12311 2202
rect 12363 2150 12375 2202
rect 12427 2150 12439 2202
rect 12491 2150 12503 2202
rect 12555 2150 12567 2202
rect 12619 2150 17992 2202
rect 18044 2150 18056 2202
rect 18108 2150 18120 2202
rect 18172 2150 18184 2202
rect 18236 2150 18248 2202
rect 18300 2150 23673 2202
rect 23725 2150 23737 2202
rect 23789 2150 23801 2202
rect 23853 2150 23865 2202
rect 23917 2150 23929 2202
rect 23981 2150 23987 2202
rect 1104 2128 23987 2150
rect 7282 1028 7288 1080
rect 7340 1068 7346 1080
rect 10410 1068 10416 1080
rect 7340 1040 10416 1068
rect 7340 1028 7346 1040
rect 10410 1028 10416 1040
rect 10468 1028 10474 1080
rect 16942 1028 16948 1080
rect 17000 1068 17006 1080
rect 18506 1068 18512 1080
rect 17000 1040 18512 1068
rect 17000 1028 17006 1040
rect 18506 1028 18512 1040
rect 18564 1028 18570 1080
rect 18874 1028 18880 1080
rect 18932 1068 18938 1080
rect 20714 1068 20720 1080
rect 18932 1040 20720 1068
rect 18932 1028 18938 1040
rect 20714 1028 20720 1040
rect 20772 1028 20778 1080
rect 1486 960 1492 1012
rect 1544 1000 1550 1012
rect 5810 1000 5816 1012
rect 1544 972 5816 1000
rect 1544 960 1550 972
rect 5810 960 5816 972
rect 5868 960 5874 1012
rect 7926 960 7932 1012
rect 7984 1000 7990 1012
rect 10318 1000 10324 1012
rect 7984 972 10324 1000
rect 7984 960 7990 972
rect 10318 960 10324 972
rect 10376 960 10382 1012
rect 18230 960 18236 1012
rect 18288 1000 18294 1012
rect 20070 1000 20076 1012
rect 18288 972 20076 1000
rect 18288 960 18294 972
rect 20070 960 20076 972
rect 20128 960 20134 1012
rect 20806 960 20812 1012
rect 20864 1000 20870 1012
rect 22646 1000 22652 1012
rect 20864 972 22652 1000
rect 20864 960 20870 972
rect 22646 960 22652 972
rect 22704 960 22710 1012
rect 3142 892 3148 944
rect 3200 932 3206 944
rect 4706 932 4712 944
rect 3200 904 4712 932
rect 3200 892 3206 904
rect 4706 892 4712 904
rect 4764 892 4770 944
rect 8570 892 8576 944
rect 8628 932 8634 944
rect 9766 932 9772 944
rect 8628 904 9772 932
rect 8628 892 8634 904
rect 9766 892 9772 904
rect 9824 892 9830 944
rect 17586 892 17592 944
rect 17644 932 17650 944
rect 19426 932 19432 944
rect 17644 904 19432 932
rect 17644 892 17650 904
rect 19426 892 19432 904
rect 19484 892 19490 944
rect 20162 892 20168 944
rect 20220 932 20226 944
rect 22002 932 22008 944
rect 20220 904 22008 932
rect 20220 892 20226 904
rect 22002 892 22008 904
rect 22060 892 22066 944
<< via1 >>
rect 3790 22278 3842 22330
rect 3854 22278 3906 22330
rect 3918 22278 3970 22330
rect 3982 22278 4034 22330
rect 4046 22278 4098 22330
rect 9471 22278 9523 22330
rect 9535 22278 9587 22330
rect 9599 22278 9651 22330
rect 9663 22278 9715 22330
rect 9727 22278 9779 22330
rect 15152 22278 15204 22330
rect 15216 22278 15268 22330
rect 15280 22278 15332 22330
rect 15344 22278 15396 22330
rect 15408 22278 15460 22330
rect 20833 22278 20885 22330
rect 20897 22278 20949 22330
rect 20961 22278 21013 22330
rect 21025 22278 21077 22330
rect 21089 22278 21141 22330
rect 12716 22108 12768 22160
rect 12072 22040 12124 22092
rect 15660 22040 15712 22092
rect 2044 22015 2096 22024
rect 2044 21981 2053 22015
rect 2053 21981 2087 22015
rect 2087 21981 2096 22015
rect 2044 21972 2096 21981
rect 4528 22015 4580 22024
rect 4528 21981 4537 22015
rect 4537 21981 4571 22015
rect 4571 21981 4580 22015
rect 4528 21972 4580 21981
rect 11980 21972 12032 22024
rect 2596 21904 2648 21956
rect 7472 21904 7524 21956
rect 12532 21972 12584 22024
rect 20444 22015 20496 22024
rect 20444 21981 20453 22015
rect 20453 21981 20487 22015
rect 20487 21981 20496 22015
rect 20444 21972 20496 21981
rect 20720 21972 20772 22024
rect 3240 21836 3292 21888
rect 6092 21836 6144 21888
rect 7380 21836 7432 21888
rect 13176 21947 13228 21956
rect 13176 21913 13185 21947
rect 13185 21913 13219 21947
rect 13219 21913 13228 21947
rect 13176 21904 13228 21913
rect 17408 21904 17460 21956
rect 22652 21947 22704 21956
rect 22652 21913 22661 21947
rect 22661 21913 22695 21947
rect 22695 21913 22704 21947
rect 22652 21904 22704 21913
rect 13084 21836 13136 21888
rect 14740 21836 14792 21888
rect 15844 21836 15896 21888
rect 18880 21836 18932 21888
rect 19248 21836 19300 21888
rect 22836 21836 22888 21888
rect 6630 21734 6682 21786
rect 6694 21734 6746 21786
rect 6758 21734 6810 21786
rect 6822 21734 6874 21786
rect 6886 21734 6938 21786
rect 12311 21734 12363 21786
rect 12375 21734 12427 21786
rect 12439 21734 12491 21786
rect 12503 21734 12555 21786
rect 12567 21734 12619 21786
rect 17992 21734 18044 21786
rect 18056 21734 18108 21786
rect 18120 21734 18172 21786
rect 18184 21734 18236 21786
rect 18248 21734 18300 21786
rect 23673 21734 23725 21786
rect 23737 21734 23789 21786
rect 23801 21734 23853 21786
rect 23865 21734 23917 21786
rect 23929 21734 23981 21786
rect 3700 21564 3752 21616
rect 4528 21564 4580 21616
rect 4160 21539 4212 21548
rect 4160 21505 4169 21539
rect 4169 21505 4203 21539
rect 4203 21505 4212 21539
rect 4160 21496 4212 21505
rect 5724 21539 5776 21548
rect 19248 21675 19300 21684
rect 19248 21641 19257 21675
rect 19257 21641 19291 21675
rect 19291 21641 19300 21675
rect 19248 21632 19300 21641
rect 15016 21564 15068 21616
rect 15936 21607 15988 21616
rect 15936 21573 15945 21607
rect 15945 21573 15979 21607
rect 15979 21573 15988 21607
rect 15936 21564 15988 21573
rect 5724 21505 5742 21539
rect 5742 21505 5776 21539
rect 5724 21496 5776 21505
rect 6092 21496 6144 21548
rect 9956 21496 10008 21548
rect 12164 21496 12216 21548
rect 12440 21539 12492 21548
rect 12440 21505 12449 21539
rect 12449 21505 12483 21539
rect 12483 21505 12492 21539
rect 12440 21496 12492 21505
rect 12532 21539 12584 21548
rect 12532 21505 12541 21539
rect 12541 21505 12575 21539
rect 12575 21505 12584 21539
rect 12532 21496 12584 21505
rect 12716 21539 12768 21548
rect 12716 21505 12725 21539
rect 12725 21505 12759 21539
rect 12759 21505 12768 21539
rect 12716 21496 12768 21505
rect 13084 21496 13136 21548
rect 14188 21539 14240 21548
rect 14188 21505 14197 21539
rect 14197 21505 14231 21539
rect 14231 21505 14240 21539
rect 14188 21496 14240 21505
rect 14648 21539 14700 21548
rect 14648 21505 14657 21539
rect 14657 21505 14691 21539
rect 14691 21505 14700 21539
rect 14648 21496 14700 21505
rect 15844 21496 15896 21548
rect 17408 21496 17460 21548
rect 17868 21539 17920 21548
rect 17868 21505 17877 21539
rect 17877 21505 17911 21539
rect 17911 21505 17920 21539
rect 17868 21496 17920 21505
rect 19432 21564 19484 21616
rect 18144 21539 18196 21548
rect 18144 21505 18153 21539
rect 18153 21505 18187 21539
rect 18187 21505 18196 21539
rect 18144 21496 18196 21505
rect 19708 21496 19760 21548
rect 4436 21292 4488 21344
rect 4620 21335 4672 21344
rect 4620 21301 4629 21335
rect 4629 21301 4663 21335
rect 4663 21301 4672 21335
rect 4620 21292 4672 21301
rect 8208 21428 8260 21480
rect 13820 21428 13872 21480
rect 14096 21428 14148 21480
rect 11980 21360 12032 21412
rect 14648 21360 14700 21412
rect 14832 21360 14884 21412
rect 7196 21292 7248 21344
rect 8116 21292 8168 21344
rect 9864 21292 9916 21344
rect 13268 21292 13320 21344
rect 15752 21335 15804 21344
rect 15752 21301 15761 21335
rect 15761 21301 15795 21335
rect 15795 21301 15804 21335
rect 15752 21292 15804 21301
rect 16028 21292 16080 21344
rect 17132 21360 17184 21412
rect 18880 21471 18932 21480
rect 18880 21437 18889 21471
rect 18889 21437 18923 21471
rect 18923 21437 18932 21471
rect 18880 21428 18932 21437
rect 22284 21632 22336 21684
rect 22376 21675 22428 21684
rect 22376 21641 22385 21675
rect 22385 21641 22419 21675
rect 22419 21641 22428 21675
rect 22376 21632 22428 21641
rect 22652 21632 22704 21684
rect 20720 21607 20772 21616
rect 20720 21573 20729 21607
rect 20729 21573 20763 21607
rect 20763 21573 20772 21607
rect 20720 21564 20772 21573
rect 20260 21539 20312 21548
rect 20260 21505 20269 21539
rect 20269 21505 20303 21539
rect 20303 21505 20312 21539
rect 20260 21496 20312 21505
rect 20444 21496 20496 21548
rect 20720 21428 20772 21480
rect 3790 21190 3842 21242
rect 3854 21190 3906 21242
rect 3918 21190 3970 21242
rect 3982 21190 4034 21242
rect 4046 21190 4098 21242
rect 9471 21190 9523 21242
rect 9535 21190 9587 21242
rect 9599 21190 9651 21242
rect 9663 21190 9715 21242
rect 9727 21190 9779 21242
rect 15152 21190 15204 21242
rect 15216 21190 15268 21242
rect 15280 21190 15332 21242
rect 15344 21190 15396 21242
rect 15408 21190 15460 21242
rect 20833 21190 20885 21242
rect 20897 21190 20949 21242
rect 20961 21190 21013 21242
rect 21025 21190 21077 21242
rect 21089 21190 21141 21242
rect 14188 21088 14240 21140
rect 8392 21020 8444 21072
rect 12440 20952 12492 21004
rect 14280 21020 14332 21072
rect 15016 21088 15068 21140
rect 17132 21131 17184 21140
rect 17132 21097 17141 21131
rect 17141 21097 17175 21131
rect 17175 21097 17184 21131
rect 17132 21088 17184 21097
rect 18144 21088 18196 21140
rect 19524 21088 19576 21140
rect 17408 21063 17460 21072
rect 17408 21029 17417 21063
rect 17417 21029 17451 21063
rect 17451 21029 17460 21063
rect 17408 21020 17460 21029
rect 2044 20884 2096 20936
rect 2504 20884 2556 20936
rect 5816 20884 5868 20936
rect 7196 20927 7248 20936
rect 7196 20893 7205 20927
rect 7205 20893 7239 20927
rect 7239 20893 7248 20927
rect 7196 20884 7248 20893
rect 9128 20884 9180 20936
rect 2320 20816 2372 20868
rect 7104 20816 7156 20868
rect 2688 20748 2740 20800
rect 5632 20748 5684 20800
rect 8484 20791 8536 20800
rect 8484 20757 8493 20791
rect 8493 20757 8527 20791
rect 8527 20757 8536 20791
rect 8484 20748 8536 20757
rect 10968 20816 11020 20868
rect 11060 20748 11112 20800
rect 12716 20884 12768 20936
rect 12900 20927 12952 20936
rect 12900 20893 12909 20927
rect 12909 20893 12943 20927
rect 12943 20893 12952 20927
rect 12900 20884 12952 20893
rect 13268 20884 13320 20936
rect 14556 20927 14608 20936
rect 14556 20893 14565 20927
rect 14565 20893 14599 20927
rect 14599 20893 14608 20927
rect 14556 20884 14608 20893
rect 14740 20927 14792 20936
rect 14740 20893 14749 20927
rect 14749 20893 14783 20927
rect 14783 20893 14792 20927
rect 14740 20884 14792 20893
rect 16304 20952 16356 21004
rect 14372 20816 14424 20868
rect 15660 20884 15712 20936
rect 16212 20927 16264 20936
rect 16212 20893 16221 20927
rect 16221 20893 16255 20927
rect 16255 20893 16264 20927
rect 16212 20884 16264 20893
rect 17408 20884 17460 20936
rect 17500 20927 17552 20936
rect 17500 20893 17509 20927
rect 17509 20893 17543 20927
rect 17543 20893 17552 20927
rect 17500 20884 17552 20893
rect 17868 21020 17920 21072
rect 19340 21020 19392 21072
rect 18880 20952 18932 21004
rect 18144 20884 18196 20936
rect 14280 20748 14332 20800
rect 14924 20791 14976 20800
rect 14924 20757 14933 20791
rect 14933 20757 14967 20791
rect 14967 20757 14976 20791
rect 14924 20748 14976 20757
rect 18328 20816 18380 20868
rect 18236 20748 18288 20800
rect 19524 20884 19576 20936
rect 19616 20927 19668 20936
rect 19616 20893 19625 20927
rect 19625 20893 19659 20927
rect 19659 20893 19668 20927
rect 19616 20884 19668 20893
rect 19800 20884 19852 20936
rect 20168 20884 20220 20936
rect 20628 20884 20680 20936
rect 22652 20995 22704 21004
rect 22652 20961 22661 20995
rect 22661 20961 22695 20995
rect 22695 20961 22704 20995
rect 22652 20952 22704 20961
rect 20076 20816 20128 20868
rect 21916 20859 21968 20868
rect 21916 20825 21925 20859
rect 21925 20825 21959 20859
rect 21959 20825 21968 20859
rect 21916 20816 21968 20825
rect 20260 20748 20312 20800
rect 6630 20646 6682 20698
rect 6694 20646 6746 20698
rect 6758 20646 6810 20698
rect 6822 20646 6874 20698
rect 6886 20646 6938 20698
rect 12311 20646 12363 20698
rect 12375 20646 12427 20698
rect 12439 20646 12491 20698
rect 12503 20646 12555 20698
rect 12567 20646 12619 20698
rect 17992 20646 18044 20698
rect 18056 20646 18108 20698
rect 18120 20646 18172 20698
rect 18184 20646 18236 20698
rect 18248 20646 18300 20698
rect 23673 20646 23725 20698
rect 23737 20646 23789 20698
rect 23801 20646 23853 20698
rect 23865 20646 23917 20698
rect 23929 20646 23981 20698
rect 2044 20544 2096 20596
rect 4160 20544 4212 20596
rect 11060 20587 11112 20596
rect 11060 20553 11069 20587
rect 11069 20553 11103 20587
rect 11103 20553 11112 20587
rect 11060 20544 11112 20553
rect 13636 20544 13688 20596
rect 13084 20476 13136 20528
rect 14096 20476 14148 20528
rect 4344 20451 4396 20460
rect 4344 20417 4353 20451
rect 4353 20417 4387 20451
rect 4387 20417 4396 20451
rect 4344 20408 4396 20417
rect 11428 20408 11480 20460
rect 8208 20383 8260 20392
rect 8208 20349 8217 20383
rect 8217 20349 8251 20383
rect 8251 20349 8260 20383
rect 8208 20340 8260 20349
rect 11244 20272 11296 20324
rect 13084 20340 13136 20392
rect 13728 20451 13780 20460
rect 13728 20417 13737 20451
rect 13737 20417 13771 20451
rect 13771 20417 13780 20451
rect 13728 20408 13780 20417
rect 13820 20451 13872 20460
rect 13820 20417 13829 20451
rect 13829 20417 13863 20451
rect 13863 20417 13872 20451
rect 13820 20408 13872 20417
rect 14280 20451 14332 20460
rect 14280 20417 14289 20451
rect 14289 20417 14323 20451
rect 14323 20417 14332 20451
rect 14280 20408 14332 20417
rect 15200 20476 15252 20528
rect 14924 20408 14976 20460
rect 18328 20544 18380 20596
rect 20720 20587 20772 20596
rect 20720 20553 20729 20587
rect 20729 20553 20763 20587
rect 20763 20553 20772 20587
rect 20720 20544 20772 20553
rect 22652 20587 22704 20596
rect 22652 20553 22661 20587
rect 22661 20553 22695 20587
rect 22695 20553 22704 20587
rect 22652 20544 22704 20553
rect 15660 20476 15712 20528
rect 16396 20476 16448 20528
rect 15752 20408 15804 20460
rect 20260 20476 20312 20528
rect 15568 20340 15620 20392
rect 22008 20451 22060 20460
rect 22008 20417 22017 20451
rect 22017 20417 22051 20451
rect 22051 20417 22060 20451
rect 22008 20408 22060 20417
rect 22284 20408 22336 20460
rect 22836 20451 22888 20460
rect 22836 20417 22845 20451
rect 22845 20417 22879 20451
rect 22879 20417 22888 20451
rect 22836 20408 22888 20417
rect 22560 20340 22612 20392
rect 15752 20272 15804 20324
rect 16120 20272 16172 20324
rect 20168 20272 20220 20324
rect 20536 20272 20588 20324
rect 9128 20204 9180 20256
rect 11060 20204 11112 20256
rect 14924 20247 14976 20256
rect 14924 20213 14933 20247
rect 14933 20213 14967 20247
rect 14967 20213 14976 20247
rect 14924 20204 14976 20213
rect 3790 20102 3842 20154
rect 3854 20102 3906 20154
rect 3918 20102 3970 20154
rect 3982 20102 4034 20154
rect 4046 20102 4098 20154
rect 9471 20102 9523 20154
rect 9535 20102 9587 20154
rect 9599 20102 9651 20154
rect 9663 20102 9715 20154
rect 9727 20102 9779 20154
rect 15152 20102 15204 20154
rect 15216 20102 15268 20154
rect 15280 20102 15332 20154
rect 15344 20102 15396 20154
rect 15408 20102 15460 20154
rect 20833 20102 20885 20154
rect 20897 20102 20949 20154
rect 20961 20102 21013 20154
rect 21025 20102 21077 20154
rect 21089 20102 21141 20154
rect 11428 20043 11480 20052
rect 11428 20009 11437 20043
rect 11437 20009 11471 20043
rect 11471 20009 11480 20043
rect 11428 20000 11480 20009
rect 12072 20000 12124 20052
rect 14280 20000 14332 20052
rect 4160 19864 4212 19916
rect 7196 19839 7248 19848
rect 7196 19805 7205 19839
rect 7205 19805 7239 19839
rect 7239 19805 7248 19839
rect 7196 19796 7248 19805
rect 8208 19796 8260 19848
rect 9128 19839 9180 19848
rect 9128 19805 9137 19839
rect 9137 19805 9171 19839
rect 9171 19805 9180 19839
rect 9128 19796 9180 19805
rect 11336 19796 11388 19848
rect 15016 20000 15068 20052
rect 15568 20043 15620 20052
rect 15568 20009 15577 20043
rect 15577 20009 15611 20043
rect 15611 20009 15620 20043
rect 15568 20000 15620 20009
rect 19432 20043 19484 20052
rect 19432 20009 19441 20043
rect 19441 20009 19475 20043
rect 19475 20009 19484 20043
rect 19432 20000 19484 20009
rect 14556 19932 14608 19984
rect 22284 19932 22336 19984
rect 11980 19864 12032 19916
rect 15108 19907 15160 19916
rect 15108 19873 15117 19907
rect 15117 19873 15151 19907
rect 15151 19873 15160 19907
rect 15108 19864 15160 19873
rect 15660 19864 15712 19916
rect 16120 19864 16172 19916
rect 2964 19728 3016 19780
rect 6184 19728 6236 19780
rect 8484 19728 8536 19780
rect 2412 19660 2464 19712
rect 5356 19703 5408 19712
rect 5356 19669 5365 19703
rect 5365 19669 5399 19703
rect 5399 19669 5408 19703
rect 5356 19660 5408 19669
rect 9220 19660 9272 19712
rect 10324 19660 10376 19712
rect 13452 19839 13504 19848
rect 13452 19805 13461 19839
rect 13461 19805 13495 19839
rect 13495 19805 13504 19839
rect 13452 19796 13504 19805
rect 14372 19839 14424 19848
rect 14372 19805 14381 19839
rect 14381 19805 14415 19839
rect 14415 19805 14424 19839
rect 14372 19796 14424 19805
rect 14556 19839 14608 19848
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 17408 19796 17460 19848
rect 18328 19796 18380 19848
rect 22008 19864 22060 19916
rect 20076 19796 20128 19848
rect 16304 19728 16356 19780
rect 13912 19660 13964 19712
rect 14464 19703 14516 19712
rect 14464 19669 14473 19703
rect 14473 19669 14507 19703
rect 14507 19669 14516 19703
rect 14464 19660 14516 19669
rect 18788 19660 18840 19712
rect 6630 19558 6682 19610
rect 6694 19558 6746 19610
rect 6758 19558 6810 19610
rect 6822 19558 6874 19610
rect 6886 19558 6938 19610
rect 12311 19558 12363 19610
rect 12375 19558 12427 19610
rect 12439 19558 12491 19610
rect 12503 19558 12555 19610
rect 12567 19558 12619 19610
rect 17992 19558 18044 19610
rect 18056 19558 18108 19610
rect 18120 19558 18172 19610
rect 18184 19558 18236 19610
rect 18248 19558 18300 19610
rect 23673 19558 23725 19610
rect 23737 19558 23789 19610
rect 23801 19558 23853 19610
rect 23865 19558 23917 19610
rect 23929 19558 23981 19610
rect 10692 19456 10744 19508
rect 12900 19456 12952 19508
rect 16212 19456 16264 19508
rect 17500 19456 17552 19508
rect 4620 19431 4672 19440
rect 4620 19397 4629 19431
rect 4629 19397 4663 19431
rect 4663 19397 4672 19431
rect 4620 19388 4672 19397
rect 12440 19388 12492 19440
rect 13728 19388 13780 19440
rect 4160 19320 4212 19372
rect 4344 19320 4396 19372
rect 7656 19320 7708 19372
rect 8208 19363 8260 19372
rect 8208 19329 8217 19363
rect 8217 19329 8251 19363
rect 8251 19329 8260 19363
rect 8208 19320 8260 19329
rect 5264 19252 5316 19304
rect 11336 19320 11388 19372
rect 11704 19320 11756 19372
rect 12624 19363 12676 19372
rect 12624 19329 12633 19363
rect 12633 19329 12667 19363
rect 12667 19329 12676 19363
rect 12624 19320 12676 19329
rect 12900 19320 12952 19372
rect 15108 19388 15160 19440
rect 18512 19456 18564 19508
rect 18788 19456 18840 19508
rect 22008 19456 22060 19508
rect 18604 19388 18656 19440
rect 18880 19388 18932 19440
rect 14556 19320 14608 19372
rect 12440 19252 12492 19304
rect 12532 19295 12584 19304
rect 12532 19261 12540 19295
rect 12540 19261 12574 19295
rect 12574 19261 12584 19295
rect 12532 19252 12584 19261
rect 14740 19295 14792 19304
rect 14740 19261 14749 19295
rect 14749 19261 14783 19295
rect 14783 19261 14792 19295
rect 14740 19252 14792 19261
rect 16212 19252 16264 19304
rect 17132 19252 17184 19304
rect 17224 19295 17276 19304
rect 17224 19261 17233 19295
rect 17233 19261 17267 19295
rect 17267 19261 17276 19295
rect 17224 19252 17276 19261
rect 17408 19295 17460 19304
rect 17408 19261 17417 19295
rect 17417 19261 17451 19295
rect 17451 19261 17460 19295
rect 17408 19252 17460 19261
rect 17960 19320 18012 19372
rect 12992 19184 13044 19236
rect 13544 19227 13596 19236
rect 13544 19193 13553 19227
rect 13553 19193 13587 19227
rect 13587 19193 13596 19227
rect 13544 19184 13596 19193
rect 14004 19184 14056 19236
rect 16028 19184 16080 19236
rect 18512 19295 18564 19304
rect 18512 19261 18521 19295
rect 18521 19261 18555 19295
rect 18555 19261 18564 19295
rect 18512 19252 18564 19261
rect 19616 19320 19668 19372
rect 19708 19363 19760 19372
rect 19708 19329 19717 19363
rect 19717 19329 19751 19363
rect 19751 19329 19760 19363
rect 19708 19320 19760 19329
rect 20076 19320 20128 19372
rect 21180 19252 21232 19304
rect 19432 19184 19484 19236
rect 14556 19159 14608 19168
rect 14556 19125 14565 19159
rect 14565 19125 14599 19159
rect 14599 19125 14608 19159
rect 14556 19116 14608 19125
rect 14832 19116 14884 19168
rect 15568 19116 15620 19168
rect 15936 19116 15988 19168
rect 22284 19159 22336 19168
rect 22284 19125 22293 19159
rect 22293 19125 22327 19159
rect 22327 19125 22336 19159
rect 22284 19116 22336 19125
rect 3790 19014 3842 19066
rect 3854 19014 3906 19066
rect 3918 19014 3970 19066
rect 3982 19014 4034 19066
rect 4046 19014 4098 19066
rect 9471 19014 9523 19066
rect 9535 19014 9587 19066
rect 9599 19014 9651 19066
rect 9663 19014 9715 19066
rect 9727 19014 9779 19066
rect 15152 19014 15204 19066
rect 15216 19014 15268 19066
rect 15280 19014 15332 19066
rect 15344 19014 15396 19066
rect 15408 19014 15460 19066
rect 20833 19014 20885 19066
rect 20897 19014 20949 19066
rect 20961 19014 21013 19066
rect 21025 19014 21077 19066
rect 21089 19014 21141 19066
rect 5816 18955 5868 18964
rect 5816 18921 5825 18955
rect 5825 18921 5859 18955
rect 5859 18921 5868 18955
rect 5816 18912 5868 18921
rect 7656 18955 7708 18964
rect 7656 18921 7665 18955
rect 7665 18921 7699 18955
rect 7699 18921 7708 18955
rect 7656 18912 7708 18921
rect 13820 18912 13872 18964
rect 14556 18912 14608 18964
rect 18880 18955 18932 18964
rect 18880 18921 18889 18955
rect 18889 18921 18923 18955
rect 18923 18921 18932 18955
rect 18880 18912 18932 18921
rect 19432 18955 19484 18964
rect 19432 18921 19441 18955
rect 19441 18921 19475 18955
rect 19475 18921 19484 18955
rect 19432 18912 19484 18921
rect 12716 18844 12768 18896
rect 16028 18844 16080 18896
rect 2044 18819 2096 18828
rect 2044 18785 2053 18819
rect 2053 18785 2087 18819
rect 2087 18785 2096 18819
rect 2044 18776 2096 18785
rect 12624 18776 12676 18828
rect 12992 18819 13044 18828
rect 12992 18785 13001 18819
rect 13001 18785 13035 18819
rect 13035 18785 13044 18819
rect 12992 18776 13044 18785
rect 17224 18776 17276 18828
rect 5816 18708 5868 18760
rect 9128 18751 9180 18760
rect 9128 18717 9137 18751
rect 9137 18717 9171 18751
rect 9171 18717 9180 18751
rect 9128 18708 9180 18717
rect 12808 18751 12860 18760
rect 12808 18717 12817 18751
rect 12817 18717 12851 18751
rect 12851 18717 12860 18751
rect 12808 18708 12860 18717
rect 13084 18751 13136 18760
rect 13084 18717 13093 18751
rect 13093 18717 13127 18751
rect 13127 18717 13136 18751
rect 13084 18708 13136 18717
rect 14464 18751 14516 18760
rect 14464 18717 14473 18751
rect 14473 18717 14507 18751
rect 14507 18717 14516 18751
rect 14464 18708 14516 18717
rect 16764 18708 16816 18760
rect 18512 18776 18564 18828
rect 18236 18751 18288 18760
rect 18236 18717 18245 18751
rect 18245 18717 18279 18751
rect 18279 18717 18288 18751
rect 18236 18708 18288 18717
rect 18420 18751 18472 18760
rect 18420 18717 18427 18751
rect 18427 18717 18472 18751
rect 18420 18708 18472 18717
rect 18696 18844 18748 18896
rect 19524 18776 19576 18828
rect 18880 18708 18932 18760
rect 3332 18640 3384 18692
rect 12072 18640 12124 18692
rect 14556 18683 14608 18692
rect 14556 18649 14565 18683
rect 14565 18649 14599 18683
rect 14599 18649 14608 18683
rect 14556 18640 14608 18649
rect 14648 18683 14700 18692
rect 14648 18649 14657 18683
rect 14657 18649 14691 18683
rect 14691 18649 14700 18683
rect 14648 18640 14700 18649
rect 15108 18640 15160 18692
rect 17316 18640 17368 18692
rect 19984 18708 20036 18760
rect 20444 18708 20496 18760
rect 5448 18572 5500 18624
rect 10968 18572 11020 18624
rect 12532 18572 12584 18624
rect 13176 18572 13228 18624
rect 13268 18615 13320 18624
rect 13268 18581 13277 18615
rect 13277 18581 13311 18615
rect 13311 18581 13320 18615
rect 13268 18572 13320 18581
rect 13912 18572 13964 18624
rect 17592 18572 17644 18624
rect 19800 18572 19852 18624
rect 20168 18572 20220 18624
rect 6630 18470 6682 18522
rect 6694 18470 6746 18522
rect 6758 18470 6810 18522
rect 6822 18470 6874 18522
rect 6886 18470 6938 18522
rect 12311 18470 12363 18522
rect 12375 18470 12427 18522
rect 12439 18470 12491 18522
rect 12503 18470 12555 18522
rect 12567 18470 12619 18522
rect 17992 18470 18044 18522
rect 18056 18470 18108 18522
rect 18120 18470 18172 18522
rect 18184 18470 18236 18522
rect 18248 18470 18300 18522
rect 23673 18470 23725 18522
rect 23737 18470 23789 18522
rect 23801 18470 23853 18522
rect 23865 18470 23917 18522
rect 23929 18470 23981 18522
rect 9128 18411 9180 18420
rect 9128 18377 9137 18411
rect 9137 18377 9171 18411
rect 9171 18377 9180 18411
rect 9128 18368 9180 18377
rect 12072 18411 12124 18420
rect 12072 18377 12081 18411
rect 12081 18377 12115 18411
rect 12115 18377 12124 18411
rect 12072 18368 12124 18377
rect 13912 18368 13964 18420
rect 15108 18368 15160 18420
rect 15476 18368 15528 18420
rect 16764 18368 16816 18420
rect 3516 18300 3568 18352
rect 7656 18232 7708 18284
rect 12992 18300 13044 18352
rect 13268 18300 13320 18352
rect 3056 18207 3108 18216
rect 3056 18173 3065 18207
rect 3065 18173 3099 18207
rect 3099 18173 3108 18207
rect 3056 18164 3108 18173
rect 12072 18164 12124 18216
rect 12716 18232 12768 18284
rect 13544 18232 13596 18284
rect 5080 18028 5132 18080
rect 14096 18164 14148 18216
rect 14280 18232 14332 18284
rect 14832 18232 14884 18284
rect 15476 18232 15528 18284
rect 16028 18232 16080 18284
rect 17500 18368 17552 18420
rect 18328 18368 18380 18420
rect 18420 18368 18472 18420
rect 19340 18368 19392 18420
rect 17408 18300 17460 18352
rect 17776 18232 17828 18284
rect 15016 18207 15068 18216
rect 15016 18173 15025 18207
rect 15025 18173 15059 18207
rect 15059 18173 15068 18207
rect 15016 18164 15068 18173
rect 15108 18164 15160 18216
rect 19800 18300 19852 18352
rect 20260 18300 20312 18352
rect 19892 18275 19944 18284
rect 19892 18241 19901 18275
rect 19901 18241 19935 18275
rect 19935 18241 19944 18275
rect 19892 18232 19944 18241
rect 20076 18232 20128 18284
rect 14188 18096 14240 18148
rect 20720 18164 20772 18216
rect 14004 18028 14056 18080
rect 14740 18028 14792 18080
rect 15108 18028 15160 18080
rect 15476 18028 15528 18080
rect 17960 18096 18012 18148
rect 19156 18096 19208 18148
rect 17408 18028 17460 18080
rect 17868 18071 17920 18080
rect 17868 18037 17877 18071
rect 17877 18037 17911 18071
rect 17911 18037 17920 18071
rect 17868 18028 17920 18037
rect 18328 18028 18380 18080
rect 3790 17926 3842 17978
rect 3854 17926 3906 17978
rect 3918 17926 3970 17978
rect 3982 17926 4034 17978
rect 4046 17926 4098 17978
rect 9471 17926 9523 17978
rect 9535 17926 9587 17978
rect 9599 17926 9651 17978
rect 9663 17926 9715 17978
rect 9727 17926 9779 17978
rect 15152 17926 15204 17978
rect 15216 17926 15268 17978
rect 15280 17926 15332 17978
rect 15344 17926 15396 17978
rect 15408 17926 15460 17978
rect 20833 17926 20885 17978
rect 20897 17926 20949 17978
rect 20961 17926 21013 17978
rect 21025 17926 21077 17978
rect 21089 17926 21141 17978
rect 11704 17867 11756 17876
rect 11704 17833 11713 17867
rect 11713 17833 11747 17867
rect 11747 17833 11756 17867
rect 11704 17824 11756 17833
rect 13176 17867 13228 17876
rect 13176 17833 13185 17867
rect 13185 17833 13219 17867
rect 13219 17833 13228 17867
rect 13176 17824 13228 17833
rect 13268 17824 13320 17876
rect 20444 17824 20496 17876
rect 14556 17756 14608 17808
rect 15936 17756 15988 17808
rect 17316 17756 17368 17808
rect 13544 17731 13596 17740
rect 6552 17620 6604 17672
rect 9128 17663 9180 17672
rect 9128 17629 9137 17663
rect 9137 17629 9171 17663
rect 9171 17629 9180 17663
rect 9128 17620 9180 17629
rect 11612 17663 11664 17672
rect 11612 17629 11621 17663
rect 11621 17629 11655 17663
rect 11655 17629 11664 17663
rect 11612 17620 11664 17629
rect 11888 17620 11940 17672
rect 13544 17697 13553 17731
rect 13553 17697 13587 17731
rect 13587 17697 13596 17731
rect 13544 17688 13596 17697
rect 14188 17688 14240 17740
rect 14648 17688 14700 17740
rect 15200 17688 15252 17740
rect 16028 17688 16080 17740
rect 17592 17731 17644 17740
rect 17592 17697 17601 17731
rect 17601 17697 17635 17731
rect 17635 17697 17644 17731
rect 17592 17688 17644 17697
rect 12716 17620 12768 17672
rect 13360 17663 13412 17672
rect 13360 17629 13369 17663
rect 13369 17629 13403 17663
rect 13403 17629 13412 17663
rect 13360 17620 13412 17629
rect 7472 17552 7524 17604
rect 13820 17620 13872 17672
rect 14280 17620 14332 17672
rect 15016 17663 15068 17672
rect 15016 17629 15025 17663
rect 15025 17629 15059 17663
rect 15059 17629 15068 17663
rect 15016 17620 15068 17629
rect 15660 17663 15712 17672
rect 15660 17629 15669 17663
rect 15669 17629 15703 17663
rect 15703 17629 15712 17663
rect 15660 17620 15712 17629
rect 16212 17620 16264 17672
rect 6092 17484 6144 17536
rect 8024 17484 8076 17536
rect 11520 17484 11572 17536
rect 13728 17552 13780 17604
rect 15568 17552 15620 17604
rect 16580 17663 16632 17672
rect 16580 17629 16589 17663
rect 16589 17629 16623 17663
rect 16623 17629 16632 17663
rect 16580 17620 16632 17629
rect 16856 17663 16908 17672
rect 16856 17629 16865 17663
rect 16865 17629 16899 17663
rect 16899 17629 16908 17663
rect 16856 17620 16908 17629
rect 16672 17552 16724 17604
rect 14924 17484 14976 17536
rect 15660 17484 15712 17536
rect 16028 17484 16080 17536
rect 16120 17484 16172 17536
rect 22560 17824 22612 17876
rect 22192 17663 22244 17672
rect 22192 17629 22201 17663
rect 22201 17629 22235 17663
rect 22235 17629 22244 17663
rect 22192 17620 22244 17629
rect 22284 17663 22336 17672
rect 22284 17629 22293 17663
rect 22293 17629 22327 17663
rect 22327 17629 22336 17663
rect 22284 17620 22336 17629
rect 22376 17663 22428 17672
rect 22376 17629 22385 17663
rect 22385 17629 22419 17663
rect 22419 17629 22428 17663
rect 22376 17620 22428 17629
rect 17224 17552 17276 17604
rect 6630 17382 6682 17434
rect 6694 17382 6746 17434
rect 6758 17382 6810 17434
rect 6822 17382 6874 17434
rect 6886 17382 6938 17434
rect 12311 17382 12363 17434
rect 12375 17382 12427 17434
rect 12439 17382 12491 17434
rect 12503 17382 12555 17434
rect 12567 17382 12619 17434
rect 17992 17382 18044 17434
rect 18056 17382 18108 17434
rect 18120 17382 18172 17434
rect 18184 17382 18236 17434
rect 18248 17382 18300 17434
rect 23673 17382 23725 17434
rect 23737 17382 23789 17434
rect 23801 17382 23853 17434
rect 23865 17382 23917 17434
rect 23929 17382 23981 17434
rect 11336 17280 11388 17332
rect 12716 17280 12768 17332
rect 13084 17280 13136 17332
rect 13360 17280 13412 17332
rect 13820 17280 13872 17332
rect 11888 17212 11940 17264
rect 14924 17280 14976 17332
rect 16304 17280 16356 17332
rect 16672 17280 16724 17332
rect 17960 17280 18012 17332
rect 18880 17280 18932 17332
rect 19616 17280 19668 17332
rect 19708 17280 19760 17332
rect 3056 17144 3108 17196
rect 7932 17144 7984 17196
rect 10600 17144 10652 17196
rect 13176 17144 13228 17196
rect 2228 17076 2280 17128
rect 6552 17119 6604 17128
rect 6552 17085 6561 17119
rect 6561 17085 6595 17119
rect 6595 17085 6604 17119
rect 6552 17076 6604 17085
rect 8484 17119 8536 17128
rect 8484 17085 8493 17119
rect 8493 17085 8527 17119
rect 8527 17085 8536 17119
rect 8484 17076 8536 17085
rect 12808 17076 12860 17128
rect 13360 17187 13412 17196
rect 13360 17153 13369 17187
rect 13369 17153 13403 17187
rect 13403 17153 13412 17187
rect 13360 17144 13412 17153
rect 13820 17187 13872 17196
rect 13820 17153 13829 17187
rect 13829 17153 13863 17187
rect 13863 17153 13872 17187
rect 13820 17144 13872 17153
rect 14004 17187 14056 17196
rect 14004 17153 14013 17187
rect 14013 17153 14047 17187
rect 14047 17153 14056 17187
rect 14004 17144 14056 17153
rect 14372 17144 14424 17196
rect 16856 17212 16908 17264
rect 17316 17212 17368 17264
rect 19156 17212 19208 17264
rect 15200 17187 15252 17196
rect 15200 17153 15202 17187
rect 15202 17153 15236 17187
rect 15236 17153 15252 17187
rect 14464 17076 14516 17128
rect 15200 17144 15252 17153
rect 16120 17187 16172 17196
rect 16120 17153 16129 17187
rect 16129 17153 16163 17187
rect 16163 17153 16172 17187
rect 16120 17144 16172 17153
rect 18880 17144 18932 17196
rect 19248 17187 19300 17196
rect 19248 17153 19257 17187
rect 19257 17153 19291 17187
rect 19291 17153 19300 17187
rect 19248 17144 19300 17153
rect 19800 17144 19852 17196
rect 17500 17076 17552 17128
rect 17684 17076 17736 17128
rect 12992 17008 13044 17060
rect 13176 17008 13228 17060
rect 13544 17008 13596 17060
rect 15108 17008 15160 17060
rect 4528 16983 4580 16992
rect 4528 16949 4537 16983
rect 4537 16949 4571 16983
rect 4571 16949 4580 16983
rect 4528 16940 4580 16949
rect 8852 16940 8904 16992
rect 10232 16940 10284 16992
rect 12532 16940 12584 16992
rect 14556 16983 14608 16992
rect 14556 16949 14565 16983
rect 14565 16949 14599 16983
rect 14599 16949 14608 16983
rect 14556 16940 14608 16949
rect 15016 16940 15068 16992
rect 21824 17076 21876 17128
rect 22376 17187 22428 17196
rect 22376 17153 22385 17187
rect 22385 17153 22419 17187
rect 22419 17153 22428 17187
rect 22376 17144 22428 17153
rect 22284 17076 22336 17128
rect 21180 17008 21232 17060
rect 21272 17008 21324 17060
rect 3790 16838 3842 16890
rect 3854 16838 3906 16890
rect 3918 16838 3970 16890
rect 3982 16838 4034 16890
rect 4046 16838 4098 16890
rect 9471 16838 9523 16890
rect 9535 16838 9587 16890
rect 9599 16838 9651 16890
rect 9663 16838 9715 16890
rect 9727 16838 9779 16890
rect 15152 16838 15204 16890
rect 15216 16838 15268 16890
rect 15280 16838 15332 16890
rect 15344 16838 15396 16890
rect 15408 16838 15460 16890
rect 20833 16838 20885 16890
rect 20897 16838 20949 16890
rect 20961 16838 21013 16890
rect 21025 16838 21077 16890
rect 21089 16838 21141 16890
rect 8024 16736 8076 16788
rect 13084 16736 13136 16788
rect 11336 16711 11388 16720
rect 11336 16677 11345 16711
rect 11345 16677 11379 16711
rect 11379 16677 11388 16711
rect 11336 16668 11388 16677
rect 6552 16600 6604 16652
rect 8484 16600 8536 16652
rect 9128 16643 9180 16652
rect 9128 16609 9137 16643
rect 9137 16609 9171 16643
rect 9171 16609 9180 16643
rect 9128 16600 9180 16609
rect 12532 16643 12584 16652
rect 12532 16609 12541 16643
rect 12541 16609 12575 16643
rect 12575 16609 12584 16643
rect 12532 16600 12584 16609
rect 14372 16668 14424 16720
rect 7748 16532 7800 16584
rect 8024 16575 8076 16584
rect 8024 16541 8033 16575
rect 8033 16541 8067 16575
rect 8067 16541 8076 16575
rect 8024 16532 8076 16541
rect 12808 16643 12860 16652
rect 12808 16609 12817 16643
rect 12817 16609 12851 16643
rect 12851 16609 12860 16643
rect 12808 16600 12860 16609
rect 12900 16600 12952 16652
rect 13268 16600 13320 16652
rect 16764 16600 16816 16652
rect 17316 16600 17368 16652
rect 16488 16532 16540 16584
rect 16856 16532 16908 16584
rect 22284 16779 22336 16788
rect 22284 16745 22293 16779
rect 22293 16745 22327 16779
rect 22327 16745 22336 16779
rect 22284 16736 22336 16745
rect 17960 16668 18012 16720
rect 17776 16600 17828 16652
rect 18788 16600 18840 16652
rect 20352 16668 20404 16720
rect 17500 16575 17552 16584
rect 17500 16541 17509 16575
rect 17509 16541 17543 16575
rect 17543 16541 17552 16575
rect 17500 16532 17552 16541
rect 18604 16532 18656 16584
rect 21180 16600 21232 16652
rect 3056 16464 3108 16516
rect 3608 16464 3660 16516
rect 6276 16464 6328 16516
rect 11704 16464 11756 16516
rect 1492 16396 1544 16448
rect 3424 16396 3476 16448
rect 11428 16396 11480 16448
rect 14004 16464 14056 16516
rect 14924 16464 14976 16516
rect 15844 16464 15896 16516
rect 16948 16464 17000 16516
rect 17040 16507 17092 16516
rect 17040 16473 17049 16507
rect 17049 16473 17083 16507
rect 17083 16473 17092 16507
rect 17040 16464 17092 16473
rect 18696 16464 18748 16516
rect 12164 16396 12216 16448
rect 15384 16396 15436 16448
rect 17776 16396 17828 16448
rect 19524 16396 19576 16448
rect 19892 16464 19944 16516
rect 21456 16396 21508 16448
rect 6630 16294 6682 16346
rect 6694 16294 6746 16346
rect 6758 16294 6810 16346
rect 6822 16294 6874 16346
rect 6886 16294 6938 16346
rect 12311 16294 12363 16346
rect 12375 16294 12427 16346
rect 12439 16294 12491 16346
rect 12503 16294 12555 16346
rect 12567 16294 12619 16346
rect 17992 16294 18044 16346
rect 18056 16294 18108 16346
rect 18120 16294 18172 16346
rect 18184 16294 18236 16346
rect 18248 16294 18300 16346
rect 23673 16294 23725 16346
rect 23737 16294 23789 16346
rect 23801 16294 23853 16346
rect 23865 16294 23917 16346
rect 23929 16294 23981 16346
rect 9128 16235 9180 16244
rect 9128 16201 9137 16235
rect 9137 16201 9171 16235
rect 9171 16201 9180 16235
rect 9128 16192 9180 16201
rect 15752 16192 15804 16244
rect 4344 16167 4396 16176
rect 4344 16133 4353 16167
rect 4353 16133 4387 16167
rect 4387 16133 4396 16167
rect 4344 16124 4396 16133
rect 7656 16124 7708 16176
rect 11704 16124 11756 16176
rect 18696 16192 18748 16244
rect 20444 16192 20496 16244
rect 20720 16235 20772 16244
rect 20720 16201 20729 16235
rect 20729 16201 20763 16235
rect 20763 16201 20772 16235
rect 20720 16192 20772 16201
rect 22376 16235 22428 16244
rect 22376 16201 22385 16235
rect 22385 16201 22419 16235
rect 22419 16201 22428 16235
rect 22376 16192 22428 16201
rect 12164 16056 12216 16108
rect 15568 16099 15620 16108
rect 15568 16065 15577 16099
rect 15577 16065 15611 16099
rect 15611 16065 15620 16099
rect 15568 16056 15620 16065
rect 15660 16099 15712 16108
rect 15660 16065 15669 16099
rect 15669 16065 15703 16099
rect 15703 16065 15712 16099
rect 15660 16056 15712 16065
rect 16396 16056 16448 16108
rect 17040 16056 17092 16108
rect 17224 16056 17276 16108
rect 17592 16099 17644 16108
rect 17592 16065 17601 16099
rect 17601 16065 17635 16099
rect 17635 16065 17644 16099
rect 17592 16056 17644 16065
rect 18972 16056 19024 16108
rect 13636 15988 13688 16040
rect 15016 15988 15068 16040
rect 19064 16031 19116 16040
rect 19064 15997 19073 16031
rect 19073 15997 19107 16031
rect 19107 15997 19116 16031
rect 20260 16099 20312 16108
rect 20260 16065 20269 16099
rect 20269 16065 20303 16099
rect 20303 16065 20312 16099
rect 20260 16056 20312 16065
rect 20628 16056 20680 16108
rect 22928 16099 22980 16108
rect 22928 16065 22937 16099
rect 22937 16065 22971 16099
rect 22971 16065 22980 16099
rect 22928 16056 22980 16065
rect 19064 15988 19116 15997
rect 12624 15920 12676 15972
rect 19156 15920 19208 15972
rect 19892 15920 19944 15972
rect 3056 15895 3108 15904
rect 3056 15861 3065 15895
rect 3065 15861 3099 15895
rect 3099 15861 3108 15895
rect 3056 15852 3108 15861
rect 11244 15852 11296 15904
rect 12348 15852 12400 15904
rect 13912 15895 13964 15904
rect 13912 15861 13921 15895
rect 13921 15861 13955 15895
rect 13955 15861 13964 15895
rect 13912 15852 13964 15861
rect 17040 15852 17092 15904
rect 17316 15852 17368 15904
rect 17684 15852 17736 15904
rect 20536 15852 20588 15904
rect 20720 15852 20772 15904
rect 22376 15852 22428 15904
rect 3790 15750 3842 15802
rect 3854 15750 3906 15802
rect 3918 15750 3970 15802
rect 3982 15750 4034 15802
rect 4046 15750 4098 15802
rect 9471 15750 9523 15802
rect 9535 15750 9587 15802
rect 9599 15750 9651 15802
rect 9663 15750 9715 15802
rect 9727 15750 9779 15802
rect 15152 15750 15204 15802
rect 15216 15750 15268 15802
rect 15280 15750 15332 15802
rect 15344 15750 15396 15802
rect 15408 15750 15460 15802
rect 20833 15750 20885 15802
rect 20897 15750 20949 15802
rect 20961 15750 21013 15802
rect 21025 15750 21077 15802
rect 21089 15750 21141 15802
rect 12072 15648 12124 15700
rect 13452 15648 13504 15700
rect 10600 15580 10652 15632
rect 6552 15512 6604 15564
rect 9128 15555 9180 15564
rect 9128 15521 9137 15555
rect 9137 15521 9171 15555
rect 9171 15521 9180 15555
rect 9128 15512 9180 15521
rect 12164 15512 12216 15564
rect 12440 15512 12492 15564
rect 2412 15487 2464 15496
rect 2412 15453 2421 15487
rect 2421 15453 2455 15487
rect 2455 15453 2464 15487
rect 2412 15444 2464 15453
rect 4528 15444 4580 15496
rect 4988 15444 5040 15496
rect 8300 15444 8352 15496
rect 5172 15376 5224 15428
rect 11060 15376 11112 15428
rect 2504 15308 2556 15360
rect 10140 15308 10192 15360
rect 10416 15308 10468 15360
rect 11336 15444 11388 15496
rect 11704 15444 11756 15496
rect 13360 15487 13412 15496
rect 13360 15453 13369 15487
rect 13369 15453 13403 15487
rect 13403 15453 13412 15487
rect 13360 15444 13412 15453
rect 12624 15376 12676 15428
rect 13636 15487 13688 15496
rect 13636 15453 13645 15487
rect 13645 15453 13679 15487
rect 13679 15453 13688 15487
rect 13636 15444 13688 15453
rect 15016 15555 15068 15564
rect 15016 15521 15025 15555
rect 15025 15521 15059 15555
rect 15059 15521 15068 15555
rect 15016 15512 15068 15521
rect 14280 15444 14332 15496
rect 15476 15444 15528 15496
rect 17040 15691 17092 15700
rect 17040 15657 17049 15691
rect 17049 15657 17083 15691
rect 17083 15657 17092 15691
rect 17040 15648 17092 15657
rect 17500 15580 17552 15632
rect 15844 15376 15896 15428
rect 11428 15308 11480 15360
rect 12716 15351 12768 15360
rect 12716 15317 12725 15351
rect 12725 15317 12759 15351
rect 12759 15317 12768 15351
rect 12716 15308 12768 15317
rect 14924 15351 14976 15360
rect 14924 15317 14933 15351
rect 14933 15317 14967 15351
rect 14967 15317 14976 15351
rect 14924 15308 14976 15317
rect 15200 15308 15252 15360
rect 16396 15512 16448 15564
rect 17684 15555 17736 15564
rect 17684 15521 17693 15555
rect 17693 15521 17727 15555
rect 17727 15521 17736 15555
rect 17684 15512 17736 15521
rect 19248 15512 19300 15564
rect 19432 15623 19484 15632
rect 19432 15589 19441 15623
rect 19441 15589 19475 15623
rect 19475 15589 19484 15623
rect 19432 15580 19484 15589
rect 21824 15691 21876 15700
rect 21824 15657 21833 15691
rect 21833 15657 21867 15691
rect 21867 15657 21876 15691
rect 21824 15648 21876 15657
rect 17776 15444 17828 15496
rect 22652 15512 22704 15564
rect 16856 15376 16908 15428
rect 16672 15308 16724 15360
rect 20168 15444 20220 15496
rect 22100 15444 22152 15496
rect 22284 15487 22336 15496
rect 22284 15453 22293 15487
rect 22293 15453 22327 15487
rect 22327 15453 22336 15487
rect 22284 15444 22336 15453
rect 20720 15376 20772 15428
rect 21640 15376 21692 15428
rect 21272 15308 21324 15360
rect 22468 15308 22520 15360
rect 6630 15206 6682 15258
rect 6694 15206 6746 15258
rect 6758 15206 6810 15258
rect 6822 15206 6874 15258
rect 6886 15206 6938 15258
rect 12311 15206 12363 15258
rect 12375 15206 12427 15258
rect 12439 15206 12491 15258
rect 12503 15206 12555 15258
rect 12567 15206 12619 15258
rect 17992 15206 18044 15258
rect 18056 15206 18108 15258
rect 18120 15206 18172 15258
rect 18184 15206 18236 15258
rect 18248 15206 18300 15258
rect 23673 15206 23725 15258
rect 23737 15206 23789 15258
rect 23801 15206 23853 15258
rect 23865 15206 23917 15258
rect 23929 15206 23981 15258
rect 2964 15104 3016 15156
rect 2504 15036 2556 15088
rect 5448 15036 5500 15088
rect 7012 15036 7064 15088
rect 13544 15079 13596 15088
rect 13544 15045 13553 15079
rect 13553 15045 13587 15079
rect 13587 15045 13596 15079
rect 13544 15036 13596 15045
rect 14556 15079 14608 15088
rect 14556 15045 14565 15079
rect 14565 15045 14599 15079
rect 14599 15045 14608 15079
rect 14556 15036 14608 15045
rect 14924 15104 14976 15156
rect 15844 15104 15896 15156
rect 17316 15104 17368 15156
rect 17500 15104 17552 15156
rect 17684 15104 17736 15156
rect 18788 15104 18840 15156
rect 17868 15036 17920 15088
rect 19708 15104 19760 15156
rect 21180 15104 21232 15156
rect 1860 15011 1912 15020
rect 1860 14977 1869 15011
rect 1869 14977 1903 15011
rect 1903 14977 1912 15011
rect 1860 14968 1912 14977
rect 2044 15011 2096 15020
rect 2044 14977 2053 15011
rect 2053 14977 2087 15011
rect 2087 14977 2096 15011
rect 2044 14968 2096 14977
rect 2228 15011 2280 15020
rect 2228 14977 2237 15011
rect 2237 14977 2271 15011
rect 2271 14977 2280 15011
rect 2228 14968 2280 14977
rect 6000 14968 6052 15020
rect 7380 14968 7432 15020
rect 9128 15011 9180 15020
rect 9128 14977 9137 15011
rect 9137 14977 9171 15011
rect 9171 14977 9180 15011
rect 9128 14968 9180 14977
rect 11060 14968 11112 15020
rect 12900 15011 12952 15020
rect 12900 14977 12909 15011
rect 12909 14977 12943 15011
rect 12943 14977 12952 15011
rect 12900 14968 12952 14977
rect 14096 14968 14148 15020
rect 14280 15011 14332 15020
rect 14280 14977 14289 15011
rect 14289 14977 14323 15011
rect 14323 14977 14332 15011
rect 14280 14968 14332 14977
rect 14464 15011 14516 15020
rect 14464 14977 14473 15011
rect 14473 14977 14507 15011
rect 14507 14977 14516 15011
rect 14464 14968 14516 14977
rect 14648 15011 14700 15020
rect 14648 14977 14657 15011
rect 14657 14977 14691 15011
rect 14691 14977 14700 15011
rect 14648 14968 14700 14977
rect 15660 14968 15712 15020
rect 15936 15011 15988 15020
rect 15936 14977 15945 15011
rect 15945 14977 15979 15011
rect 15979 14977 15988 15011
rect 15936 14968 15988 14977
rect 16028 15011 16080 15020
rect 16028 14977 16037 15011
rect 16037 14977 16071 15011
rect 16071 14977 16080 15011
rect 16028 14968 16080 14977
rect 3056 14943 3108 14952
rect 3056 14909 3065 14943
rect 3065 14909 3099 14943
rect 3099 14909 3108 14943
rect 3056 14900 3108 14909
rect 6092 14900 6144 14952
rect 12072 14943 12124 14952
rect 12072 14909 12081 14943
rect 12081 14909 12115 14943
rect 12115 14909 12124 14943
rect 12072 14900 12124 14909
rect 12716 14900 12768 14952
rect 15200 14900 15252 14952
rect 16304 15011 16356 15020
rect 16304 14977 16313 15011
rect 16313 14977 16347 15011
rect 16347 14977 16356 15011
rect 16304 14968 16356 14977
rect 16672 14968 16724 15020
rect 17040 14943 17092 14952
rect 17040 14909 17049 14943
rect 17049 14909 17083 14943
rect 17083 14909 17092 14943
rect 17040 14900 17092 14909
rect 17224 15011 17276 15020
rect 17224 14977 17233 15011
rect 17233 14977 17267 15011
rect 17267 14977 17276 15011
rect 17224 14968 17276 14977
rect 17776 14900 17828 14952
rect 18788 14968 18840 15020
rect 20444 15036 20496 15088
rect 22560 15147 22612 15156
rect 22560 15113 22569 15147
rect 22569 15113 22603 15147
rect 22603 15113 22612 15147
rect 22560 15104 22612 15113
rect 18696 14900 18748 14952
rect 5908 14832 5960 14884
rect 6644 14832 6696 14884
rect 14556 14832 14608 14884
rect 5356 14764 5408 14816
rect 6552 14807 6604 14816
rect 6552 14773 6561 14807
rect 6561 14773 6595 14807
rect 6595 14773 6604 14807
rect 6552 14764 6604 14773
rect 10876 14764 10928 14816
rect 14740 14764 14792 14816
rect 15936 14832 15988 14884
rect 16856 14832 16908 14884
rect 19432 15011 19484 15020
rect 19432 14977 19441 15011
rect 19441 14977 19475 15011
rect 19475 14977 19484 15011
rect 19432 14968 19484 14977
rect 21732 14968 21784 15020
rect 20076 14900 20128 14952
rect 20536 14900 20588 14952
rect 22008 14943 22060 14952
rect 22008 14909 22017 14943
rect 22017 14909 22051 14943
rect 22051 14909 22060 14943
rect 22008 14900 22060 14909
rect 21548 14832 21600 14884
rect 21180 14764 21232 14816
rect 3790 14662 3842 14714
rect 3854 14662 3906 14714
rect 3918 14662 3970 14714
rect 3982 14662 4034 14714
rect 4046 14662 4098 14714
rect 9471 14662 9523 14714
rect 9535 14662 9587 14714
rect 9599 14662 9651 14714
rect 9663 14662 9715 14714
rect 9727 14662 9779 14714
rect 15152 14662 15204 14714
rect 15216 14662 15268 14714
rect 15280 14662 15332 14714
rect 15344 14662 15396 14714
rect 15408 14662 15460 14714
rect 20833 14662 20885 14714
rect 20897 14662 20949 14714
rect 20961 14662 21013 14714
rect 21025 14662 21077 14714
rect 21089 14662 21141 14714
rect 2320 14603 2372 14612
rect 2320 14569 2329 14603
rect 2329 14569 2363 14603
rect 2363 14569 2372 14603
rect 2320 14560 2372 14569
rect 3332 14560 3384 14612
rect 6092 14603 6144 14612
rect 6092 14569 6101 14603
rect 6101 14569 6135 14603
rect 6135 14569 6144 14603
rect 6092 14560 6144 14569
rect 7748 14560 7800 14612
rect 9220 14560 9272 14612
rect 8208 14492 8260 14544
rect 1860 14356 1912 14408
rect 2228 14356 2280 14408
rect 2872 14356 2924 14408
rect 5172 14424 5224 14476
rect 8668 14492 8720 14544
rect 1952 14331 2004 14340
rect 1952 14297 1961 14331
rect 1961 14297 1995 14331
rect 1995 14297 2004 14331
rect 1952 14288 2004 14297
rect 1676 14220 1728 14272
rect 2688 14288 2740 14340
rect 2228 14220 2280 14272
rect 3976 14263 4028 14272
rect 3976 14229 3985 14263
rect 3985 14229 4019 14263
rect 4019 14229 4028 14263
rect 3976 14220 4028 14229
rect 4344 14331 4396 14340
rect 4344 14297 4353 14331
rect 4353 14297 4387 14331
rect 4387 14297 4396 14331
rect 4344 14288 4396 14297
rect 5356 14399 5408 14408
rect 5356 14365 5365 14399
rect 5365 14365 5399 14399
rect 5399 14365 5408 14399
rect 5356 14356 5408 14365
rect 5816 14356 5868 14408
rect 6644 14399 6696 14408
rect 6644 14365 6653 14399
rect 6653 14365 6687 14399
rect 6687 14365 6696 14399
rect 6644 14356 6696 14365
rect 7288 14356 7340 14408
rect 4528 14220 4580 14272
rect 5448 14331 5500 14340
rect 5448 14297 5457 14331
rect 5457 14297 5491 14331
rect 5491 14297 5500 14331
rect 5448 14288 5500 14297
rect 6368 14331 6420 14340
rect 6368 14297 6377 14331
rect 6377 14297 6411 14331
rect 6411 14297 6420 14331
rect 6368 14288 6420 14297
rect 6460 14331 6512 14340
rect 6460 14297 6469 14331
rect 6469 14297 6503 14331
rect 6503 14297 6512 14331
rect 6460 14288 6512 14297
rect 7564 14288 7616 14340
rect 7840 14399 7892 14408
rect 7840 14365 7849 14399
rect 7849 14365 7883 14399
rect 7883 14365 7892 14399
rect 7840 14356 7892 14365
rect 8024 14356 8076 14408
rect 10784 14492 10836 14544
rect 10140 14356 10192 14408
rect 11612 14560 11664 14612
rect 13268 14560 13320 14612
rect 14280 14492 14332 14544
rect 11888 14424 11940 14476
rect 13636 14424 13688 14476
rect 14648 14560 14700 14612
rect 15476 14560 15528 14612
rect 15844 14560 15896 14612
rect 16120 14560 16172 14612
rect 19984 14560 20036 14612
rect 18880 14492 18932 14544
rect 21824 14560 21876 14612
rect 22192 14560 22244 14612
rect 20444 14492 20496 14544
rect 11704 14399 11756 14408
rect 11704 14365 11713 14399
rect 11713 14365 11747 14399
rect 11747 14365 11756 14399
rect 11704 14356 11756 14365
rect 11796 14356 11848 14408
rect 14096 14356 14148 14408
rect 14740 14399 14792 14408
rect 14740 14365 14749 14399
rect 14749 14365 14783 14399
rect 14783 14365 14792 14399
rect 14740 14356 14792 14365
rect 16304 14424 16356 14476
rect 17132 14424 17184 14476
rect 16856 14356 16908 14408
rect 19064 14424 19116 14476
rect 20720 14492 20772 14544
rect 7104 14220 7156 14272
rect 8484 14288 8536 14340
rect 8668 14220 8720 14272
rect 9220 14220 9272 14272
rect 10876 14331 10928 14340
rect 10876 14297 10885 14331
rect 10885 14297 10919 14331
rect 10919 14297 10928 14331
rect 10876 14288 10928 14297
rect 11152 14288 11204 14340
rect 13912 14288 13964 14340
rect 15108 14288 15160 14340
rect 15568 14288 15620 14340
rect 19892 14399 19944 14408
rect 19892 14365 19901 14399
rect 19901 14365 19935 14399
rect 19935 14365 19944 14399
rect 19892 14356 19944 14365
rect 13820 14220 13872 14272
rect 14556 14220 14608 14272
rect 15936 14220 15988 14272
rect 18696 14220 18748 14272
rect 19340 14220 19392 14272
rect 19616 14220 19668 14272
rect 20444 14288 20496 14340
rect 20996 14424 21048 14476
rect 21640 14399 21692 14408
rect 21640 14365 21649 14399
rect 21649 14365 21683 14399
rect 21683 14365 21692 14399
rect 21640 14356 21692 14365
rect 22008 14399 22060 14408
rect 22008 14365 22017 14399
rect 22017 14365 22051 14399
rect 22051 14365 22060 14399
rect 22008 14356 22060 14365
rect 22284 14356 22336 14408
rect 23204 14356 23256 14408
rect 20904 14263 20956 14272
rect 20904 14229 20913 14263
rect 20913 14229 20947 14263
rect 20947 14229 20956 14263
rect 20904 14220 20956 14229
rect 21456 14288 21508 14340
rect 22836 14263 22888 14272
rect 22836 14229 22845 14263
rect 22845 14229 22879 14263
rect 22879 14229 22888 14263
rect 22836 14220 22888 14229
rect 6630 14118 6682 14170
rect 6694 14118 6746 14170
rect 6758 14118 6810 14170
rect 6822 14118 6874 14170
rect 6886 14118 6938 14170
rect 12311 14118 12363 14170
rect 12375 14118 12427 14170
rect 12439 14118 12491 14170
rect 12503 14118 12555 14170
rect 12567 14118 12619 14170
rect 17992 14118 18044 14170
rect 18056 14118 18108 14170
rect 18120 14118 18172 14170
rect 18184 14118 18236 14170
rect 18248 14118 18300 14170
rect 23673 14118 23725 14170
rect 23737 14118 23789 14170
rect 23801 14118 23853 14170
rect 23865 14118 23917 14170
rect 23929 14118 23981 14170
rect 2044 14016 2096 14068
rect 2872 14059 2924 14068
rect 2872 14025 2881 14059
rect 2881 14025 2915 14059
rect 2915 14025 2924 14059
rect 2872 14016 2924 14025
rect 4436 14016 4488 14068
rect 4804 14016 4856 14068
rect 5264 14059 5316 14068
rect 5264 14025 5273 14059
rect 5273 14025 5307 14059
rect 5307 14025 5316 14059
rect 5264 14016 5316 14025
rect 6460 14016 6512 14068
rect 7564 14016 7616 14068
rect 8208 14059 8260 14068
rect 8208 14025 8217 14059
rect 8217 14025 8251 14059
rect 8251 14025 8260 14059
rect 8208 14016 8260 14025
rect 11796 14059 11848 14068
rect 11796 14025 11805 14059
rect 11805 14025 11839 14059
rect 11839 14025 11848 14059
rect 11796 14016 11848 14025
rect 12532 14016 12584 14068
rect 13268 14016 13320 14068
rect 14188 14016 14240 14068
rect 16396 14016 16448 14068
rect 16488 14016 16540 14068
rect 3056 13948 3108 14000
rect 2412 13923 2464 13932
rect 2412 13889 2421 13923
rect 2421 13889 2455 13923
rect 2455 13889 2464 13923
rect 2412 13880 2464 13889
rect 3976 13923 4028 13932
rect 5816 13948 5868 14000
rect 7380 13948 7432 14000
rect 7748 13948 7800 14000
rect 3976 13889 3994 13923
rect 3994 13889 4028 13923
rect 3976 13880 4028 13889
rect 8300 13923 8352 13932
rect 8300 13889 8309 13923
rect 8309 13889 8343 13923
rect 8343 13889 8352 13923
rect 8300 13880 8352 13889
rect 13084 13948 13136 14000
rect 11704 13923 11756 13932
rect 11704 13889 11713 13923
rect 11713 13889 11747 13923
rect 11747 13889 11756 13923
rect 11704 13880 11756 13889
rect 11888 13923 11940 13932
rect 11888 13889 11897 13923
rect 11897 13889 11931 13923
rect 11931 13889 11940 13923
rect 11888 13880 11940 13889
rect 14096 13880 14148 13932
rect 14832 13948 14884 14000
rect 14924 13880 14976 13932
rect 15108 13880 15160 13932
rect 16212 13880 16264 13932
rect 2136 13855 2188 13864
rect 2136 13821 2145 13855
rect 2145 13821 2179 13855
rect 2179 13821 2188 13855
rect 2136 13812 2188 13821
rect 4620 13744 4672 13796
rect 5540 13744 5592 13796
rect 11152 13855 11204 13864
rect 11152 13821 11161 13855
rect 11161 13821 11195 13855
rect 11195 13821 11204 13855
rect 11152 13812 11204 13821
rect 12072 13812 12124 13864
rect 13912 13855 13964 13864
rect 13912 13821 13921 13855
rect 13921 13821 13955 13855
rect 13955 13821 13964 13855
rect 13912 13812 13964 13821
rect 14280 13855 14332 13864
rect 14280 13821 14289 13855
rect 14289 13821 14323 13855
rect 14323 13821 14332 13855
rect 15016 13855 15068 13864
rect 14280 13812 14332 13821
rect 15016 13821 15025 13855
rect 15025 13821 15059 13855
rect 15059 13821 15068 13855
rect 15016 13812 15068 13821
rect 15476 13812 15528 13864
rect 17132 13923 17184 13932
rect 17132 13889 17141 13923
rect 17141 13889 17175 13923
rect 17175 13889 17184 13923
rect 17132 13880 17184 13889
rect 20260 14016 20312 14068
rect 20536 14016 20588 14068
rect 21824 14016 21876 14068
rect 19800 13923 19852 13932
rect 19800 13889 19809 13923
rect 19809 13889 19843 13923
rect 19843 13889 19852 13923
rect 19800 13880 19852 13889
rect 19984 13923 20036 13932
rect 19984 13889 19993 13923
rect 19993 13889 20027 13923
rect 20027 13889 20036 13923
rect 19984 13880 20036 13889
rect 20076 13923 20128 13932
rect 20076 13889 20085 13923
rect 20085 13889 20119 13923
rect 20119 13889 20128 13923
rect 20076 13880 20128 13889
rect 21180 13880 21232 13932
rect 7104 13787 7156 13796
rect 7104 13753 7113 13787
rect 7113 13753 7147 13787
rect 7147 13753 7156 13787
rect 7104 13744 7156 13753
rect 11520 13744 11572 13796
rect 11704 13744 11756 13796
rect 16856 13787 16908 13796
rect 16856 13753 16865 13787
rect 16865 13753 16899 13787
rect 16899 13753 16908 13787
rect 16856 13744 16908 13753
rect 19248 13812 19300 13864
rect 18420 13744 18472 13796
rect 18604 13744 18656 13796
rect 20904 13744 20956 13796
rect 20996 13744 21048 13796
rect 21272 13744 21324 13796
rect 2780 13676 2832 13728
rect 5908 13676 5960 13728
rect 6460 13676 6512 13728
rect 21916 13676 21968 13728
rect 22100 13744 22152 13796
rect 22192 13676 22244 13728
rect 22376 13719 22428 13728
rect 22376 13685 22385 13719
rect 22385 13685 22419 13719
rect 22419 13685 22428 13719
rect 22376 13676 22428 13685
rect 22744 13719 22796 13728
rect 22744 13685 22753 13719
rect 22753 13685 22787 13719
rect 22787 13685 22796 13719
rect 22744 13676 22796 13685
rect 3790 13574 3842 13626
rect 3854 13574 3906 13626
rect 3918 13574 3970 13626
rect 3982 13574 4034 13626
rect 4046 13574 4098 13626
rect 9471 13574 9523 13626
rect 9535 13574 9587 13626
rect 9599 13574 9651 13626
rect 9663 13574 9715 13626
rect 9727 13574 9779 13626
rect 15152 13574 15204 13626
rect 15216 13574 15268 13626
rect 15280 13574 15332 13626
rect 15344 13574 15396 13626
rect 15408 13574 15460 13626
rect 20833 13574 20885 13626
rect 20897 13574 20949 13626
rect 20961 13574 21013 13626
rect 21025 13574 21077 13626
rect 21089 13574 21141 13626
rect 5448 13472 5500 13524
rect 5908 13472 5960 13524
rect 7012 13472 7064 13524
rect 9220 13472 9272 13524
rect 12808 13515 12860 13524
rect 12808 13481 12817 13515
rect 12817 13481 12851 13515
rect 12851 13481 12860 13515
rect 12808 13472 12860 13481
rect 13176 13472 13228 13524
rect 13636 13472 13688 13524
rect 14188 13472 14240 13524
rect 14648 13472 14700 13524
rect 14832 13515 14884 13524
rect 14832 13481 14841 13515
rect 14841 13481 14875 13515
rect 14875 13481 14884 13515
rect 14832 13472 14884 13481
rect 14924 13472 14976 13524
rect 15384 13472 15436 13524
rect 16028 13472 16080 13524
rect 17040 13472 17092 13524
rect 19248 13472 19300 13524
rect 22928 13515 22980 13524
rect 2228 13404 2280 13456
rect 3700 13404 3752 13456
rect 4804 13404 4856 13456
rect 2136 13336 2188 13388
rect 7932 13404 7984 13456
rect 14740 13404 14792 13456
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 2320 13268 2372 13320
rect 2412 13268 2464 13320
rect 3240 13311 3292 13320
rect 3240 13277 3249 13311
rect 3249 13277 3283 13311
rect 3283 13277 3292 13311
rect 3240 13268 3292 13277
rect 7656 13336 7708 13388
rect 1860 13200 1912 13252
rect 4252 13311 4304 13320
rect 4252 13277 4261 13311
rect 4261 13277 4295 13311
rect 4295 13277 4304 13311
rect 4252 13268 4304 13277
rect 4896 13268 4948 13320
rect 5540 13268 5592 13320
rect 6552 13268 6604 13320
rect 7012 13268 7064 13320
rect 1768 13175 1820 13184
rect 1768 13141 1777 13175
rect 1777 13141 1811 13175
rect 1811 13141 1820 13175
rect 1768 13132 1820 13141
rect 2044 13132 2096 13184
rect 3424 13175 3476 13184
rect 3424 13141 3433 13175
rect 3433 13141 3467 13175
rect 3467 13141 3476 13175
rect 3424 13132 3476 13141
rect 5172 13132 5224 13184
rect 5816 13132 5868 13184
rect 6092 13175 6144 13184
rect 6092 13141 6119 13175
rect 6119 13141 6144 13175
rect 6092 13132 6144 13141
rect 7288 13200 7340 13252
rect 8208 13311 8260 13320
rect 8208 13277 8217 13311
rect 8217 13277 8251 13311
rect 8251 13277 8260 13311
rect 8208 13268 8260 13277
rect 7932 13200 7984 13252
rect 8852 13268 8904 13320
rect 10692 13311 10744 13320
rect 12900 13336 12952 13388
rect 13820 13336 13872 13388
rect 17132 13336 17184 13388
rect 17408 13336 17460 13388
rect 19524 13404 19576 13456
rect 19616 13404 19668 13456
rect 10692 13277 10731 13311
rect 10731 13277 10744 13311
rect 10692 13268 10744 13277
rect 11336 13311 11388 13320
rect 11336 13277 11345 13311
rect 11345 13277 11379 13311
rect 11379 13277 11388 13311
rect 11336 13268 11388 13277
rect 11060 13200 11112 13252
rect 11152 13200 11204 13252
rect 11704 13268 11756 13320
rect 12164 13268 12216 13320
rect 12532 13311 12584 13320
rect 12532 13277 12541 13311
rect 12541 13277 12575 13311
rect 12575 13277 12584 13311
rect 12532 13268 12584 13277
rect 13176 13268 13228 13320
rect 14004 13268 14056 13320
rect 15292 13268 15344 13320
rect 15568 13268 15620 13320
rect 16396 13311 16448 13320
rect 16396 13277 16405 13311
rect 16405 13277 16439 13311
rect 16439 13277 16448 13311
rect 16396 13268 16448 13277
rect 16580 13268 16632 13320
rect 16672 13311 16724 13320
rect 16672 13277 16681 13311
rect 16681 13277 16715 13311
rect 16715 13277 16724 13311
rect 16672 13268 16724 13277
rect 13544 13200 13596 13252
rect 10048 13132 10100 13184
rect 10508 13175 10560 13184
rect 10508 13141 10517 13175
rect 10517 13141 10551 13175
rect 10551 13141 10560 13175
rect 10508 13132 10560 13141
rect 11336 13132 11388 13184
rect 11980 13132 12032 13184
rect 14464 13243 14516 13252
rect 14464 13209 14473 13243
rect 14473 13209 14507 13243
rect 14507 13209 14516 13243
rect 14464 13200 14516 13209
rect 14924 13200 14976 13252
rect 14648 13175 14700 13184
rect 14648 13141 14657 13175
rect 14657 13141 14691 13175
rect 14691 13141 14700 13175
rect 14648 13132 14700 13141
rect 14832 13132 14884 13184
rect 15752 13132 15804 13184
rect 16212 13132 16264 13184
rect 17408 13200 17460 13252
rect 19340 13336 19392 13388
rect 18788 13268 18840 13320
rect 20812 13336 20864 13388
rect 21824 13336 21876 13388
rect 20720 13268 20772 13320
rect 22928 13481 22937 13515
rect 22937 13481 22971 13515
rect 22971 13481 22980 13515
rect 22928 13472 22980 13481
rect 19248 13200 19300 13252
rect 22836 13268 22888 13320
rect 20352 13132 20404 13184
rect 6630 13030 6682 13082
rect 6694 13030 6746 13082
rect 6758 13030 6810 13082
rect 6822 13030 6874 13082
rect 6886 13030 6938 13082
rect 12311 13030 12363 13082
rect 12375 13030 12427 13082
rect 12439 13030 12491 13082
rect 12503 13030 12555 13082
rect 12567 13030 12619 13082
rect 17992 13030 18044 13082
rect 18056 13030 18108 13082
rect 18120 13030 18172 13082
rect 18184 13030 18236 13082
rect 18248 13030 18300 13082
rect 23673 13030 23725 13082
rect 23737 13030 23789 13082
rect 23801 13030 23853 13082
rect 23865 13030 23917 13082
rect 23929 13030 23981 13082
rect 2596 12928 2648 12980
rect 2412 12860 2464 12912
rect 6092 12928 6144 12980
rect 10508 12928 10560 12980
rect 13176 12928 13228 12980
rect 13912 12971 13964 12980
rect 13912 12937 13921 12971
rect 13921 12937 13955 12971
rect 13955 12937 13964 12971
rect 13912 12928 13964 12937
rect 14372 12928 14424 12980
rect 17132 12928 17184 12980
rect 17592 12928 17644 12980
rect 18512 12928 18564 12980
rect 20076 12928 20128 12980
rect 5172 12903 5224 12912
rect 5172 12869 5181 12903
rect 5181 12869 5215 12903
rect 5215 12869 5224 12903
rect 5172 12860 5224 12869
rect 6920 12860 6972 12912
rect 7104 12860 7156 12912
rect 8852 12860 8904 12912
rect 2688 12792 2740 12844
rect 2964 12835 3016 12844
rect 2964 12801 2973 12835
rect 2973 12801 3007 12835
rect 3007 12801 3016 12835
rect 2964 12792 3016 12801
rect 3240 12792 3292 12844
rect 3424 12792 3476 12844
rect 5540 12792 5592 12844
rect 6092 12792 6144 12844
rect 6460 12792 6512 12844
rect 3148 12724 3200 12776
rect 5448 12724 5500 12776
rect 9036 12835 9088 12844
rect 9036 12801 9045 12835
rect 9045 12801 9079 12835
rect 9079 12801 9088 12835
rect 9036 12792 9088 12801
rect 9220 12835 9272 12844
rect 9220 12801 9229 12835
rect 9229 12801 9263 12835
rect 9263 12801 9272 12835
rect 9220 12792 9272 12801
rect 9956 12792 10008 12844
rect 10232 12835 10284 12844
rect 10232 12801 10241 12835
rect 10241 12801 10275 12835
rect 10275 12801 10284 12835
rect 10232 12792 10284 12801
rect 10692 12860 10744 12912
rect 11704 12903 11756 12912
rect 11704 12869 11713 12903
rect 11713 12869 11747 12903
rect 11747 12869 11756 12903
rect 11704 12860 11756 12869
rect 12716 12903 12768 12912
rect 12716 12869 12725 12903
rect 12725 12869 12759 12903
rect 12759 12869 12768 12903
rect 12716 12860 12768 12869
rect 13728 12860 13780 12912
rect 11980 12835 12032 12844
rect 11980 12801 11989 12835
rect 11989 12801 12023 12835
rect 12023 12801 12032 12835
rect 11980 12792 12032 12801
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 10692 12724 10744 12776
rect 14188 12835 14240 12844
rect 14188 12801 14197 12835
rect 14197 12801 14231 12835
rect 14231 12801 14240 12835
rect 14188 12792 14240 12801
rect 15384 12860 15436 12912
rect 15476 12903 15528 12912
rect 15476 12869 15485 12903
rect 15485 12869 15519 12903
rect 15519 12869 15528 12903
rect 15476 12860 15528 12869
rect 14832 12792 14884 12844
rect 14464 12724 14516 12776
rect 15292 12792 15344 12844
rect 16028 12860 16080 12912
rect 16304 12860 16356 12912
rect 15752 12792 15804 12844
rect 21824 12860 21876 12912
rect 16948 12835 17000 12844
rect 16948 12801 16958 12835
rect 16958 12801 16992 12835
rect 16992 12801 17000 12835
rect 16948 12792 17000 12801
rect 17132 12835 17184 12844
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 17224 12835 17276 12844
rect 17224 12801 17233 12835
rect 17233 12801 17267 12835
rect 17267 12801 17276 12835
rect 17224 12792 17276 12801
rect 17408 12792 17460 12844
rect 19064 12792 19116 12844
rect 21640 12792 21692 12844
rect 22100 12792 22152 12844
rect 22468 12835 22520 12844
rect 22468 12801 22477 12835
rect 22477 12801 22511 12835
rect 22511 12801 22520 12835
rect 22468 12792 22520 12801
rect 18236 12724 18288 12776
rect 18512 12767 18564 12776
rect 18512 12733 18521 12767
rect 18521 12733 18555 12767
rect 18555 12733 18564 12767
rect 18512 12724 18564 12733
rect 18788 12767 18840 12776
rect 18788 12733 18797 12767
rect 18797 12733 18831 12767
rect 18831 12733 18840 12767
rect 18788 12724 18840 12733
rect 2780 12699 2832 12708
rect 2780 12665 2789 12699
rect 2789 12665 2823 12699
rect 2823 12665 2832 12699
rect 2780 12656 2832 12665
rect 3056 12656 3108 12708
rect 3424 12656 3476 12708
rect 2044 12588 2096 12640
rect 2504 12588 2556 12640
rect 2596 12588 2648 12640
rect 2964 12588 3016 12640
rect 5264 12588 5316 12640
rect 6000 12656 6052 12708
rect 6460 12656 6512 12708
rect 8024 12656 8076 12708
rect 11888 12656 11940 12708
rect 9312 12631 9364 12640
rect 9312 12597 9321 12631
rect 9321 12597 9355 12631
rect 9355 12597 9364 12631
rect 9312 12588 9364 12597
rect 11152 12588 11204 12640
rect 13452 12656 13504 12708
rect 13268 12588 13320 12640
rect 15476 12588 15528 12640
rect 17040 12656 17092 12708
rect 18604 12656 18656 12708
rect 19156 12656 19208 12708
rect 16580 12588 16632 12640
rect 17868 12588 17920 12640
rect 20352 12588 20404 12640
rect 22928 12631 22980 12640
rect 22928 12597 22937 12631
rect 22937 12597 22971 12631
rect 22971 12597 22980 12631
rect 22928 12588 22980 12597
rect 3790 12486 3842 12538
rect 3854 12486 3906 12538
rect 3918 12486 3970 12538
rect 3982 12486 4034 12538
rect 4046 12486 4098 12538
rect 9471 12486 9523 12538
rect 9535 12486 9587 12538
rect 9599 12486 9651 12538
rect 9663 12486 9715 12538
rect 9727 12486 9779 12538
rect 15152 12486 15204 12538
rect 15216 12486 15268 12538
rect 15280 12486 15332 12538
rect 15344 12486 15396 12538
rect 15408 12486 15460 12538
rect 20833 12486 20885 12538
rect 20897 12486 20949 12538
rect 20961 12486 21013 12538
rect 21025 12486 21077 12538
rect 21089 12486 21141 12538
rect 1768 12427 1820 12436
rect 1768 12393 1777 12427
rect 1777 12393 1811 12427
rect 1811 12393 1820 12427
rect 1768 12384 1820 12393
rect 1952 12384 2004 12436
rect 2412 12427 2464 12436
rect 2412 12393 2421 12427
rect 2421 12393 2455 12427
rect 2455 12393 2464 12427
rect 2412 12384 2464 12393
rect 2596 12427 2648 12436
rect 2596 12393 2605 12427
rect 2605 12393 2639 12427
rect 2639 12393 2648 12427
rect 2596 12384 2648 12393
rect 4804 12384 4856 12436
rect 5264 12384 5316 12436
rect 5632 12384 5684 12436
rect 7288 12384 7340 12436
rect 7564 12427 7616 12436
rect 7564 12393 7573 12427
rect 7573 12393 7607 12427
rect 7607 12393 7616 12427
rect 7564 12384 7616 12393
rect 8116 12427 8168 12436
rect 8116 12393 8125 12427
rect 8125 12393 8159 12427
rect 8159 12393 8168 12427
rect 8116 12384 8168 12393
rect 14648 12384 14700 12436
rect 7012 12316 7064 12368
rect 8208 12316 8260 12368
rect 1952 12291 2004 12300
rect 1952 12257 1961 12291
rect 1961 12257 1995 12291
rect 1995 12257 2004 12291
rect 1952 12248 2004 12257
rect 2136 12248 2188 12300
rect 4528 12248 4580 12300
rect 3700 12180 3752 12232
rect 4436 12180 4488 12232
rect 6920 12223 6972 12232
rect 6920 12189 6929 12223
rect 6929 12189 6963 12223
rect 6963 12189 6972 12223
rect 7380 12223 7432 12232
rect 6920 12180 6972 12189
rect 7380 12189 7389 12223
rect 7389 12189 7423 12223
rect 7423 12189 7432 12223
rect 7380 12180 7432 12189
rect 7564 12223 7616 12232
rect 7564 12189 7573 12223
rect 7573 12189 7607 12223
rect 7607 12189 7616 12223
rect 7564 12180 7616 12189
rect 7932 12180 7984 12232
rect 2780 12155 2832 12164
rect 2780 12121 2789 12155
rect 2789 12121 2823 12155
rect 2823 12121 2832 12155
rect 2780 12112 2832 12121
rect 2964 12112 3016 12164
rect 3240 12044 3292 12096
rect 3792 12044 3844 12096
rect 5448 12044 5500 12096
rect 7104 12112 7156 12164
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 9220 12316 9272 12368
rect 10324 12316 10376 12368
rect 13820 12316 13872 12368
rect 11612 12248 11664 12300
rect 12992 12248 13044 12300
rect 14556 12248 14608 12300
rect 16948 12384 17000 12436
rect 17500 12384 17552 12436
rect 18328 12384 18380 12436
rect 19340 12384 19392 12436
rect 19524 12384 19576 12436
rect 19708 12427 19760 12436
rect 19708 12393 19717 12427
rect 19717 12393 19751 12427
rect 19751 12393 19760 12427
rect 19708 12384 19760 12393
rect 21824 12384 21876 12436
rect 15200 12316 15252 12368
rect 15568 12316 15620 12368
rect 14924 12248 14976 12300
rect 15844 12316 15896 12368
rect 16672 12316 16724 12368
rect 16580 12248 16632 12300
rect 9588 12180 9640 12232
rect 9864 12180 9916 12232
rect 12072 12180 12124 12232
rect 12716 12180 12768 12232
rect 8484 12112 8536 12164
rect 10232 12112 10284 12164
rect 11888 12112 11940 12164
rect 12992 12112 13044 12164
rect 8576 12087 8628 12096
rect 8576 12053 8585 12087
rect 8585 12053 8619 12087
rect 8619 12053 8628 12087
rect 8576 12044 8628 12053
rect 9220 12087 9272 12096
rect 9220 12053 9229 12087
rect 9229 12053 9263 12087
rect 9263 12053 9272 12087
rect 9220 12044 9272 12053
rect 10508 12087 10560 12096
rect 10508 12053 10517 12087
rect 10517 12053 10551 12087
rect 10551 12053 10560 12087
rect 10508 12044 10560 12053
rect 13268 12223 13320 12232
rect 13268 12189 13277 12223
rect 13277 12189 13311 12223
rect 13311 12189 13320 12223
rect 13268 12180 13320 12189
rect 13728 12180 13780 12232
rect 14372 12180 14424 12232
rect 14464 12223 14516 12232
rect 14464 12189 14473 12223
rect 14473 12189 14507 12223
rect 14507 12189 14516 12223
rect 14464 12180 14516 12189
rect 15568 12223 15620 12232
rect 15568 12189 15577 12223
rect 15577 12189 15611 12223
rect 15611 12189 15620 12223
rect 15568 12180 15620 12189
rect 15660 12223 15712 12232
rect 15660 12189 15669 12223
rect 15669 12189 15703 12223
rect 15703 12189 15712 12223
rect 15660 12180 15712 12189
rect 15844 12223 15896 12232
rect 15844 12189 15853 12223
rect 15853 12189 15887 12223
rect 15887 12189 15896 12223
rect 15844 12180 15896 12189
rect 13544 12112 13596 12164
rect 16028 12112 16080 12164
rect 16488 12223 16540 12232
rect 16488 12189 16497 12223
rect 16497 12189 16531 12223
rect 16531 12189 16540 12223
rect 16488 12180 16540 12189
rect 16672 12223 16724 12232
rect 16672 12189 16681 12223
rect 16681 12189 16715 12223
rect 16715 12189 16724 12223
rect 16672 12180 16724 12189
rect 17040 12316 17092 12368
rect 19616 12316 19668 12368
rect 17776 12291 17828 12300
rect 17776 12257 17785 12291
rect 17785 12257 17819 12291
rect 17819 12257 17828 12291
rect 17776 12248 17828 12257
rect 17868 12291 17920 12300
rect 17868 12257 17877 12291
rect 17877 12257 17911 12291
rect 17911 12257 17920 12291
rect 17868 12248 17920 12257
rect 19340 12248 19392 12300
rect 19800 12248 19852 12300
rect 17408 12180 17460 12232
rect 19064 12112 19116 12164
rect 14280 12044 14332 12096
rect 17316 12044 17368 12096
rect 17776 12044 17828 12096
rect 20076 12223 20128 12232
rect 20076 12189 20085 12223
rect 20085 12189 20119 12223
rect 20119 12189 20128 12223
rect 20076 12180 20128 12189
rect 21088 12291 21140 12300
rect 21088 12257 21097 12291
rect 21097 12257 21131 12291
rect 21131 12257 21140 12291
rect 21088 12248 21140 12257
rect 21272 12316 21324 12368
rect 21456 12316 21508 12368
rect 21548 12316 21600 12368
rect 22468 12316 22520 12368
rect 20352 12223 20404 12232
rect 20352 12189 20361 12223
rect 20361 12189 20395 12223
rect 20395 12189 20404 12223
rect 20352 12180 20404 12189
rect 20720 12180 20772 12232
rect 21180 12180 21232 12232
rect 21456 12223 21508 12232
rect 21456 12189 21465 12223
rect 21465 12189 21499 12223
rect 21499 12189 21508 12223
rect 21456 12180 21508 12189
rect 21916 12248 21968 12300
rect 22928 12248 22980 12300
rect 20536 12044 20588 12096
rect 22008 12112 22060 12164
rect 22744 12180 22796 12232
rect 23020 12223 23072 12232
rect 23020 12189 23029 12223
rect 23029 12189 23063 12223
rect 23063 12189 23072 12223
rect 23020 12180 23072 12189
rect 23204 12223 23256 12232
rect 23204 12189 23213 12223
rect 23213 12189 23247 12223
rect 23247 12189 23256 12223
rect 23204 12180 23256 12189
rect 22468 12112 22520 12164
rect 22652 12112 22704 12164
rect 22376 12044 22428 12096
rect 6630 11942 6682 11994
rect 6694 11942 6746 11994
rect 6758 11942 6810 11994
rect 6822 11942 6874 11994
rect 6886 11942 6938 11994
rect 12311 11942 12363 11994
rect 12375 11942 12427 11994
rect 12439 11942 12491 11994
rect 12503 11942 12555 11994
rect 12567 11942 12619 11994
rect 17992 11942 18044 11994
rect 18056 11942 18108 11994
rect 18120 11942 18172 11994
rect 18184 11942 18236 11994
rect 18248 11942 18300 11994
rect 23673 11942 23725 11994
rect 23737 11942 23789 11994
rect 23801 11942 23853 11994
rect 23865 11942 23917 11994
rect 23929 11942 23981 11994
rect 4344 11883 4396 11892
rect 4344 11849 4353 11883
rect 4353 11849 4387 11883
rect 4387 11849 4396 11883
rect 4344 11840 4396 11849
rect 4804 11840 4856 11892
rect 5080 11840 5132 11892
rect 5816 11840 5868 11892
rect 6184 11840 6236 11892
rect 7196 11840 7248 11892
rect 11428 11840 11480 11892
rect 12072 11840 12124 11892
rect 13268 11840 13320 11892
rect 1860 11772 1912 11824
rect 3516 11772 3568 11824
rect 5908 11772 5960 11824
rect 6460 11772 6512 11824
rect 10508 11772 10560 11824
rect 12164 11772 12216 11824
rect 12716 11772 12768 11824
rect 13912 11815 13964 11824
rect 13912 11781 13921 11815
rect 13921 11781 13955 11815
rect 13955 11781 13964 11815
rect 13912 11772 13964 11781
rect 14096 11772 14148 11824
rect 14188 11772 14240 11824
rect 14556 11840 14608 11892
rect 15384 11840 15436 11892
rect 15936 11840 15988 11892
rect 16580 11772 16632 11824
rect 5356 11747 5408 11756
rect 5356 11713 5365 11747
rect 5365 11713 5399 11747
rect 5399 11713 5408 11747
rect 5356 11704 5408 11713
rect 5448 11747 5500 11756
rect 5448 11713 5457 11747
rect 5457 11713 5491 11747
rect 5491 11713 5500 11747
rect 5448 11704 5500 11713
rect 5540 11747 5592 11756
rect 5540 11713 5549 11747
rect 5549 11713 5583 11747
rect 5583 11713 5592 11747
rect 5540 11704 5592 11713
rect 6736 11747 6788 11756
rect 6736 11713 6745 11747
rect 6745 11713 6779 11747
rect 6779 11713 6788 11747
rect 6736 11704 6788 11713
rect 6920 11747 6972 11756
rect 6920 11713 6929 11747
rect 6929 11713 6963 11747
rect 6963 11713 6972 11747
rect 6920 11704 6972 11713
rect 2780 11636 2832 11688
rect 3700 11679 3752 11688
rect 3700 11645 3709 11679
rect 3709 11645 3743 11679
rect 3743 11645 3752 11679
rect 3700 11636 3752 11645
rect 3792 11679 3844 11688
rect 3792 11645 3801 11679
rect 3801 11645 3835 11679
rect 3835 11645 3844 11679
rect 3792 11636 3844 11645
rect 4160 11679 4212 11688
rect 4160 11645 4169 11679
rect 4169 11645 4203 11679
rect 4203 11645 4212 11679
rect 4160 11636 4212 11645
rect 5816 11679 5868 11688
rect 5816 11645 5825 11679
rect 5825 11645 5859 11679
rect 5859 11645 5868 11679
rect 5816 11636 5868 11645
rect 5908 11636 5960 11688
rect 7196 11679 7248 11688
rect 7196 11645 7205 11679
rect 7205 11645 7239 11679
rect 7239 11645 7248 11679
rect 7196 11636 7248 11645
rect 8760 11747 8812 11756
rect 8760 11713 8769 11747
rect 8769 11713 8803 11747
rect 8803 11713 8812 11747
rect 8760 11704 8812 11713
rect 8852 11747 8904 11756
rect 8852 11713 8861 11747
rect 8861 11713 8895 11747
rect 8895 11713 8904 11747
rect 8852 11704 8904 11713
rect 8944 11636 8996 11688
rect 10048 11747 10100 11756
rect 10048 11713 10057 11747
rect 10057 11713 10091 11747
rect 10091 11713 10100 11747
rect 10048 11704 10100 11713
rect 10140 11704 10192 11756
rect 12072 11704 12124 11756
rect 13820 11704 13872 11756
rect 14464 11704 14516 11756
rect 15016 11704 15068 11756
rect 15844 11704 15896 11756
rect 17316 11840 17368 11892
rect 17408 11883 17460 11892
rect 17408 11849 17417 11883
rect 17417 11849 17451 11883
rect 17451 11849 17460 11883
rect 17408 11840 17460 11849
rect 19984 11840 20036 11892
rect 22008 11840 22060 11892
rect 17040 11704 17092 11756
rect 5172 11568 5224 11620
rect 5540 11568 5592 11620
rect 6920 11568 6972 11620
rect 7288 11568 7340 11620
rect 10232 11636 10284 11688
rect 13360 11679 13412 11688
rect 13360 11645 13369 11679
rect 13369 11645 13403 11679
rect 13403 11645 13412 11679
rect 13360 11636 13412 11645
rect 14004 11636 14056 11688
rect 14280 11568 14332 11620
rect 16764 11636 16816 11688
rect 17592 11704 17644 11756
rect 20536 11704 20588 11756
rect 22560 11772 22612 11824
rect 22744 11815 22796 11824
rect 22744 11781 22753 11815
rect 22753 11781 22787 11815
rect 22787 11781 22796 11815
rect 22744 11772 22796 11781
rect 21364 11704 21416 11756
rect 17868 11679 17920 11688
rect 17868 11645 17877 11679
rect 17877 11645 17911 11679
rect 17911 11645 17920 11679
rect 17868 11636 17920 11645
rect 20168 11636 20220 11688
rect 20444 11636 20496 11688
rect 23020 11636 23072 11688
rect 16856 11568 16908 11620
rect 19800 11568 19852 11620
rect 20260 11568 20312 11620
rect 21364 11568 21416 11620
rect 3700 11500 3752 11552
rect 9128 11500 9180 11552
rect 9588 11500 9640 11552
rect 11244 11500 11296 11552
rect 11704 11500 11756 11552
rect 16212 11543 16264 11552
rect 16212 11509 16221 11543
rect 16221 11509 16255 11543
rect 16255 11509 16264 11543
rect 16212 11500 16264 11509
rect 16304 11500 16356 11552
rect 18696 11500 18748 11552
rect 19708 11500 19760 11552
rect 20444 11500 20496 11552
rect 3790 11398 3842 11450
rect 3854 11398 3906 11450
rect 3918 11398 3970 11450
rect 3982 11398 4034 11450
rect 4046 11398 4098 11450
rect 9471 11398 9523 11450
rect 9535 11398 9587 11450
rect 9599 11398 9651 11450
rect 9663 11398 9715 11450
rect 9727 11398 9779 11450
rect 15152 11398 15204 11450
rect 15216 11398 15268 11450
rect 15280 11398 15332 11450
rect 15344 11398 15396 11450
rect 15408 11398 15460 11450
rect 20833 11398 20885 11450
rect 20897 11398 20949 11450
rect 20961 11398 21013 11450
rect 21025 11398 21077 11450
rect 21089 11398 21141 11450
rect 1952 11296 2004 11348
rect 5448 11296 5500 11348
rect 7932 11296 7984 11348
rect 13084 11296 13136 11348
rect 4160 11228 4212 11280
rect 5632 11228 5684 11280
rect 6644 11228 6696 11280
rect 1584 11135 1636 11144
rect 1584 11101 1593 11135
rect 1593 11101 1627 11135
rect 1627 11101 1636 11135
rect 1584 11092 1636 11101
rect 1860 11092 1912 11144
rect 3700 11160 3752 11212
rect 4436 11160 4488 11212
rect 2780 11092 2832 11144
rect 4528 11092 4580 11144
rect 5448 11092 5500 11144
rect 6092 11092 6144 11144
rect 11612 11228 11664 11280
rect 13544 11296 13596 11348
rect 14556 11296 14608 11348
rect 14740 11296 14792 11348
rect 8944 11160 8996 11212
rect 10324 11160 10376 11212
rect 10416 11160 10468 11212
rect 14096 11160 14148 11212
rect 16488 11296 16540 11348
rect 16672 11296 16724 11348
rect 18328 11296 18380 11348
rect 20076 11339 20128 11348
rect 20076 11305 20085 11339
rect 20085 11305 20119 11339
rect 20119 11305 20128 11339
rect 20076 11296 20128 11305
rect 20352 11296 20404 11348
rect 15660 11228 15712 11280
rect 6368 11024 6420 11076
rect 9036 11092 9088 11144
rect 9404 11092 9456 11144
rect 11704 11092 11756 11144
rect 15752 11160 15804 11212
rect 16028 11160 16080 11212
rect 9864 11024 9916 11076
rect 10140 11067 10192 11076
rect 10140 11033 10149 11067
rect 10149 11033 10183 11067
rect 10183 11033 10192 11067
rect 10140 11024 10192 11033
rect 11612 11067 11664 11076
rect 11612 11033 11621 11067
rect 11621 11033 11655 11067
rect 11655 11033 11664 11067
rect 11612 11024 11664 11033
rect 11796 11067 11848 11076
rect 11796 11033 11805 11067
rect 11805 11033 11839 11067
rect 11839 11033 11848 11067
rect 11796 11024 11848 11033
rect 13268 11024 13320 11076
rect 13820 11024 13872 11076
rect 14924 11024 14976 11076
rect 15292 11135 15344 11144
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 16304 11135 16356 11144
rect 16304 11101 16313 11135
rect 16313 11101 16347 11135
rect 16347 11101 16356 11135
rect 16304 11092 16356 11101
rect 17040 11135 17092 11144
rect 17040 11101 17049 11135
rect 17049 11101 17083 11135
rect 17083 11101 17092 11135
rect 17040 11092 17092 11101
rect 17500 11160 17552 11212
rect 18512 11160 18564 11212
rect 6000 10956 6052 11008
rect 6276 10956 6328 11008
rect 11244 10956 11296 11008
rect 16212 11024 16264 11076
rect 16488 11024 16540 11076
rect 17776 11092 17828 11144
rect 22376 11228 22428 11280
rect 23204 11228 23256 11280
rect 21916 11203 21968 11212
rect 21916 11169 21925 11203
rect 21925 11169 21959 11203
rect 21959 11169 21968 11203
rect 21916 11160 21968 11169
rect 22284 11160 22336 11212
rect 16948 10956 17000 11008
rect 18420 11024 18472 11076
rect 18512 11024 18564 11076
rect 19800 11135 19852 11144
rect 19800 11101 19809 11135
rect 19809 11101 19843 11135
rect 19843 11101 19852 11135
rect 19800 11092 19852 11101
rect 21364 11092 21416 11144
rect 21732 11092 21784 11144
rect 22100 11092 22152 11144
rect 22468 11135 22520 11144
rect 22468 11101 22477 11135
rect 22477 11101 22511 11135
rect 22511 11101 22520 11135
rect 22468 11092 22520 11101
rect 22652 11135 22704 11144
rect 22652 11101 22661 11135
rect 22661 11101 22695 11135
rect 22695 11101 22704 11135
rect 22652 11092 22704 11101
rect 18788 11024 18840 11076
rect 19064 11024 19116 11076
rect 19248 10956 19300 11008
rect 19524 11067 19576 11076
rect 19524 11033 19533 11067
rect 19533 11033 19567 11067
rect 19567 11033 19576 11067
rect 19524 11024 19576 11033
rect 6630 10854 6682 10906
rect 6694 10854 6746 10906
rect 6758 10854 6810 10906
rect 6822 10854 6874 10906
rect 6886 10854 6938 10906
rect 12311 10854 12363 10906
rect 12375 10854 12427 10906
rect 12439 10854 12491 10906
rect 12503 10854 12555 10906
rect 12567 10854 12619 10906
rect 17992 10854 18044 10906
rect 18056 10854 18108 10906
rect 18120 10854 18172 10906
rect 18184 10854 18236 10906
rect 18248 10854 18300 10906
rect 23673 10854 23725 10906
rect 23737 10854 23789 10906
rect 23801 10854 23853 10906
rect 23865 10854 23917 10906
rect 23929 10854 23981 10906
rect 1584 10752 1636 10804
rect 2964 10752 3016 10804
rect 5080 10752 5132 10804
rect 5356 10752 5408 10804
rect 6552 10752 6604 10804
rect 8760 10752 8812 10804
rect 9312 10752 9364 10804
rect 11704 10752 11756 10804
rect 12716 10752 12768 10804
rect 13728 10752 13780 10804
rect 2228 10727 2280 10736
rect 2228 10693 2237 10727
rect 2237 10693 2271 10727
rect 2271 10693 2280 10727
rect 2228 10684 2280 10693
rect 2504 10684 2556 10736
rect 4436 10684 4488 10736
rect 2320 10616 2372 10668
rect 2964 10659 3016 10668
rect 2964 10625 2973 10659
rect 2973 10625 3007 10659
rect 3007 10625 3016 10659
rect 2964 10616 3016 10625
rect 3148 10616 3200 10668
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 6184 10616 6236 10668
rect 7012 10684 7064 10736
rect 7104 10659 7156 10668
rect 7104 10625 7113 10659
rect 7113 10625 7147 10659
rect 7147 10625 7156 10659
rect 7104 10616 7156 10625
rect 7656 10616 7708 10668
rect 8668 10616 8720 10668
rect 10140 10684 10192 10736
rect 9128 10659 9180 10668
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 9128 10616 9180 10625
rect 9956 10616 10008 10668
rect 10324 10616 10376 10668
rect 1676 10548 1728 10600
rect 2412 10548 2464 10600
rect 4160 10548 4212 10600
rect 5816 10591 5868 10600
rect 5816 10557 5825 10591
rect 5825 10557 5859 10591
rect 5859 10557 5868 10591
rect 5816 10548 5868 10557
rect 7012 10591 7064 10600
rect 7012 10557 7021 10591
rect 7021 10557 7055 10591
rect 7055 10557 7064 10591
rect 7012 10548 7064 10557
rect 7196 10591 7248 10600
rect 7196 10557 7205 10591
rect 7205 10557 7239 10591
rect 7239 10557 7248 10591
rect 7196 10548 7248 10557
rect 10600 10548 10652 10600
rect 7472 10480 7524 10532
rect 2596 10412 2648 10464
rect 3700 10412 3752 10464
rect 5724 10412 5776 10464
rect 10508 10412 10560 10464
rect 10600 10455 10652 10464
rect 10600 10421 10609 10455
rect 10609 10421 10643 10455
rect 10643 10421 10652 10455
rect 10600 10412 10652 10421
rect 10876 10412 10928 10464
rect 12072 10659 12124 10668
rect 12072 10625 12081 10659
rect 12081 10625 12115 10659
rect 12115 10625 12124 10659
rect 12072 10616 12124 10625
rect 12256 10659 12308 10668
rect 12256 10625 12265 10659
rect 12265 10625 12299 10659
rect 12299 10625 12308 10659
rect 12256 10616 12308 10625
rect 13268 10684 13320 10736
rect 14004 10616 14056 10668
rect 14280 10659 14332 10668
rect 14280 10625 14287 10659
rect 14287 10625 14332 10659
rect 14280 10616 14332 10625
rect 13268 10548 13320 10600
rect 15292 10752 15344 10804
rect 15568 10752 15620 10804
rect 15200 10616 15252 10668
rect 15844 10659 15896 10668
rect 15844 10625 15853 10659
rect 15853 10625 15887 10659
rect 15887 10625 15896 10659
rect 15844 10616 15896 10625
rect 17132 10752 17184 10804
rect 16580 10684 16632 10736
rect 18420 10752 18472 10804
rect 21364 10795 21416 10804
rect 21364 10761 21373 10795
rect 21373 10761 21407 10795
rect 21407 10761 21416 10795
rect 21364 10752 21416 10761
rect 16856 10659 16908 10668
rect 16856 10625 16865 10659
rect 16865 10625 16899 10659
rect 16899 10625 16908 10659
rect 16856 10616 16908 10625
rect 13176 10523 13228 10532
rect 13176 10489 13185 10523
rect 13185 10489 13219 10523
rect 13219 10489 13228 10523
rect 13176 10480 13228 10489
rect 14188 10480 14240 10532
rect 14372 10412 14424 10464
rect 15568 10412 15620 10464
rect 17316 10616 17368 10668
rect 19432 10684 19484 10736
rect 18604 10659 18656 10668
rect 18604 10625 18613 10659
rect 18613 10625 18647 10659
rect 18647 10625 18656 10659
rect 18604 10616 18656 10625
rect 18696 10616 18748 10668
rect 21180 10616 21232 10668
rect 18052 10412 18104 10464
rect 18328 10412 18380 10464
rect 19248 10412 19300 10464
rect 22100 10591 22152 10600
rect 22100 10557 22109 10591
rect 22109 10557 22143 10591
rect 22143 10557 22152 10591
rect 22100 10548 22152 10557
rect 22376 10480 22428 10532
rect 19616 10412 19668 10464
rect 20720 10412 20772 10464
rect 21732 10412 21784 10464
rect 22560 10455 22612 10464
rect 22560 10421 22569 10455
rect 22569 10421 22603 10455
rect 22603 10421 22612 10455
rect 22560 10412 22612 10421
rect 3790 10310 3842 10362
rect 3854 10310 3906 10362
rect 3918 10310 3970 10362
rect 3982 10310 4034 10362
rect 4046 10310 4098 10362
rect 9471 10310 9523 10362
rect 9535 10310 9587 10362
rect 9599 10310 9651 10362
rect 9663 10310 9715 10362
rect 9727 10310 9779 10362
rect 15152 10310 15204 10362
rect 15216 10310 15268 10362
rect 15280 10310 15332 10362
rect 15344 10310 15396 10362
rect 15408 10310 15460 10362
rect 20833 10310 20885 10362
rect 20897 10310 20949 10362
rect 20961 10310 21013 10362
rect 21025 10310 21077 10362
rect 21089 10310 21141 10362
rect 4252 10208 4304 10260
rect 5632 10208 5684 10260
rect 7380 10208 7432 10260
rect 10140 10208 10192 10260
rect 13636 10208 13688 10260
rect 17868 10208 17920 10260
rect 18052 10208 18104 10260
rect 18696 10208 18748 10260
rect 22468 10208 22520 10260
rect 2504 10140 2556 10192
rect 3240 10183 3292 10192
rect 3240 10149 3249 10183
rect 3249 10149 3283 10183
rect 3283 10149 3292 10183
rect 3240 10140 3292 10149
rect 2780 10072 2832 10124
rect 2320 9936 2372 9988
rect 2780 9868 2832 9920
rect 4436 10072 4488 10124
rect 5816 10072 5868 10124
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 4160 10047 4212 10056
rect 4160 10013 4169 10047
rect 4169 10013 4203 10047
rect 4203 10013 4212 10047
rect 4160 10004 4212 10013
rect 4620 10004 4672 10056
rect 4988 10047 5040 10056
rect 4988 10013 4997 10047
rect 4997 10013 5031 10047
rect 5031 10013 5040 10047
rect 4988 10004 5040 10013
rect 5172 10004 5224 10056
rect 6552 10072 6604 10124
rect 10876 10140 10928 10192
rect 13268 10183 13320 10192
rect 13268 10149 13277 10183
rect 13277 10149 13311 10183
rect 13311 10149 13320 10183
rect 13268 10140 13320 10149
rect 14280 10140 14332 10192
rect 9864 10072 9916 10124
rect 10048 10072 10100 10124
rect 13176 10072 13228 10124
rect 16212 10140 16264 10192
rect 17592 10140 17644 10192
rect 7104 10004 7156 10056
rect 8944 10004 8996 10056
rect 9128 10004 9180 10056
rect 11704 10047 11756 10056
rect 11704 10013 11713 10047
rect 11713 10013 11747 10047
rect 11747 10013 11756 10047
rect 11704 10004 11756 10013
rect 11980 10047 12032 10056
rect 11980 10013 11989 10047
rect 11989 10013 12023 10047
rect 12023 10013 12032 10047
rect 11980 10004 12032 10013
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 14372 10047 14424 10056
rect 14372 10013 14381 10047
rect 14381 10013 14415 10047
rect 14415 10013 14424 10047
rect 14372 10004 14424 10013
rect 15108 10004 15160 10056
rect 15476 10004 15528 10056
rect 7564 9936 7616 9988
rect 11796 9936 11848 9988
rect 14832 9936 14884 9988
rect 15568 9936 15620 9988
rect 16212 9936 16264 9988
rect 19156 10072 19208 10124
rect 20812 10072 20864 10124
rect 16580 10047 16632 10056
rect 16580 10013 16589 10047
rect 16589 10013 16623 10047
rect 16623 10013 16632 10047
rect 16580 10004 16632 10013
rect 16856 10004 16908 10056
rect 16948 9979 17000 9988
rect 16948 9945 16957 9979
rect 16957 9945 16991 9979
rect 16991 9945 17000 9979
rect 16948 9936 17000 9945
rect 18328 10047 18380 10056
rect 18328 10013 18337 10047
rect 18337 10013 18371 10047
rect 18371 10013 18380 10047
rect 18328 10004 18380 10013
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 18512 10047 18564 10056
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 18512 10004 18564 10013
rect 19432 10004 19484 10056
rect 20260 10004 20312 10056
rect 20628 10004 20680 10056
rect 21088 10004 21140 10056
rect 21364 10047 21416 10056
rect 21364 10013 21373 10047
rect 21373 10013 21407 10047
rect 21407 10013 21416 10047
rect 21364 10004 21416 10013
rect 6368 9911 6420 9920
rect 6368 9877 6377 9911
rect 6377 9877 6411 9911
rect 6411 9877 6420 9911
rect 6368 9868 6420 9877
rect 8944 9868 8996 9920
rect 13268 9868 13320 9920
rect 16580 9868 16632 9920
rect 20168 9868 20220 9920
rect 22284 9868 22336 9920
rect 6630 9766 6682 9818
rect 6694 9766 6746 9818
rect 6758 9766 6810 9818
rect 6822 9766 6874 9818
rect 6886 9766 6938 9818
rect 12311 9766 12363 9818
rect 12375 9766 12427 9818
rect 12439 9766 12491 9818
rect 12503 9766 12555 9818
rect 12567 9766 12619 9818
rect 17992 9766 18044 9818
rect 18056 9766 18108 9818
rect 18120 9766 18172 9818
rect 18184 9766 18236 9818
rect 18248 9766 18300 9818
rect 23673 9766 23725 9818
rect 23737 9766 23789 9818
rect 23801 9766 23853 9818
rect 23865 9766 23917 9818
rect 23929 9766 23981 9818
rect 2228 9707 2280 9716
rect 2228 9673 2237 9707
rect 2237 9673 2271 9707
rect 2271 9673 2280 9707
rect 2228 9664 2280 9673
rect 4068 9664 4120 9716
rect 6184 9664 6236 9716
rect 7012 9707 7064 9716
rect 7012 9673 7021 9707
rect 7021 9673 7055 9707
rect 7055 9673 7064 9707
rect 7012 9664 7064 9673
rect 3608 9596 3660 9648
rect 5540 9596 5592 9648
rect 2136 9571 2188 9580
rect 2136 9537 2148 9571
rect 2148 9537 2182 9571
rect 2182 9537 2188 9571
rect 2136 9528 2188 9537
rect 2320 9528 2372 9580
rect 2596 9528 2648 9580
rect 3240 9571 3292 9580
rect 3240 9537 3249 9571
rect 3249 9537 3283 9571
rect 3283 9537 3292 9571
rect 3240 9528 3292 9537
rect 4712 9528 4764 9580
rect 4988 9528 5040 9580
rect 5264 9571 5316 9580
rect 5264 9537 5273 9571
rect 5273 9537 5307 9571
rect 5307 9537 5316 9571
rect 5264 9528 5316 9537
rect 5908 9528 5960 9580
rect 7104 9528 7156 9580
rect 8484 9664 8536 9716
rect 9404 9664 9456 9716
rect 11244 9664 11296 9716
rect 11520 9664 11572 9716
rect 13268 9664 13320 9716
rect 14188 9664 14240 9716
rect 5724 9460 5776 9512
rect 4160 9392 4212 9444
rect 7012 9392 7064 9444
rect 7380 9571 7432 9580
rect 7380 9537 7425 9571
rect 7425 9537 7432 9571
rect 7380 9528 7432 9537
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 7656 9460 7708 9512
rect 8116 9392 8168 9444
rect 8852 9392 8904 9444
rect 8944 9392 8996 9444
rect 9312 9392 9364 9444
rect 9864 9528 9916 9580
rect 9772 9503 9824 9512
rect 9772 9469 9781 9503
rect 9781 9469 9815 9503
rect 9815 9469 9824 9503
rect 9772 9460 9824 9469
rect 10324 9503 10376 9512
rect 10324 9469 10333 9503
rect 10333 9469 10367 9503
rect 10367 9469 10376 9503
rect 10324 9460 10376 9469
rect 1676 9367 1728 9376
rect 1676 9333 1685 9367
rect 1685 9333 1719 9367
rect 1719 9333 1728 9367
rect 1676 9324 1728 9333
rect 2964 9324 3016 9376
rect 3332 9324 3384 9376
rect 4896 9324 4948 9376
rect 5356 9324 5408 9376
rect 7748 9324 7800 9376
rect 7932 9324 7984 9376
rect 10232 9324 10284 9376
rect 10508 9392 10560 9444
rect 11060 9596 11112 9648
rect 10968 9528 11020 9580
rect 12716 9596 12768 9648
rect 13728 9639 13780 9648
rect 13728 9605 13737 9639
rect 13737 9605 13771 9639
rect 13771 9605 13780 9639
rect 13728 9596 13780 9605
rect 13820 9596 13872 9648
rect 13912 9528 13964 9580
rect 14924 9596 14976 9648
rect 16304 9596 16356 9648
rect 17224 9596 17276 9648
rect 21088 9664 21140 9716
rect 22100 9664 22152 9716
rect 17684 9596 17736 9648
rect 14740 9528 14792 9580
rect 15108 9571 15160 9580
rect 15108 9537 15117 9571
rect 15117 9537 15151 9571
rect 15151 9537 15160 9571
rect 15108 9528 15160 9537
rect 16764 9528 16816 9580
rect 13360 9460 13412 9512
rect 14464 9392 14516 9444
rect 10876 9324 10928 9376
rect 12532 9324 12584 9376
rect 14832 9324 14884 9376
rect 16028 9460 16080 9512
rect 16396 9460 16448 9512
rect 18420 9571 18472 9580
rect 18420 9537 18429 9571
rect 18429 9537 18463 9571
rect 18463 9537 18472 9571
rect 18420 9528 18472 9537
rect 21180 9596 21232 9648
rect 21272 9596 21324 9648
rect 21548 9596 21600 9648
rect 19340 9571 19392 9580
rect 19340 9537 19349 9571
rect 19349 9537 19383 9571
rect 19383 9537 19392 9571
rect 19340 9528 19392 9537
rect 18328 9460 18380 9512
rect 18880 9460 18932 9512
rect 19248 9460 19300 9512
rect 20628 9528 20680 9580
rect 20812 9571 20864 9580
rect 20812 9537 20821 9571
rect 20821 9537 20855 9571
rect 20855 9537 20864 9571
rect 20812 9528 20864 9537
rect 21732 9528 21784 9580
rect 22008 9571 22060 9580
rect 22008 9537 22017 9571
rect 22017 9537 22051 9571
rect 22051 9537 22060 9571
rect 22008 9528 22060 9537
rect 20444 9460 20496 9512
rect 21180 9460 21232 9512
rect 22284 9392 22336 9444
rect 16856 9324 16908 9376
rect 17132 9367 17184 9376
rect 17132 9333 17141 9367
rect 17141 9333 17175 9367
rect 17175 9333 17184 9367
rect 17132 9324 17184 9333
rect 17224 9324 17276 9376
rect 18604 9324 18656 9376
rect 19432 9324 19484 9376
rect 21640 9324 21692 9376
rect 22100 9324 22152 9376
rect 22376 9324 22428 9376
rect 22652 9324 22704 9376
rect 3790 9222 3842 9274
rect 3854 9222 3906 9274
rect 3918 9222 3970 9274
rect 3982 9222 4034 9274
rect 4046 9222 4098 9274
rect 9471 9222 9523 9274
rect 9535 9222 9587 9274
rect 9599 9222 9651 9274
rect 9663 9222 9715 9274
rect 9727 9222 9779 9274
rect 15152 9222 15204 9274
rect 15216 9222 15268 9274
rect 15280 9222 15332 9274
rect 15344 9222 15396 9274
rect 15408 9222 15460 9274
rect 20833 9222 20885 9274
rect 20897 9222 20949 9274
rect 20961 9222 21013 9274
rect 21025 9222 21077 9274
rect 21089 9222 21141 9274
rect 5172 9163 5224 9172
rect 5172 9129 5181 9163
rect 5181 9129 5215 9163
rect 5215 9129 5224 9163
rect 5172 9120 5224 9129
rect 5356 9120 5408 9172
rect 6828 9120 6880 9172
rect 7196 9120 7248 9172
rect 9220 9120 9272 9172
rect 4528 9052 4580 9104
rect 2228 8984 2280 9036
rect 2412 8984 2464 9036
rect 2136 8916 2188 8968
rect 2504 8848 2556 8900
rect 2872 8916 2924 8968
rect 5172 8984 5224 9036
rect 6184 8984 6236 9036
rect 6828 9027 6880 9036
rect 6828 8993 6837 9027
rect 6837 8993 6871 9027
rect 6871 8993 6880 9027
rect 6828 8984 6880 8993
rect 7656 8984 7708 9036
rect 7840 8984 7892 9036
rect 10324 8984 10376 9036
rect 10600 8984 10652 9036
rect 6460 8916 6512 8968
rect 4160 8848 4212 8900
rect 4252 8891 4304 8900
rect 4252 8857 4261 8891
rect 4261 8857 4295 8891
rect 4295 8857 4304 8891
rect 4252 8848 4304 8857
rect 5080 8891 5132 8900
rect 5080 8857 5089 8891
rect 5089 8857 5123 8891
rect 5123 8857 5132 8891
rect 5080 8848 5132 8857
rect 5264 8848 5316 8900
rect 5448 8848 5500 8900
rect 7012 8916 7064 8968
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 8024 8848 8076 8900
rect 9588 8891 9640 8900
rect 9588 8857 9597 8891
rect 9597 8857 9631 8891
rect 9631 8857 9640 8891
rect 9588 8848 9640 8857
rect 11704 8959 11756 8968
rect 11704 8925 11713 8959
rect 11713 8925 11747 8959
rect 11747 8925 11756 8959
rect 11704 8916 11756 8925
rect 12164 8984 12216 9036
rect 11980 8959 12032 8968
rect 11980 8925 11989 8959
rect 11989 8925 12023 8959
rect 12023 8925 12032 8959
rect 11980 8916 12032 8925
rect 12532 8959 12584 8968
rect 12532 8925 12541 8959
rect 12541 8925 12575 8959
rect 12575 8925 12584 8959
rect 12532 8916 12584 8925
rect 14004 9052 14056 9104
rect 17868 9120 17920 9172
rect 15568 9052 15620 9104
rect 13360 8984 13412 9036
rect 14372 8984 14424 9036
rect 14556 9027 14608 9036
rect 14556 8993 14565 9027
rect 14565 8993 14599 9027
rect 14599 8993 14608 9027
rect 14556 8984 14608 8993
rect 14832 8984 14884 9036
rect 16488 8984 16540 9036
rect 13268 8959 13320 8968
rect 13268 8925 13277 8959
rect 13277 8925 13311 8959
rect 13311 8925 13320 8959
rect 13268 8916 13320 8925
rect 12808 8848 12860 8900
rect 13820 8916 13872 8968
rect 14280 8916 14332 8968
rect 14464 8959 14516 8968
rect 14464 8925 14473 8959
rect 14473 8925 14507 8959
rect 14507 8925 14516 8959
rect 14464 8916 14516 8925
rect 14740 8959 14792 8968
rect 14740 8925 14749 8959
rect 14749 8925 14783 8959
rect 14783 8925 14792 8959
rect 14740 8916 14792 8925
rect 14924 8959 14976 8968
rect 14924 8925 14933 8959
rect 14933 8925 14967 8959
rect 14967 8925 14976 8959
rect 14924 8916 14976 8925
rect 16028 8916 16080 8968
rect 18604 9052 18656 9104
rect 19156 9052 19208 9104
rect 19616 9052 19668 9104
rect 16856 9027 16908 9036
rect 16856 8993 16865 9027
rect 16865 8993 16899 9027
rect 16899 8993 16908 9027
rect 16856 8984 16908 8993
rect 17592 8984 17644 9036
rect 20996 9120 21048 9172
rect 20536 9052 20588 9104
rect 21088 9052 21140 9104
rect 18052 8916 18104 8968
rect 18696 8916 18748 8968
rect 20812 8984 20864 9036
rect 21272 9027 21324 9036
rect 21272 8993 21281 9027
rect 21281 8993 21315 9027
rect 21315 8993 21324 9027
rect 21272 8984 21324 8993
rect 22192 9120 22244 9172
rect 3056 8780 3108 8832
rect 3700 8780 3752 8832
rect 4068 8780 4120 8832
rect 10600 8780 10652 8832
rect 11336 8780 11388 8832
rect 15660 8780 15712 8832
rect 18328 8848 18380 8900
rect 19800 8848 19852 8900
rect 20536 8959 20588 8968
rect 20536 8925 20545 8959
rect 20545 8925 20579 8959
rect 20579 8925 20588 8959
rect 20536 8916 20588 8925
rect 21088 8916 21140 8968
rect 21824 8984 21876 9036
rect 22836 9120 22888 9172
rect 22744 9052 22796 9104
rect 21456 8959 21508 8968
rect 21456 8925 21465 8959
rect 21465 8925 21499 8959
rect 21499 8925 21508 8959
rect 21456 8916 21508 8925
rect 22468 8959 22520 8968
rect 22468 8925 22477 8959
rect 22477 8925 22511 8959
rect 22511 8925 22520 8959
rect 22468 8916 22520 8925
rect 23204 8916 23256 8968
rect 22836 8848 22888 8900
rect 16948 8780 17000 8832
rect 17868 8823 17920 8832
rect 17868 8789 17877 8823
rect 17877 8789 17911 8823
rect 17911 8789 17920 8823
rect 17868 8780 17920 8789
rect 18052 8780 18104 8832
rect 21364 8780 21416 8832
rect 21640 8823 21692 8832
rect 21640 8789 21649 8823
rect 21649 8789 21683 8823
rect 21683 8789 21692 8823
rect 21640 8780 21692 8789
rect 6630 8678 6682 8730
rect 6694 8678 6746 8730
rect 6758 8678 6810 8730
rect 6822 8678 6874 8730
rect 6886 8678 6938 8730
rect 12311 8678 12363 8730
rect 12375 8678 12427 8730
rect 12439 8678 12491 8730
rect 12503 8678 12555 8730
rect 12567 8678 12619 8730
rect 17992 8678 18044 8730
rect 18056 8678 18108 8730
rect 18120 8678 18172 8730
rect 18184 8678 18236 8730
rect 18248 8678 18300 8730
rect 23673 8678 23725 8730
rect 23737 8678 23789 8730
rect 23801 8678 23853 8730
rect 23865 8678 23917 8730
rect 23929 8678 23981 8730
rect 7104 8576 7156 8628
rect 7748 8576 7800 8628
rect 2596 8440 2648 8492
rect 2964 8440 3016 8492
rect 4068 8508 4120 8560
rect 5172 8551 5224 8560
rect 5172 8517 5181 8551
rect 5181 8517 5215 8551
rect 5215 8517 5224 8551
rect 5172 8508 5224 8517
rect 6460 8508 6512 8560
rect 2504 8372 2556 8424
rect 3240 8415 3292 8424
rect 3240 8381 3249 8415
rect 3249 8381 3283 8415
rect 3283 8381 3292 8415
rect 3240 8372 3292 8381
rect 5356 8440 5408 8492
rect 2688 8304 2740 8356
rect 4528 8304 4580 8356
rect 4712 8304 4764 8356
rect 6552 8372 6604 8424
rect 8208 8508 8260 8560
rect 7656 8440 7708 8492
rect 8300 8440 8352 8492
rect 10140 8576 10192 8628
rect 12532 8576 12584 8628
rect 12164 8508 12216 8560
rect 14464 8576 14516 8628
rect 15476 8619 15528 8628
rect 15476 8585 15485 8619
rect 15485 8585 15519 8619
rect 15519 8585 15528 8619
rect 15476 8576 15528 8585
rect 15568 8619 15620 8628
rect 15568 8585 15577 8619
rect 15577 8585 15611 8619
rect 15611 8585 15620 8619
rect 15568 8576 15620 8585
rect 16212 8619 16264 8628
rect 16212 8585 16221 8619
rect 16221 8585 16255 8619
rect 16255 8585 16264 8619
rect 16212 8576 16264 8585
rect 16580 8576 16632 8628
rect 16948 8576 17000 8628
rect 18328 8576 18380 8628
rect 18972 8576 19024 8628
rect 19892 8576 19944 8628
rect 14372 8508 14424 8560
rect 16396 8508 16448 8560
rect 19064 8508 19116 8560
rect 6828 8304 6880 8356
rect 10048 8304 10100 8356
rect 11152 8440 11204 8492
rect 11428 8440 11480 8492
rect 11796 8440 11848 8492
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 13176 8440 13228 8492
rect 13268 8440 13320 8492
rect 10416 8415 10468 8424
rect 10416 8381 10425 8415
rect 10425 8381 10459 8415
rect 10459 8381 10468 8415
rect 10416 8372 10468 8381
rect 10600 8372 10652 8424
rect 13912 8440 13964 8492
rect 14004 8483 14056 8492
rect 14004 8449 14013 8483
rect 14013 8449 14047 8483
rect 14047 8449 14056 8483
rect 14004 8440 14056 8449
rect 14096 8483 14148 8492
rect 14096 8449 14105 8483
rect 14105 8449 14139 8483
rect 14139 8449 14148 8483
rect 14096 8440 14148 8449
rect 14188 8440 14240 8492
rect 11612 8304 11664 8356
rect 14556 8372 14608 8424
rect 15660 8440 15712 8492
rect 13820 8304 13872 8356
rect 16948 8372 17000 8424
rect 17500 8440 17552 8492
rect 18144 8483 18196 8492
rect 18144 8449 18153 8483
rect 18153 8449 18187 8483
rect 18187 8449 18196 8483
rect 18144 8440 18196 8449
rect 19156 8440 19208 8492
rect 19616 8508 19668 8560
rect 19432 8483 19484 8492
rect 19432 8449 19441 8483
rect 19441 8449 19475 8483
rect 19475 8449 19484 8483
rect 19432 8440 19484 8449
rect 17776 8372 17828 8424
rect 16764 8304 16816 8356
rect 17960 8304 18012 8356
rect 19892 8372 19944 8424
rect 20720 8576 20772 8628
rect 20628 8508 20680 8560
rect 20996 8551 21048 8560
rect 20996 8517 21005 8551
rect 21005 8517 21039 8551
rect 21039 8517 21048 8551
rect 20996 8508 21048 8517
rect 21088 8508 21140 8560
rect 20260 8483 20312 8492
rect 20260 8449 20269 8483
rect 20269 8449 20303 8483
rect 20303 8449 20312 8483
rect 20260 8440 20312 8449
rect 20352 8440 20404 8492
rect 21548 8440 21600 8492
rect 22284 8483 22336 8492
rect 22284 8449 22293 8483
rect 22293 8449 22327 8483
rect 22327 8449 22336 8483
rect 22284 8440 22336 8449
rect 22560 8440 22612 8492
rect 23020 8440 23072 8492
rect 21180 8372 21232 8424
rect 22376 8415 22428 8424
rect 22376 8381 22385 8415
rect 22385 8381 22419 8415
rect 22419 8381 22428 8415
rect 22376 8372 22428 8381
rect 2044 8236 2096 8288
rect 3056 8279 3108 8288
rect 3056 8245 3065 8279
rect 3065 8245 3099 8279
rect 3099 8245 3108 8279
rect 3056 8236 3108 8245
rect 3700 8236 3752 8288
rect 4160 8236 4212 8288
rect 5908 8236 5960 8288
rect 7656 8236 7708 8288
rect 7748 8279 7800 8288
rect 7748 8245 7757 8279
rect 7757 8245 7791 8279
rect 7791 8245 7800 8279
rect 7748 8236 7800 8245
rect 8484 8236 8536 8288
rect 8852 8236 8904 8288
rect 9588 8236 9640 8288
rect 10784 8236 10836 8288
rect 11060 8236 11112 8288
rect 19524 8236 19576 8288
rect 20352 8236 20404 8288
rect 3790 8134 3842 8186
rect 3854 8134 3906 8186
rect 3918 8134 3970 8186
rect 3982 8134 4034 8186
rect 4046 8134 4098 8186
rect 9471 8134 9523 8186
rect 9535 8134 9587 8186
rect 9599 8134 9651 8186
rect 9663 8134 9715 8186
rect 9727 8134 9779 8186
rect 15152 8134 15204 8186
rect 15216 8134 15268 8186
rect 15280 8134 15332 8186
rect 15344 8134 15396 8186
rect 15408 8134 15460 8186
rect 20833 8134 20885 8186
rect 20897 8134 20949 8186
rect 20961 8134 21013 8186
rect 21025 8134 21077 8186
rect 21089 8134 21141 8186
rect 2780 8032 2832 8084
rect 3056 8032 3108 8084
rect 4252 8032 4304 8084
rect 7380 8032 7432 8084
rect 8116 8075 8168 8084
rect 8116 8041 8125 8075
rect 8125 8041 8159 8075
rect 8159 8041 8168 8075
rect 8116 8032 8168 8041
rect 4160 7964 4212 8016
rect 5172 7964 5224 8016
rect 6920 7964 6972 8016
rect 9128 7964 9180 8016
rect 2504 7828 2556 7880
rect 3424 7828 3476 7880
rect 4528 7871 4580 7880
rect 4528 7837 4537 7871
rect 4537 7837 4571 7871
rect 4571 7837 4580 7871
rect 4528 7828 4580 7837
rect 2596 7760 2648 7812
rect 2780 7760 2832 7812
rect 8116 7896 8168 7948
rect 9772 8032 9824 8084
rect 10600 8032 10652 8084
rect 11704 8032 11756 8084
rect 12072 8032 12124 8084
rect 10048 7964 10100 8016
rect 5080 7828 5132 7880
rect 5356 7828 5408 7880
rect 6920 7871 6972 7880
rect 6920 7837 6929 7871
rect 6929 7837 6963 7871
rect 6963 7837 6972 7871
rect 6920 7828 6972 7837
rect 7748 7871 7800 7880
rect 7748 7837 7757 7871
rect 7757 7837 7791 7871
rect 7791 7837 7800 7871
rect 7748 7828 7800 7837
rect 9128 7871 9180 7880
rect 5908 7760 5960 7812
rect 6184 7760 6236 7812
rect 5356 7692 5408 7744
rect 7380 7760 7432 7812
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 9128 7828 9180 7837
rect 10232 7896 10284 7948
rect 13728 8075 13780 8084
rect 13728 8041 13737 8075
rect 13737 8041 13771 8075
rect 13771 8041 13780 8075
rect 13728 8032 13780 8041
rect 14740 8032 14792 8084
rect 15476 8032 15528 8084
rect 15844 8075 15896 8084
rect 15844 8041 15853 8075
rect 15853 8041 15887 8075
rect 15887 8041 15896 8075
rect 15844 8032 15896 8041
rect 17132 8032 17184 8084
rect 18420 8075 18472 8084
rect 18420 8041 18429 8075
rect 18429 8041 18463 8075
rect 18463 8041 18472 8075
rect 18420 8032 18472 8041
rect 16856 7964 16908 8016
rect 17040 7964 17092 8016
rect 17408 7964 17460 8016
rect 20536 8032 20588 8084
rect 22744 8075 22796 8084
rect 22744 8041 22753 8075
rect 22753 8041 22787 8075
rect 22787 8041 22796 8075
rect 22744 8032 22796 8041
rect 8392 7760 8444 7812
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 15660 7896 15712 7948
rect 17316 7896 17368 7948
rect 22284 7964 22336 8016
rect 20260 7896 20312 7948
rect 11428 7828 11480 7880
rect 8944 7692 8996 7744
rect 11336 7760 11388 7812
rect 12164 7828 12216 7880
rect 12808 7871 12860 7880
rect 12808 7837 12817 7871
rect 12817 7837 12851 7871
rect 12851 7837 12860 7871
rect 12808 7828 12860 7837
rect 12716 7760 12768 7812
rect 13084 7803 13136 7812
rect 13084 7769 13093 7803
rect 13093 7769 13127 7803
rect 13127 7769 13136 7803
rect 13084 7760 13136 7769
rect 14648 7871 14700 7880
rect 14648 7837 14657 7871
rect 14657 7837 14691 7871
rect 14691 7837 14700 7871
rect 14648 7828 14700 7837
rect 15200 7828 15252 7880
rect 15568 7828 15620 7880
rect 15936 7828 15988 7880
rect 16856 7871 16908 7880
rect 16856 7837 16865 7871
rect 16865 7837 16899 7871
rect 16899 7837 16908 7871
rect 16856 7828 16908 7837
rect 16488 7760 16540 7812
rect 17224 7871 17276 7880
rect 17224 7837 17233 7871
rect 17233 7837 17267 7871
rect 17267 7837 17276 7871
rect 17224 7828 17276 7837
rect 17408 7871 17460 7880
rect 17408 7837 17417 7871
rect 17417 7837 17451 7871
rect 17451 7837 17460 7871
rect 17408 7828 17460 7837
rect 17776 7828 17828 7880
rect 18144 7760 18196 7812
rect 18696 7828 18748 7880
rect 19616 7871 19668 7880
rect 19616 7837 19625 7871
rect 19625 7837 19659 7871
rect 19659 7837 19668 7871
rect 19616 7828 19668 7837
rect 19984 7760 20036 7812
rect 12992 7692 13044 7744
rect 15016 7692 15068 7744
rect 15568 7692 15620 7744
rect 16764 7692 16816 7744
rect 19432 7692 19484 7744
rect 20720 7828 20772 7880
rect 21180 7828 21232 7880
rect 20168 7760 20220 7812
rect 22560 7692 22612 7744
rect 6630 7590 6682 7642
rect 6694 7590 6746 7642
rect 6758 7590 6810 7642
rect 6822 7590 6874 7642
rect 6886 7590 6938 7642
rect 12311 7590 12363 7642
rect 12375 7590 12427 7642
rect 12439 7590 12491 7642
rect 12503 7590 12555 7642
rect 12567 7590 12619 7642
rect 17992 7590 18044 7642
rect 18056 7590 18108 7642
rect 18120 7590 18172 7642
rect 18184 7590 18236 7642
rect 18248 7590 18300 7642
rect 23673 7590 23725 7642
rect 23737 7590 23789 7642
rect 23801 7590 23853 7642
rect 23865 7590 23917 7642
rect 23929 7590 23981 7642
rect 2136 7488 2188 7540
rect 4528 7488 4580 7540
rect 2320 7420 2372 7472
rect 2780 7395 2832 7404
rect 2780 7361 2789 7395
rect 2789 7361 2823 7395
rect 2823 7361 2832 7395
rect 2780 7352 2832 7361
rect 4160 7352 4212 7404
rect 1860 7284 1912 7336
rect 3148 7284 3200 7336
rect 8392 7531 8444 7540
rect 8392 7497 8401 7531
rect 8401 7497 8435 7531
rect 8435 7497 8444 7531
rect 8392 7488 8444 7497
rect 9128 7488 9180 7540
rect 9864 7488 9916 7540
rect 10232 7531 10284 7540
rect 10232 7497 10241 7531
rect 10241 7497 10275 7531
rect 10275 7497 10284 7531
rect 10232 7488 10284 7497
rect 10324 7488 10376 7540
rect 15016 7488 15068 7540
rect 15200 7531 15252 7540
rect 15200 7497 15209 7531
rect 15209 7497 15243 7531
rect 15243 7497 15252 7531
rect 15200 7488 15252 7497
rect 21732 7488 21784 7540
rect 22744 7488 22796 7540
rect 5356 7420 5408 7472
rect 4896 7352 4948 7404
rect 6552 7352 6604 7404
rect 7012 7395 7064 7404
rect 7012 7361 7021 7395
rect 7021 7361 7055 7395
rect 7055 7361 7064 7395
rect 8484 7420 8536 7472
rect 7012 7352 7064 7361
rect 7748 7352 7800 7404
rect 8116 7395 8168 7404
rect 8116 7361 8125 7395
rect 8125 7361 8159 7395
rect 8159 7361 8168 7395
rect 8116 7352 8168 7361
rect 8852 7395 8904 7404
rect 8852 7361 8861 7395
rect 8861 7361 8895 7395
rect 8895 7361 8904 7395
rect 8852 7352 8904 7361
rect 9036 7395 9088 7404
rect 9036 7361 9045 7395
rect 9045 7361 9079 7395
rect 9079 7361 9088 7395
rect 9036 7352 9088 7361
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 10968 7420 11020 7472
rect 11152 7463 11204 7472
rect 11152 7429 11161 7463
rect 11161 7429 11195 7463
rect 11195 7429 11204 7463
rect 11152 7420 11204 7429
rect 12256 7420 12308 7472
rect 14648 7420 14700 7472
rect 17408 7420 17460 7472
rect 17592 7463 17644 7472
rect 17592 7429 17601 7463
rect 17601 7429 17635 7463
rect 17635 7429 17644 7463
rect 17592 7420 17644 7429
rect 7932 7284 7984 7336
rect 8944 7284 8996 7336
rect 10416 7352 10468 7404
rect 12072 7352 12124 7404
rect 14096 7352 14148 7404
rect 14280 7395 14332 7404
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 15844 7352 15896 7404
rect 16764 7352 16816 7404
rect 17040 7395 17092 7404
rect 17040 7361 17046 7395
rect 17046 7361 17092 7395
rect 17040 7352 17092 7361
rect 18328 7352 18380 7404
rect 18972 7352 19024 7404
rect 19156 7352 19208 7404
rect 11428 7284 11480 7336
rect 16580 7284 16632 7336
rect 19708 7284 19760 7336
rect 20260 7284 20312 7336
rect 20444 7284 20496 7336
rect 2412 7148 2464 7200
rect 5264 7191 5316 7200
rect 5264 7157 5273 7191
rect 5273 7157 5307 7191
rect 5307 7157 5316 7191
rect 5264 7148 5316 7157
rect 5816 7191 5868 7200
rect 5816 7157 5825 7191
rect 5825 7157 5859 7191
rect 5859 7157 5868 7191
rect 5816 7148 5868 7157
rect 6276 7148 6328 7200
rect 6552 7148 6604 7200
rect 8300 7216 8352 7268
rect 8852 7216 8904 7268
rect 17132 7259 17184 7268
rect 17132 7225 17141 7259
rect 17141 7225 17175 7259
rect 17175 7225 17184 7259
rect 17132 7216 17184 7225
rect 22468 7216 22520 7268
rect 22836 7352 22888 7404
rect 8116 7191 8168 7200
rect 8116 7157 8125 7191
rect 8125 7157 8159 7191
rect 8159 7157 8168 7191
rect 8116 7148 8168 7157
rect 10324 7148 10376 7200
rect 12716 7191 12768 7200
rect 12716 7157 12725 7191
rect 12725 7157 12759 7191
rect 12759 7157 12768 7191
rect 12716 7148 12768 7157
rect 13360 7148 13412 7200
rect 15016 7148 15068 7200
rect 22744 7148 22796 7200
rect 3790 7046 3842 7098
rect 3854 7046 3906 7098
rect 3918 7046 3970 7098
rect 3982 7046 4034 7098
rect 4046 7046 4098 7098
rect 9471 7046 9523 7098
rect 9535 7046 9587 7098
rect 9599 7046 9651 7098
rect 9663 7046 9715 7098
rect 9727 7046 9779 7098
rect 15152 7046 15204 7098
rect 15216 7046 15268 7098
rect 15280 7046 15332 7098
rect 15344 7046 15396 7098
rect 15408 7046 15460 7098
rect 20833 7046 20885 7098
rect 20897 7046 20949 7098
rect 20961 7046 21013 7098
rect 21025 7046 21077 7098
rect 21089 7046 21141 7098
rect 2780 6944 2832 6996
rect 9036 6944 9088 6996
rect 10416 6944 10468 6996
rect 13084 6944 13136 6996
rect 16580 6944 16632 6996
rect 2136 6740 2188 6792
rect 4528 6808 4580 6860
rect 4620 6808 4672 6860
rect 2688 6604 2740 6656
rect 3148 6604 3200 6656
rect 4252 6604 4304 6656
rect 5264 6808 5316 6860
rect 5724 6740 5776 6792
rect 5816 6783 5868 6792
rect 5816 6749 5825 6783
rect 5825 6749 5859 6783
rect 5859 6749 5868 6783
rect 5816 6740 5868 6749
rect 8392 6876 8444 6928
rect 5448 6672 5500 6724
rect 7840 6740 7892 6792
rect 8208 6808 8260 6860
rect 11704 6876 11756 6928
rect 6828 6715 6880 6724
rect 6828 6681 6837 6715
rect 6837 6681 6871 6715
rect 6871 6681 6880 6715
rect 6828 6672 6880 6681
rect 5540 6604 5592 6656
rect 5724 6604 5776 6656
rect 8116 6740 8168 6792
rect 8300 6783 8352 6792
rect 8300 6749 8309 6783
rect 8309 6749 8343 6783
rect 8343 6749 8352 6783
rect 8300 6740 8352 6749
rect 9956 6851 10008 6860
rect 9956 6817 9965 6851
rect 9965 6817 9999 6851
rect 9999 6817 10008 6851
rect 9956 6808 10008 6817
rect 10048 6808 10100 6860
rect 10324 6851 10376 6860
rect 10324 6817 10333 6851
rect 10333 6817 10367 6851
rect 10367 6817 10376 6851
rect 10324 6808 10376 6817
rect 12164 6808 12216 6860
rect 12992 6876 13044 6928
rect 13728 6876 13780 6928
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 10876 6740 10928 6792
rect 10968 6740 11020 6792
rect 12072 6740 12124 6792
rect 13452 6783 13504 6792
rect 13452 6749 13461 6783
rect 13461 6749 13495 6783
rect 13495 6749 13504 6783
rect 13452 6740 13504 6749
rect 13912 6808 13964 6860
rect 14096 6740 14148 6792
rect 14280 6740 14332 6792
rect 17040 6808 17092 6860
rect 18328 6808 18380 6860
rect 18972 6808 19024 6860
rect 16120 6740 16172 6792
rect 19064 6740 19116 6792
rect 19340 6740 19392 6792
rect 19432 6783 19484 6792
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 19248 6672 19300 6724
rect 20628 6740 20680 6792
rect 21272 6783 21324 6792
rect 21272 6749 21281 6783
rect 21281 6749 21315 6783
rect 21315 6749 21324 6783
rect 21272 6740 21324 6749
rect 9680 6604 9732 6656
rect 10324 6604 10376 6656
rect 10600 6604 10652 6656
rect 11612 6604 11664 6656
rect 12256 6604 12308 6656
rect 13176 6604 13228 6656
rect 15568 6604 15620 6656
rect 18880 6604 18932 6656
rect 20536 6604 20588 6656
rect 21548 6740 21600 6792
rect 22192 6851 22244 6860
rect 22192 6817 22201 6851
rect 22201 6817 22235 6851
rect 22235 6817 22244 6851
rect 22192 6808 22244 6817
rect 22652 6851 22704 6860
rect 22652 6817 22661 6851
rect 22661 6817 22695 6851
rect 22695 6817 22704 6851
rect 22652 6808 22704 6817
rect 21640 6672 21692 6724
rect 22744 6783 22796 6792
rect 22744 6749 22753 6783
rect 22753 6749 22787 6783
rect 22787 6749 22796 6783
rect 22744 6740 22796 6749
rect 22100 6604 22152 6656
rect 6630 6502 6682 6554
rect 6694 6502 6746 6554
rect 6758 6502 6810 6554
rect 6822 6502 6874 6554
rect 6886 6502 6938 6554
rect 12311 6502 12363 6554
rect 12375 6502 12427 6554
rect 12439 6502 12491 6554
rect 12503 6502 12555 6554
rect 12567 6502 12619 6554
rect 17992 6502 18044 6554
rect 18056 6502 18108 6554
rect 18120 6502 18172 6554
rect 18184 6502 18236 6554
rect 18248 6502 18300 6554
rect 23673 6502 23725 6554
rect 23737 6502 23789 6554
rect 23801 6502 23853 6554
rect 23865 6502 23917 6554
rect 23929 6502 23981 6554
rect 9680 6400 9732 6452
rect 10048 6400 10100 6452
rect 4344 6332 4396 6384
rect 2228 6307 2280 6316
rect 2228 6273 2237 6307
rect 2237 6273 2271 6307
rect 2271 6273 2280 6307
rect 2228 6264 2280 6273
rect 2412 6307 2464 6316
rect 2412 6273 2421 6307
rect 2421 6273 2455 6307
rect 2455 6273 2464 6307
rect 2412 6264 2464 6273
rect 2688 6307 2740 6316
rect 2688 6273 2697 6307
rect 2697 6273 2731 6307
rect 2731 6273 2740 6307
rect 2688 6264 2740 6273
rect 2964 6307 3016 6316
rect 2964 6273 2973 6307
rect 2973 6273 3007 6307
rect 3007 6273 3016 6307
rect 2964 6264 3016 6273
rect 3056 6307 3108 6316
rect 3056 6273 3065 6307
rect 3065 6273 3099 6307
rect 3099 6273 3108 6307
rect 3056 6264 3108 6273
rect 4436 6264 4488 6316
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 5448 6264 5500 6316
rect 5908 6264 5960 6316
rect 6644 6264 6696 6316
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 8208 6264 8260 6316
rect 12072 6332 12124 6384
rect 2136 6128 2188 6180
rect 7748 6196 7800 6248
rect 8944 6307 8996 6316
rect 8944 6273 8953 6307
rect 8953 6273 8987 6307
rect 8987 6273 8996 6307
rect 8944 6264 8996 6273
rect 11060 6196 11112 6248
rect 12256 6196 12308 6248
rect 18328 6400 18380 6452
rect 18788 6400 18840 6452
rect 22376 6400 22428 6452
rect 23020 6443 23072 6452
rect 23020 6409 23029 6443
rect 23029 6409 23063 6443
rect 23063 6409 23072 6443
rect 23020 6400 23072 6409
rect 13176 6375 13228 6384
rect 13176 6341 13185 6375
rect 13185 6341 13219 6375
rect 13219 6341 13228 6375
rect 13176 6332 13228 6341
rect 13452 6264 13504 6316
rect 3056 6128 3108 6180
rect 4160 6128 4212 6180
rect 4896 6128 4948 6180
rect 4988 6128 5040 6180
rect 16488 6332 16540 6384
rect 19616 6332 19668 6384
rect 15568 6264 15620 6316
rect 17132 6264 17184 6316
rect 17408 6307 17460 6316
rect 17408 6273 17417 6307
rect 17417 6273 17451 6307
rect 17451 6273 17460 6307
rect 17408 6264 17460 6273
rect 14096 6239 14148 6248
rect 14096 6205 14105 6239
rect 14105 6205 14139 6239
rect 14139 6205 14148 6239
rect 14096 6196 14148 6205
rect 14556 6196 14608 6248
rect 14740 6239 14792 6248
rect 14740 6205 14749 6239
rect 14749 6205 14783 6239
rect 14783 6205 14792 6239
rect 14740 6196 14792 6205
rect 15016 6196 15068 6248
rect 15568 6128 15620 6180
rect 4252 6060 4304 6112
rect 4436 6060 4488 6112
rect 5816 6060 5868 6112
rect 6368 6060 6420 6112
rect 9312 6060 9364 6112
rect 9404 6060 9456 6112
rect 13544 6060 13596 6112
rect 13636 6103 13688 6112
rect 13636 6069 13645 6103
rect 13645 6069 13679 6103
rect 13679 6069 13688 6103
rect 13636 6060 13688 6069
rect 14004 6103 14056 6112
rect 14004 6069 14013 6103
rect 14013 6069 14047 6103
rect 14047 6069 14056 6103
rect 14004 6060 14056 6069
rect 15476 6060 15528 6112
rect 15752 6239 15804 6248
rect 15752 6205 15761 6239
rect 15761 6205 15795 6239
rect 15795 6205 15804 6239
rect 15752 6196 15804 6205
rect 16764 6196 16816 6248
rect 15936 6128 15988 6180
rect 18236 6196 18288 6248
rect 18788 6307 18840 6316
rect 18788 6273 18797 6307
rect 18797 6273 18831 6307
rect 18831 6273 18840 6307
rect 18788 6264 18840 6273
rect 20444 6375 20496 6384
rect 20444 6341 20453 6375
rect 20453 6341 20487 6375
rect 20487 6341 20496 6375
rect 20444 6332 20496 6341
rect 19984 6307 20036 6316
rect 19984 6273 19993 6307
rect 19993 6273 20027 6307
rect 20027 6273 20036 6307
rect 19984 6264 20036 6273
rect 22468 6332 22520 6384
rect 21272 6307 21324 6316
rect 21272 6273 21281 6307
rect 21281 6273 21315 6307
rect 21315 6273 21324 6307
rect 21272 6264 21324 6273
rect 22008 6307 22060 6316
rect 22008 6273 22017 6307
rect 22017 6273 22051 6307
rect 22051 6273 22060 6307
rect 22008 6264 22060 6273
rect 23204 6307 23256 6316
rect 19156 6196 19208 6248
rect 19432 6196 19484 6248
rect 20168 6196 20220 6248
rect 23204 6273 23213 6307
rect 23213 6273 23247 6307
rect 23247 6273 23256 6307
rect 23204 6264 23256 6273
rect 17500 6128 17552 6180
rect 18972 6128 19024 6180
rect 23296 6239 23348 6248
rect 23296 6205 23305 6239
rect 23305 6205 23339 6239
rect 23339 6205 23348 6239
rect 23296 6196 23348 6205
rect 16672 6060 16724 6112
rect 22652 6060 22704 6112
rect 22836 6060 22888 6112
rect 3790 5958 3842 6010
rect 3854 5958 3906 6010
rect 3918 5958 3970 6010
rect 3982 5958 4034 6010
rect 4046 5958 4098 6010
rect 9471 5958 9523 6010
rect 9535 5958 9587 6010
rect 9599 5958 9651 6010
rect 9663 5958 9715 6010
rect 9727 5958 9779 6010
rect 15152 5958 15204 6010
rect 15216 5958 15268 6010
rect 15280 5958 15332 6010
rect 15344 5958 15396 6010
rect 15408 5958 15460 6010
rect 20833 5958 20885 6010
rect 20897 5958 20949 6010
rect 20961 5958 21013 6010
rect 21025 5958 21077 6010
rect 21089 5958 21141 6010
rect 2136 5899 2188 5908
rect 2136 5865 2145 5899
rect 2145 5865 2179 5899
rect 2179 5865 2188 5899
rect 2136 5856 2188 5865
rect 2228 5856 2280 5908
rect 5540 5856 5592 5908
rect 2688 5788 2740 5840
rect 3056 5788 3108 5840
rect 4344 5788 4396 5840
rect 6368 5788 6420 5840
rect 2228 5584 2280 5636
rect 2504 5652 2556 5704
rect 3056 5652 3108 5704
rect 6092 5720 6144 5772
rect 7932 5788 7984 5840
rect 8392 5856 8444 5908
rect 9220 5899 9272 5908
rect 9220 5865 9229 5899
rect 9229 5865 9263 5899
rect 9263 5865 9272 5899
rect 9220 5856 9272 5865
rect 11980 5856 12032 5908
rect 12164 5856 12216 5908
rect 15936 5856 15988 5908
rect 16396 5899 16448 5908
rect 16396 5865 16405 5899
rect 16405 5865 16439 5899
rect 16439 5865 16448 5899
rect 16396 5856 16448 5865
rect 18788 5856 18840 5908
rect 19892 5856 19944 5908
rect 21272 5899 21324 5908
rect 21272 5865 21281 5899
rect 21281 5865 21315 5899
rect 21315 5865 21324 5899
rect 21272 5856 21324 5865
rect 22468 5856 22520 5908
rect 8300 5788 8352 5840
rect 8484 5788 8536 5840
rect 9588 5788 9640 5840
rect 11336 5788 11388 5840
rect 11796 5788 11848 5840
rect 11888 5788 11940 5840
rect 4160 5695 4212 5704
rect 4160 5661 4169 5695
rect 4169 5661 4203 5695
rect 4203 5661 4212 5695
rect 4160 5652 4212 5661
rect 4436 5652 4488 5704
rect 4712 5652 4764 5704
rect 4988 5652 5040 5704
rect 2872 5584 2924 5636
rect 3608 5584 3660 5636
rect 2044 5516 2096 5568
rect 2412 5516 2464 5568
rect 3240 5516 3292 5568
rect 4068 5516 4120 5568
rect 5540 5584 5592 5636
rect 6552 5652 6604 5704
rect 6644 5627 6696 5636
rect 6644 5593 6653 5627
rect 6653 5593 6687 5627
rect 6687 5593 6696 5627
rect 6644 5584 6696 5593
rect 5632 5516 5684 5568
rect 5724 5559 5776 5568
rect 5724 5525 5759 5559
rect 5759 5525 5776 5559
rect 5724 5516 5776 5525
rect 6460 5516 6512 5568
rect 6828 5559 6880 5568
rect 6828 5525 6837 5559
rect 6837 5525 6871 5559
rect 6871 5525 6880 5559
rect 6828 5516 6880 5525
rect 8208 5763 8260 5772
rect 8208 5729 8217 5763
rect 8217 5729 8251 5763
rect 8251 5729 8260 5763
rect 8208 5720 8260 5729
rect 8300 5652 8352 5704
rect 10508 5652 10560 5704
rect 10600 5695 10652 5704
rect 10600 5661 10609 5695
rect 10609 5661 10643 5695
rect 10643 5661 10652 5695
rect 10600 5652 10652 5661
rect 11060 5695 11112 5704
rect 11060 5661 11069 5695
rect 11069 5661 11103 5695
rect 11103 5661 11112 5695
rect 11060 5652 11112 5661
rect 12256 5720 12308 5772
rect 20076 5788 20128 5840
rect 20168 5831 20220 5840
rect 20168 5797 20177 5831
rect 20177 5797 20211 5831
rect 20211 5797 20220 5831
rect 20168 5788 20220 5797
rect 13636 5720 13688 5772
rect 17132 5720 17184 5772
rect 11336 5695 11388 5704
rect 11336 5661 11345 5695
rect 11345 5661 11379 5695
rect 11379 5661 11388 5695
rect 11336 5652 11388 5661
rect 11428 5695 11480 5704
rect 11428 5661 11437 5695
rect 11437 5661 11471 5695
rect 11471 5661 11480 5695
rect 11428 5652 11480 5661
rect 11704 5584 11756 5636
rect 11796 5516 11848 5568
rect 13360 5695 13412 5704
rect 13360 5661 13369 5695
rect 13369 5661 13403 5695
rect 13403 5661 13412 5695
rect 13360 5652 13412 5661
rect 14740 5652 14792 5704
rect 15108 5695 15160 5704
rect 15108 5661 15117 5695
rect 15117 5661 15151 5695
rect 15151 5661 15160 5695
rect 15108 5652 15160 5661
rect 16028 5652 16080 5704
rect 16304 5652 16356 5704
rect 16580 5695 16632 5704
rect 16580 5661 16589 5695
rect 16589 5661 16623 5695
rect 16623 5661 16632 5695
rect 16580 5652 16632 5661
rect 16948 5652 17000 5704
rect 17500 5763 17552 5772
rect 17500 5729 17509 5763
rect 17509 5729 17543 5763
rect 17543 5729 17552 5763
rect 17500 5720 17552 5729
rect 18236 5763 18288 5772
rect 18236 5729 18245 5763
rect 18245 5729 18279 5763
rect 18279 5729 18288 5763
rect 18236 5720 18288 5729
rect 19800 5720 19852 5772
rect 17316 5652 17368 5704
rect 19616 5652 19668 5704
rect 20628 5763 20680 5772
rect 20628 5729 20637 5763
rect 20637 5729 20671 5763
rect 20671 5729 20680 5763
rect 20628 5720 20680 5729
rect 22284 5763 22336 5772
rect 22284 5729 22293 5763
rect 22293 5729 22327 5763
rect 22327 5729 22336 5763
rect 22284 5720 22336 5729
rect 22928 5763 22980 5772
rect 22928 5729 22937 5763
rect 22937 5729 22971 5763
rect 22971 5729 22980 5763
rect 22928 5720 22980 5729
rect 14924 5584 14976 5636
rect 12716 5516 12768 5568
rect 15844 5584 15896 5636
rect 22100 5695 22152 5704
rect 22100 5661 22109 5695
rect 22109 5661 22143 5695
rect 22143 5661 22152 5695
rect 22100 5652 22152 5661
rect 22560 5652 22612 5704
rect 20628 5584 20680 5636
rect 6630 5414 6682 5466
rect 6694 5414 6746 5466
rect 6758 5414 6810 5466
rect 6822 5414 6874 5466
rect 6886 5414 6938 5466
rect 12311 5414 12363 5466
rect 12375 5414 12427 5466
rect 12439 5414 12491 5466
rect 12503 5414 12555 5466
rect 12567 5414 12619 5466
rect 17992 5414 18044 5466
rect 18056 5414 18108 5466
rect 18120 5414 18172 5466
rect 18184 5414 18236 5466
rect 18248 5414 18300 5466
rect 23673 5414 23725 5466
rect 23737 5414 23789 5466
rect 23801 5414 23853 5466
rect 23865 5414 23917 5466
rect 23929 5414 23981 5466
rect 4620 5312 4672 5364
rect 6368 5312 6420 5364
rect 2228 5176 2280 5228
rect 2504 5244 2556 5296
rect 3700 5244 3752 5296
rect 4068 5244 4120 5296
rect 3148 5176 3200 5228
rect 2688 5108 2740 5160
rect 2872 5108 2924 5160
rect 3516 5151 3568 5160
rect 3516 5117 3525 5151
rect 3525 5117 3559 5151
rect 3559 5117 3568 5151
rect 3516 5108 3568 5117
rect 4528 5176 4580 5228
rect 5080 5176 5132 5228
rect 5816 5176 5868 5228
rect 11336 5312 11388 5364
rect 12716 5312 12768 5364
rect 13268 5312 13320 5364
rect 14740 5312 14792 5364
rect 14924 5312 14976 5364
rect 15476 5312 15528 5364
rect 16304 5312 16356 5364
rect 16856 5312 16908 5364
rect 19248 5355 19300 5364
rect 19248 5321 19257 5355
rect 19257 5321 19291 5355
rect 19291 5321 19300 5355
rect 19248 5312 19300 5321
rect 19984 5312 20036 5364
rect 7104 5244 7156 5296
rect 9220 5244 9272 5296
rect 7012 5176 7064 5228
rect 8300 5176 8352 5228
rect 8852 5176 8904 5228
rect 4988 5151 5040 5160
rect 4988 5117 4997 5151
rect 4997 5117 5031 5151
rect 5031 5117 5040 5151
rect 4988 5108 5040 5117
rect 5724 5151 5776 5160
rect 5724 5117 5733 5151
rect 5733 5117 5767 5151
rect 5767 5117 5776 5151
rect 5724 5108 5776 5117
rect 6092 5108 6144 5160
rect 6920 5040 6972 5092
rect 6644 5015 6696 5024
rect 6644 4981 6653 5015
rect 6653 4981 6687 5015
rect 6687 4981 6696 5015
rect 6644 4972 6696 4981
rect 8576 5108 8628 5160
rect 9864 5176 9916 5228
rect 15292 5287 15344 5296
rect 15292 5253 15301 5287
rect 15301 5253 15335 5287
rect 15335 5253 15344 5287
rect 15292 5244 15344 5253
rect 16948 5244 17000 5296
rect 17500 5287 17552 5296
rect 17500 5253 17509 5287
rect 17509 5253 17543 5287
rect 17543 5253 17552 5287
rect 17500 5244 17552 5253
rect 21180 5355 21232 5364
rect 21180 5321 21189 5355
rect 21189 5321 21223 5355
rect 21223 5321 21232 5355
rect 21180 5312 21232 5321
rect 22836 5312 22888 5364
rect 9588 5151 9640 5160
rect 9588 5117 9597 5151
rect 9597 5117 9631 5151
rect 9631 5117 9640 5151
rect 9588 5108 9640 5117
rect 8024 5040 8076 5092
rect 10508 5219 10560 5228
rect 10508 5185 10517 5219
rect 10517 5185 10551 5219
rect 10551 5185 10560 5219
rect 10508 5176 10560 5185
rect 10692 5219 10744 5228
rect 10692 5185 10701 5219
rect 10701 5185 10735 5219
rect 10735 5185 10744 5219
rect 10692 5176 10744 5185
rect 10876 5176 10928 5228
rect 11796 5176 11848 5228
rect 11980 5176 12032 5228
rect 12716 5219 12768 5228
rect 12716 5185 12725 5219
rect 12725 5185 12759 5219
rect 12759 5185 12768 5219
rect 12716 5176 12768 5185
rect 12808 5219 12860 5228
rect 12808 5185 12817 5219
rect 12817 5185 12851 5219
rect 12851 5185 12860 5219
rect 12808 5176 12860 5185
rect 12900 5176 12952 5228
rect 14004 5176 14056 5228
rect 14648 5176 14700 5228
rect 15476 5176 15528 5228
rect 15844 5176 15896 5228
rect 18144 5219 18196 5228
rect 18144 5185 18153 5219
rect 18153 5185 18187 5219
rect 18187 5185 18196 5219
rect 18144 5176 18196 5185
rect 18328 5176 18380 5228
rect 18420 5219 18472 5228
rect 18420 5185 18429 5219
rect 18429 5185 18463 5219
rect 18463 5185 18472 5219
rect 18420 5176 18472 5185
rect 20260 5176 20312 5228
rect 20628 5176 20680 5228
rect 22100 5244 22152 5296
rect 22928 5244 22980 5296
rect 21272 5219 21324 5228
rect 21272 5185 21281 5219
rect 21281 5185 21315 5219
rect 21315 5185 21324 5219
rect 21272 5176 21324 5185
rect 22836 5176 22888 5228
rect 20444 5108 20496 5160
rect 12900 5040 12952 5092
rect 15476 5040 15528 5092
rect 8760 4972 8812 5024
rect 13360 4972 13412 5024
rect 13636 4972 13688 5024
rect 13912 4972 13964 5024
rect 15292 4972 15344 5024
rect 17500 5040 17552 5092
rect 19800 5040 19852 5092
rect 17316 5015 17368 5024
rect 17316 4981 17325 5015
rect 17325 4981 17359 5015
rect 17359 4981 17368 5015
rect 17316 4972 17368 4981
rect 3790 4870 3842 4922
rect 3854 4870 3906 4922
rect 3918 4870 3970 4922
rect 3982 4870 4034 4922
rect 4046 4870 4098 4922
rect 9471 4870 9523 4922
rect 9535 4870 9587 4922
rect 9599 4870 9651 4922
rect 9663 4870 9715 4922
rect 9727 4870 9779 4922
rect 15152 4870 15204 4922
rect 15216 4870 15268 4922
rect 15280 4870 15332 4922
rect 15344 4870 15396 4922
rect 15408 4870 15460 4922
rect 20833 4870 20885 4922
rect 20897 4870 20949 4922
rect 20961 4870 21013 4922
rect 21025 4870 21077 4922
rect 21089 4870 21141 4922
rect 7748 4768 7800 4820
rect 9128 4768 9180 4820
rect 11520 4768 11572 4820
rect 12072 4811 12124 4820
rect 12072 4777 12081 4811
rect 12081 4777 12115 4811
rect 12115 4777 12124 4811
rect 12072 4768 12124 4777
rect 12164 4768 12216 4820
rect 12716 4768 12768 4820
rect 13912 4768 13964 4820
rect 15016 4811 15068 4820
rect 15016 4777 15025 4811
rect 15025 4777 15059 4811
rect 15059 4777 15068 4811
rect 15016 4768 15068 4777
rect 15568 4811 15620 4820
rect 15568 4777 15577 4811
rect 15577 4777 15611 4811
rect 15611 4777 15620 4811
rect 15568 4768 15620 4777
rect 15936 4768 15988 4820
rect 16580 4768 16632 4820
rect 16764 4768 16816 4820
rect 18144 4768 18196 4820
rect 20260 4811 20312 4820
rect 20260 4777 20269 4811
rect 20269 4777 20303 4811
rect 20303 4777 20312 4811
rect 20260 4768 20312 4777
rect 20628 4768 20680 4820
rect 5632 4700 5684 4752
rect 7104 4700 7156 4752
rect 8208 4700 8260 4752
rect 12900 4700 12952 4752
rect 13636 4700 13688 4752
rect 7196 4632 7248 4684
rect 1676 4564 1728 4616
rect 3700 4564 3752 4616
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 4344 4607 4396 4616
rect 4344 4573 4353 4607
rect 4353 4573 4387 4607
rect 4387 4573 4396 4607
rect 4344 4564 4396 4573
rect 4620 4564 4672 4616
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 6920 4607 6972 4616
rect 6920 4573 6929 4607
rect 6929 4573 6963 4607
rect 6963 4573 6972 4607
rect 6920 4564 6972 4573
rect 7380 4632 7432 4684
rect 8484 4632 8536 4684
rect 9312 4632 9364 4684
rect 10140 4632 10192 4684
rect 2136 4539 2188 4548
rect 2136 4505 2145 4539
rect 2145 4505 2179 4539
rect 2179 4505 2188 4539
rect 2136 4496 2188 4505
rect 2780 4496 2832 4548
rect 3516 4496 3568 4548
rect 4068 4539 4120 4548
rect 4068 4505 4077 4539
rect 4077 4505 4111 4539
rect 4111 4505 4120 4539
rect 4068 4496 4120 4505
rect 4436 4539 4488 4548
rect 4436 4505 4445 4539
rect 4445 4505 4479 4539
rect 4479 4505 4488 4539
rect 4436 4496 4488 4505
rect 5264 4539 5316 4548
rect 5264 4505 5273 4539
rect 5273 4505 5307 4539
rect 5307 4505 5316 4539
rect 5264 4496 5316 4505
rect 6276 4539 6328 4548
rect 6276 4505 6285 4539
rect 6285 4505 6319 4539
rect 6319 4505 6328 4539
rect 6276 4496 6328 4505
rect 4528 4428 4580 4480
rect 4988 4428 5040 4480
rect 7472 4607 7524 4616
rect 7472 4573 7481 4607
rect 7481 4573 7515 4607
rect 7515 4573 7524 4607
rect 7472 4564 7524 4573
rect 8116 4607 8168 4616
rect 8116 4573 8125 4607
rect 8125 4573 8159 4607
rect 8159 4573 8168 4607
rect 8116 4564 8168 4573
rect 10232 4564 10284 4616
rect 12256 4607 12308 4616
rect 12256 4573 12265 4607
rect 12265 4573 12299 4607
rect 12299 4573 12308 4607
rect 12256 4564 12308 4573
rect 12716 4564 12768 4616
rect 14556 4607 14608 4616
rect 14556 4573 14565 4607
rect 14565 4573 14599 4607
rect 14599 4573 14608 4607
rect 14556 4564 14608 4573
rect 14740 4564 14792 4616
rect 18420 4700 18472 4752
rect 7196 4428 7248 4480
rect 9036 4428 9088 4480
rect 9956 4539 10008 4548
rect 9956 4505 9965 4539
rect 9965 4505 9999 4539
rect 9999 4505 10008 4539
rect 9956 4496 10008 4505
rect 11336 4496 11388 4548
rect 16488 4632 16540 4684
rect 16580 4632 16632 4684
rect 15936 4607 15988 4616
rect 15936 4573 15945 4607
rect 15945 4573 15979 4607
rect 15979 4573 15988 4607
rect 15936 4564 15988 4573
rect 16028 4564 16080 4616
rect 17868 4607 17920 4616
rect 17868 4573 17877 4607
rect 17877 4573 17911 4607
rect 17911 4573 17920 4607
rect 17868 4564 17920 4573
rect 21456 4632 21508 4684
rect 22284 4564 22336 4616
rect 22744 4607 22796 4616
rect 22744 4573 22753 4607
rect 22753 4573 22787 4607
rect 22787 4573 22796 4607
rect 22744 4564 22796 4573
rect 22928 4607 22980 4616
rect 22928 4573 22937 4607
rect 22937 4573 22971 4607
rect 22971 4573 22980 4607
rect 22928 4564 22980 4573
rect 16120 4496 16172 4548
rect 10048 4428 10100 4480
rect 10784 4428 10836 4480
rect 11060 4428 11112 4480
rect 12164 4428 12216 4480
rect 14556 4428 14608 4480
rect 16488 4428 16540 4480
rect 17224 4428 17276 4480
rect 6630 4326 6682 4378
rect 6694 4326 6746 4378
rect 6758 4326 6810 4378
rect 6822 4326 6874 4378
rect 6886 4326 6938 4378
rect 12311 4326 12363 4378
rect 12375 4326 12427 4378
rect 12439 4326 12491 4378
rect 12503 4326 12555 4378
rect 12567 4326 12619 4378
rect 17992 4326 18044 4378
rect 18056 4326 18108 4378
rect 18120 4326 18172 4378
rect 18184 4326 18236 4378
rect 18248 4326 18300 4378
rect 23673 4326 23725 4378
rect 23737 4326 23789 4378
rect 23801 4326 23853 4378
rect 23865 4326 23917 4378
rect 23929 4326 23981 4378
rect 2228 4224 2280 4276
rect 3056 4224 3108 4276
rect 4252 4224 4304 4276
rect 5264 4224 5316 4276
rect 6092 4224 6144 4276
rect 7104 4224 7156 4276
rect 8116 4224 8168 4276
rect 13452 4224 13504 4276
rect 13544 4224 13596 4276
rect 17960 4267 18012 4276
rect 3700 4199 3752 4208
rect 3700 4165 3709 4199
rect 3709 4165 3743 4199
rect 3743 4165 3752 4199
rect 3700 4156 3752 4165
rect 4068 4156 4120 4208
rect 1952 4131 2004 4140
rect 1952 4097 1961 4131
rect 1961 4097 1995 4131
rect 1995 4097 2004 4131
rect 1952 4088 2004 4097
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 2504 4088 2556 4140
rect 2596 4020 2648 4072
rect 3884 4131 3936 4140
rect 3884 4097 3893 4131
rect 3893 4097 3927 4131
rect 3927 4097 3936 4131
rect 3884 4088 3936 4097
rect 3700 4020 3752 4072
rect 4528 4088 4580 4140
rect 5540 4156 5592 4208
rect 7012 4156 7064 4208
rect 14740 4156 14792 4208
rect 17960 4233 17969 4267
rect 17969 4233 18003 4267
rect 18003 4233 18012 4267
rect 17960 4224 18012 4233
rect 22652 4267 22704 4276
rect 22652 4233 22661 4267
rect 22661 4233 22695 4267
rect 22695 4233 22704 4267
rect 22652 4224 22704 4233
rect 15384 4156 15436 4208
rect 4160 4020 4212 4072
rect 5264 4088 5316 4140
rect 4896 4063 4948 4072
rect 4896 4029 4905 4063
rect 4905 4029 4939 4063
rect 4939 4029 4948 4063
rect 4896 4020 4948 4029
rect 2044 3952 2096 4004
rect 2872 3952 2924 4004
rect 3608 3952 3660 4004
rect 3884 3952 3936 4004
rect 2320 3884 2372 3936
rect 4252 3884 4304 3936
rect 4620 3952 4672 4004
rect 6460 4088 6512 4140
rect 7840 4088 7892 4140
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 8760 4131 8812 4140
rect 8760 4097 8769 4131
rect 8769 4097 8803 4131
rect 8803 4097 8812 4131
rect 8760 4088 8812 4097
rect 7196 4063 7248 4072
rect 7196 4029 7205 4063
rect 7205 4029 7239 4063
rect 7239 4029 7248 4063
rect 7196 4020 7248 4029
rect 7932 4020 7984 4072
rect 9220 4131 9272 4140
rect 9220 4097 9229 4131
rect 9229 4097 9263 4131
rect 9263 4097 9272 4131
rect 9220 4088 9272 4097
rect 14556 4088 14608 4140
rect 15844 4088 15896 4140
rect 18696 4156 18748 4208
rect 16120 4134 16172 4143
rect 16120 4100 16129 4134
rect 16129 4100 16163 4134
rect 16163 4100 16172 4134
rect 16120 4091 16172 4100
rect 9128 4020 9180 4072
rect 11612 4020 11664 4072
rect 7472 3952 7524 4004
rect 8484 3952 8536 4004
rect 12164 3952 12216 4004
rect 13728 3952 13780 4004
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 17316 4088 17368 4140
rect 17960 4020 18012 4072
rect 18880 4020 18932 4072
rect 19248 4088 19300 4140
rect 19524 4131 19576 4140
rect 19524 4097 19533 4131
rect 19533 4097 19567 4131
rect 19567 4097 19576 4131
rect 19524 4088 19576 4097
rect 19800 4131 19852 4140
rect 19800 4097 19809 4131
rect 19809 4097 19843 4131
rect 19843 4097 19852 4131
rect 19800 4088 19852 4097
rect 22928 4156 22980 4208
rect 22744 4131 22796 4140
rect 22744 4097 22753 4131
rect 22753 4097 22787 4131
rect 22787 4097 22796 4131
rect 22744 4088 22796 4097
rect 7104 3884 7156 3936
rect 8392 3884 8444 3936
rect 8852 3927 8904 3936
rect 8852 3893 8861 3927
rect 8861 3893 8895 3927
rect 8895 3893 8904 3927
rect 8852 3884 8904 3893
rect 9864 3884 9916 3936
rect 10324 3927 10376 3936
rect 10324 3893 10333 3927
rect 10333 3893 10367 3927
rect 10367 3893 10376 3927
rect 10324 3884 10376 3893
rect 10416 3884 10468 3936
rect 11704 3927 11756 3936
rect 11704 3893 11713 3927
rect 11713 3893 11747 3927
rect 11747 3893 11756 3927
rect 11704 3884 11756 3893
rect 11796 3884 11848 3936
rect 15660 3927 15712 3936
rect 15660 3893 15669 3927
rect 15669 3893 15703 3927
rect 15703 3893 15712 3927
rect 15660 3884 15712 3893
rect 17316 3884 17368 3936
rect 3790 3782 3842 3834
rect 3854 3782 3906 3834
rect 3918 3782 3970 3834
rect 3982 3782 4034 3834
rect 4046 3782 4098 3834
rect 9471 3782 9523 3834
rect 9535 3782 9587 3834
rect 9599 3782 9651 3834
rect 9663 3782 9715 3834
rect 9727 3782 9779 3834
rect 15152 3782 15204 3834
rect 15216 3782 15268 3834
rect 15280 3782 15332 3834
rect 15344 3782 15396 3834
rect 15408 3782 15460 3834
rect 20833 3782 20885 3834
rect 20897 3782 20949 3834
rect 20961 3782 21013 3834
rect 21025 3782 21077 3834
rect 21089 3782 21141 3834
rect 2504 3723 2556 3732
rect 2504 3689 2513 3723
rect 2513 3689 2547 3723
rect 2547 3689 2556 3723
rect 2504 3680 2556 3689
rect 2872 3612 2924 3664
rect 2964 3612 3016 3664
rect 2596 3587 2648 3596
rect 2596 3553 2605 3587
rect 2605 3553 2639 3587
rect 2639 3553 2648 3587
rect 2596 3544 2648 3553
rect 4436 3680 4488 3732
rect 8576 3723 8628 3732
rect 8576 3689 8585 3723
rect 8585 3689 8619 3723
rect 8619 3689 8628 3723
rect 8576 3680 8628 3689
rect 10784 3680 10836 3732
rect 12808 3680 12860 3732
rect 14832 3680 14884 3732
rect 17592 3680 17644 3732
rect 17776 3680 17828 3732
rect 17960 3723 18012 3732
rect 17960 3689 17969 3723
rect 17969 3689 18003 3723
rect 18003 3689 18012 3723
rect 17960 3680 18012 3689
rect 8208 3612 8260 3664
rect 9956 3612 10008 3664
rect 11888 3612 11940 3664
rect 2504 3476 2556 3528
rect 3516 3544 3568 3596
rect 4712 3544 4764 3596
rect 3056 3476 3108 3528
rect 3240 3408 3292 3460
rect 2228 3340 2280 3392
rect 4804 3476 4856 3528
rect 5724 3544 5776 3596
rect 5816 3544 5868 3596
rect 10508 3544 10560 3596
rect 12716 3544 12768 3596
rect 4068 3408 4120 3460
rect 4252 3408 4304 3460
rect 5264 3519 5316 3528
rect 5264 3485 5273 3519
rect 5273 3485 5307 3519
rect 5307 3485 5316 3519
rect 5264 3476 5316 3485
rect 6276 3476 6328 3528
rect 6552 3519 6604 3528
rect 6552 3485 6561 3519
rect 6561 3485 6595 3519
rect 6595 3485 6604 3519
rect 6552 3476 6604 3485
rect 7840 3519 7892 3528
rect 7840 3485 7849 3519
rect 7849 3485 7883 3519
rect 7883 3485 7892 3519
rect 7840 3476 7892 3485
rect 8116 3476 8168 3528
rect 9220 3476 9272 3528
rect 9956 3519 10008 3528
rect 9956 3485 9965 3519
rect 9965 3485 9999 3519
rect 9999 3485 10008 3519
rect 9956 3476 10008 3485
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 11060 3519 11112 3528
rect 11060 3485 11069 3519
rect 11069 3485 11103 3519
rect 11103 3485 11112 3519
rect 11060 3476 11112 3485
rect 4620 3340 4672 3392
rect 5080 3408 5132 3460
rect 5632 3340 5684 3392
rect 6184 3408 6236 3460
rect 8300 3408 8352 3460
rect 11152 3408 11204 3460
rect 11428 3451 11480 3460
rect 11428 3417 11437 3451
rect 11437 3417 11471 3451
rect 11471 3417 11480 3451
rect 11428 3408 11480 3417
rect 12900 3519 12952 3528
rect 12900 3485 12909 3519
rect 12909 3485 12943 3519
rect 12943 3485 12952 3519
rect 12900 3476 12952 3485
rect 17868 3612 17920 3664
rect 14372 3544 14424 3596
rect 20076 3587 20128 3596
rect 20076 3553 20085 3587
rect 20085 3553 20119 3587
rect 20119 3553 20128 3587
rect 20076 3544 20128 3553
rect 23388 3544 23440 3596
rect 14280 3519 14332 3528
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14280 3476 14332 3485
rect 15016 3476 15068 3528
rect 15660 3476 15712 3528
rect 18420 3476 18472 3528
rect 22744 3476 22796 3528
rect 15200 3408 15252 3460
rect 16028 3408 16080 3460
rect 8116 3340 8168 3392
rect 8944 3340 8996 3392
rect 10140 3340 10192 3392
rect 11244 3340 11296 3392
rect 11336 3383 11388 3392
rect 11336 3349 11345 3383
rect 11345 3349 11379 3383
rect 11379 3349 11388 3383
rect 11336 3340 11388 3349
rect 11520 3340 11572 3392
rect 13268 3340 13320 3392
rect 15476 3340 15528 3392
rect 15568 3340 15620 3392
rect 15844 3340 15896 3392
rect 16764 3340 16816 3392
rect 17408 3383 17460 3392
rect 17408 3349 17417 3383
rect 17417 3349 17451 3383
rect 17451 3349 17460 3383
rect 17408 3340 17460 3349
rect 18880 3340 18932 3392
rect 19984 3383 20036 3392
rect 19984 3349 19993 3383
rect 19993 3349 20027 3383
rect 20027 3349 20036 3383
rect 19984 3340 20036 3349
rect 20628 3383 20680 3392
rect 20628 3349 20637 3383
rect 20637 3349 20671 3383
rect 20671 3349 20680 3383
rect 20628 3340 20680 3349
rect 6630 3238 6682 3290
rect 6694 3238 6746 3290
rect 6758 3238 6810 3290
rect 6822 3238 6874 3290
rect 6886 3238 6938 3290
rect 12311 3238 12363 3290
rect 12375 3238 12427 3290
rect 12439 3238 12491 3290
rect 12503 3238 12555 3290
rect 12567 3238 12619 3290
rect 17992 3238 18044 3290
rect 18056 3238 18108 3290
rect 18120 3238 18172 3290
rect 18184 3238 18236 3290
rect 18248 3238 18300 3290
rect 23673 3238 23725 3290
rect 23737 3238 23789 3290
rect 23801 3238 23853 3290
rect 23865 3238 23917 3290
rect 23929 3238 23981 3290
rect 2228 3043 2280 3052
rect 2228 3009 2237 3043
rect 2237 3009 2271 3043
rect 2271 3009 2280 3043
rect 2228 3000 2280 3009
rect 2320 3000 2372 3052
rect 2964 3136 3016 3188
rect 5448 3179 5500 3188
rect 5448 3145 5457 3179
rect 5457 3145 5491 3179
rect 5491 3145 5500 3179
rect 5448 3136 5500 3145
rect 5724 3136 5776 3188
rect 6552 3136 6604 3188
rect 8116 3136 8168 3188
rect 9128 3136 9180 3188
rect 11520 3136 11572 3188
rect 11888 3179 11940 3188
rect 11888 3145 11897 3179
rect 11897 3145 11931 3179
rect 11931 3145 11940 3179
rect 11888 3136 11940 3145
rect 12716 3136 12768 3188
rect 16120 3136 16172 3188
rect 17408 3136 17460 3188
rect 2596 3068 2648 3120
rect 2688 3068 2740 3120
rect 3700 3068 3752 3120
rect 2596 2975 2648 2984
rect 2596 2941 2605 2975
rect 2605 2941 2639 2975
rect 2639 2941 2648 2975
rect 2596 2932 2648 2941
rect 4160 3000 4212 3052
rect 4620 3000 4672 3052
rect 5908 3068 5960 3120
rect 6276 3068 6328 3120
rect 5448 3000 5500 3052
rect 5724 3000 5776 3052
rect 6184 3000 6236 3052
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 4712 2932 4764 2984
rect 1860 2864 1912 2916
rect 2688 2864 2740 2916
rect 2964 2907 3016 2916
rect 2964 2873 2973 2907
rect 2973 2873 3007 2907
rect 3007 2873 3016 2907
rect 2964 2864 3016 2873
rect 4528 2864 4580 2916
rect 6552 2864 6604 2916
rect 4896 2796 4948 2848
rect 7932 3000 7984 3052
rect 8484 3000 8536 3052
rect 8944 3000 8996 3052
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 10140 3111 10192 3120
rect 10140 3077 10149 3111
rect 10149 3077 10183 3111
rect 10183 3077 10192 3111
rect 10140 3068 10192 3077
rect 10508 3068 10560 3120
rect 15568 3068 15620 3120
rect 11336 3000 11388 3052
rect 11612 3000 11664 3052
rect 13268 3043 13320 3052
rect 13268 3009 13277 3043
rect 13277 3009 13311 3043
rect 13311 3009 13320 3043
rect 13268 3000 13320 3009
rect 13452 3043 13504 3052
rect 13452 3009 13461 3043
rect 13461 3009 13495 3043
rect 13495 3009 13504 3043
rect 13452 3000 13504 3009
rect 13728 3000 13780 3052
rect 7472 2975 7524 2984
rect 7472 2941 7481 2975
rect 7481 2941 7515 2975
rect 7515 2941 7524 2975
rect 7472 2932 7524 2941
rect 8116 2975 8168 2984
rect 8116 2941 8125 2975
rect 8125 2941 8159 2975
rect 8159 2941 8168 2975
rect 8116 2932 8168 2941
rect 11060 2932 11112 2984
rect 11152 2932 11204 2984
rect 12164 2975 12216 2984
rect 12164 2941 12173 2975
rect 12173 2941 12207 2975
rect 12207 2941 12216 2975
rect 12164 2932 12216 2941
rect 14280 3000 14332 3052
rect 14556 3043 14608 3052
rect 14556 3009 14565 3043
rect 14565 3009 14599 3043
rect 14599 3009 14608 3043
rect 14556 3000 14608 3009
rect 14924 3043 14976 3052
rect 14924 3009 14933 3043
rect 14933 3009 14967 3043
rect 14967 3009 14976 3043
rect 14924 3000 14976 3009
rect 15936 3068 15988 3120
rect 15844 3043 15896 3052
rect 15844 3009 15853 3043
rect 15853 3009 15887 3043
rect 15887 3009 15896 3043
rect 15844 3000 15896 3009
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 15200 2932 15252 2984
rect 15568 2932 15620 2984
rect 17224 3043 17276 3052
rect 17224 3009 17233 3043
rect 17233 3009 17267 3043
rect 17267 3009 17276 3043
rect 17224 3000 17276 3009
rect 17316 3043 17368 3052
rect 17316 3009 17351 3043
rect 17351 3009 17368 3043
rect 17316 3000 17368 3009
rect 17500 3043 17552 3052
rect 17500 3009 17509 3043
rect 17509 3009 17543 3043
rect 17543 3009 17552 3043
rect 17500 3000 17552 3009
rect 17592 3000 17644 3052
rect 18880 3000 18932 3052
rect 19248 3043 19300 3052
rect 19248 3009 19257 3043
rect 19257 3009 19291 3043
rect 19291 3009 19300 3043
rect 19248 3000 19300 3009
rect 19524 3068 19576 3120
rect 19984 3136 20036 3188
rect 20628 3111 20680 3120
rect 20628 3077 20637 3111
rect 20637 3077 20671 3111
rect 20671 3077 20680 3111
rect 20628 3068 20680 3077
rect 19800 3043 19852 3052
rect 19800 3009 19809 3043
rect 19809 3009 19843 3043
rect 19843 3009 19852 3043
rect 19800 3000 19852 3009
rect 17868 2932 17920 2984
rect 8392 2864 8444 2916
rect 17132 2864 17184 2916
rect 8116 2796 8168 2848
rect 8576 2796 8628 2848
rect 9312 2796 9364 2848
rect 10508 2796 10560 2848
rect 10784 2796 10836 2848
rect 17408 2796 17460 2848
rect 17776 2796 17828 2848
rect 19524 2864 19576 2916
rect 21456 2796 21508 2848
rect 22100 2796 22152 2848
rect 3790 2694 3842 2746
rect 3854 2694 3906 2746
rect 3918 2694 3970 2746
rect 3982 2694 4034 2746
rect 4046 2694 4098 2746
rect 9471 2694 9523 2746
rect 9535 2694 9587 2746
rect 9599 2694 9651 2746
rect 9663 2694 9715 2746
rect 9727 2694 9779 2746
rect 15152 2694 15204 2746
rect 15216 2694 15268 2746
rect 15280 2694 15332 2746
rect 15344 2694 15396 2746
rect 15408 2694 15460 2746
rect 20833 2694 20885 2746
rect 20897 2694 20949 2746
rect 20961 2694 21013 2746
rect 21025 2694 21077 2746
rect 21089 2694 21141 2746
rect 5724 2592 5776 2644
rect 8852 2592 8904 2644
rect 9128 2635 9180 2644
rect 9128 2601 9137 2635
rect 9137 2601 9171 2635
rect 9171 2601 9180 2635
rect 9128 2592 9180 2601
rect 12900 2592 12952 2644
rect 15752 2592 15804 2644
rect 17040 2592 17092 2644
rect 4528 2567 4580 2576
rect 4528 2533 4537 2567
rect 4537 2533 4571 2567
rect 4571 2533 4580 2567
rect 4528 2524 4580 2533
rect 4620 2567 4672 2576
rect 4620 2533 4629 2567
rect 4629 2533 4663 2567
rect 4663 2533 4672 2567
rect 4620 2524 4672 2533
rect 15476 2567 15528 2576
rect 15476 2533 15485 2567
rect 15485 2533 15519 2567
rect 15519 2533 15528 2567
rect 15476 2524 15528 2533
rect 3148 2456 3200 2508
rect 5264 2456 5316 2508
rect 8024 2456 8076 2508
rect 8116 2499 8168 2508
rect 8116 2465 8125 2499
rect 8125 2465 8159 2499
rect 8159 2465 8168 2499
rect 8116 2456 8168 2465
rect 10692 2456 10744 2508
rect 11796 2456 11848 2508
rect 14648 2456 14700 2508
rect 16580 2456 16632 2508
rect 3424 2431 3476 2440
rect 3424 2397 3433 2431
rect 3433 2397 3467 2431
rect 3467 2397 3476 2431
rect 3424 2388 3476 2397
rect 3700 2388 3752 2440
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 5908 2431 5960 2440
rect 5908 2397 5917 2431
rect 5917 2397 5951 2431
rect 5951 2397 5960 2431
rect 5908 2388 5960 2397
rect 7104 2388 7156 2440
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 10968 2388 11020 2440
rect 11428 2388 11480 2440
rect 11980 2388 12032 2440
rect 12716 2388 12768 2440
rect 13084 2388 13136 2440
rect 13820 2388 13872 2440
rect 15568 2388 15620 2440
rect 17132 2431 17184 2440
rect 17132 2397 17141 2431
rect 17141 2397 17175 2431
rect 17175 2397 17184 2431
rect 17132 2388 17184 2397
rect 17408 2431 17460 2440
rect 17408 2397 17417 2431
rect 17417 2397 17451 2431
rect 17451 2397 17460 2431
rect 17408 2388 17460 2397
rect 18512 2431 18564 2440
rect 18512 2397 18521 2431
rect 18521 2397 18555 2431
rect 18555 2397 18564 2431
rect 18512 2388 18564 2397
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 20720 2431 20772 2440
rect 20720 2397 20729 2431
rect 20729 2397 20763 2431
rect 20763 2397 20772 2431
rect 20720 2388 20772 2397
rect 22008 2431 22060 2440
rect 22008 2397 22017 2431
rect 22017 2397 22051 2431
rect 22051 2397 22060 2431
rect 22008 2388 22060 2397
rect 22652 2431 22704 2440
rect 22652 2397 22661 2431
rect 22661 2397 22695 2431
rect 22695 2397 22704 2431
rect 22652 2388 22704 2397
rect 3148 2363 3200 2372
rect 3148 2329 3157 2363
rect 3157 2329 3191 2363
rect 3191 2329 3200 2363
rect 3148 2320 3200 2329
rect 5540 2320 5592 2372
rect 6000 2320 6052 2372
rect 16764 2320 16816 2372
rect 3424 2252 3476 2304
rect 6630 2150 6682 2202
rect 6694 2150 6746 2202
rect 6758 2150 6810 2202
rect 6822 2150 6874 2202
rect 6886 2150 6938 2202
rect 12311 2150 12363 2202
rect 12375 2150 12427 2202
rect 12439 2150 12491 2202
rect 12503 2150 12555 2202
rect 12567 2150 12619 2202
rect 17992 2150 18044 2202
rect 18056 2150 18108 2202
rect 18120 2150 18172 2202
rect 18184 2150 18236 2202
rect 18248 2150 18300 2202
rect 23673 2150 23725 2202
rect 23737 2150 23789 2202
rect 23801 2150 23853 2202
rect 23865 2150 23917 2202
rect 23929 2150 23981 2202
rect 7288 1028 7340 1080
rect 10416 1028 10468 1080
rect 16948 1028 17000 1080
rect 18512 1028 18564 1080
rect 18880 1028 18932 1080
rect 20720 1028 20772 1080
rect 1492 960 1544 1012
rect 5816 960 5868 1012
rect 7932 960 7984 1012
rect 10324 960 10376 1012
rect 18236 960 18288 1012
rect 20076 960 20128 1012
rect 20812 960 20864 1012
rect 22652 960 22704 1012
rect 3148 892 3200 944
rect 4712 892 4764 944
rect 8576 892 8628 944
rect 9772 892 9824 944
rect 17592 892 17644 944
rect 19432 892 19484 944
rect 20168 892 20220 944
rect 22008 892 22060 944
<< metal2 >>
rect 2502 24200 2558 25000
rect 7470 24200 7526 25000
rect 12438 24200 12494 25000
rect 17406 24200 17462 25000
rect 22374 24200 22430 25000
rect 2044 22024 2096 22030
rect 2044 21966 2096 21972
rect 2056 20942 2084 21966
rect 2516 20942 2544 24200
rect 3790 22332 4098 22341
rect 3790 22330 3796 22332
rect 3852 22330 3876 22332
rect 3932 22330 3956 22332
rect 4012 22330 4036 22332
rect 4092 22330 4098 22332
rect 3852 22278 3854 22330
rect 4034 22278 4036 22330
rect 3790 22276 3796 22278
rect 3852 22276 3876 22278
rect 3932 22276 3956 22278
rect 4012 22276 4036 22278
rect 4092 22276 4098 22278
rect 3790 22267 4098 22276
rect 4528 22024 4580 22030
rect 4528 21966 4580 21972
rect 2596 21956 2648 21962
rect 2596 21898 2648 21904
rect 2044 20936 2096 20942
rect 2044 20878 2096 20884
rect 2504 20936 2556 20942
rect 2504 20878 2556 20884
rect 2056 20602 2084 20878
rect 2320 20868 2372 20874
rect 2320 20810 2372 20816
rect 2044 20596 2096 20602
rect 2044 20538 2096 20544
rect 2056 18834 2084 20538
rect 2044 18828 2096 18834
rect 2044 18770 2096 18776
rect 2228 17128 2280 17134
rect 2228 17070 2280 17076
rect 1492 16448 1544 16454
rect 1492 16390 1544 16396
rect 1504 9489 1532 16390
rect 2240 15026 2268 17070
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 2228 15020 2280 15026
rect 2228 14962 2280 14968
rect 1872 14414 1900 14962
rect 1860 14408 1912 14414
rect 1860 14350 1912 14356
rect 1676 14272 1728 14278
rect 1676 14214 1728 14220
rect 1688 13326 1716 14214
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1596 10810 1624 11086
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1688 10606 1716 13262
rect 1872 13258 1900 14350
rect 1952 14340 2004 14346
rect 1952 14282 2004 14288
rect 1860 13252 1912 13258
rect 1860 13194 1912 13200
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1780 12442 1808 13126
rect 1964 12442 1992 14282
rect 2056 14074 2084 14962
rect 2240 14414 2268 14962
rect 2332 14618 2360 20810
rect 2412 19712 2464 19718
rect 2412 19654 2464 19660
rect 2424 15502 2452 19654
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2504 15360 2556 15366
rect 2504 15302 2556 15308
rect 2516 15094 2544 15302
rect 2504 15088 2556 15094
rect 2504 15030 2556 15036
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 2044 14068 2096 14074
rect 2044 14010 2096 14016
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 2148 13394 2176 13806
rect 2240 13462 2268 14214
rect 2412 13932 2464 13938
rect 2412 13874 2464 13880
rect 2228 13456 2280 13462
rect 2228 13398 2280 13404
rect 2136 13388 2188 13394
rect 2136 13330 2188 13336
rect 2044 13184 2096 13190
rect 2044 13126 2096 13132
rect 2056 12646 2084 13126
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 2148 12306 2176 13330
rect 1952 12300 2004 12306
rect 1952 12242 2004 12248
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 1860 11824 1912 11830
rect 1860 11766 1912 11772
rect 1872 11150 1900 11766
rect 1964 11354 1992 12242
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1674 9616 1730 9625
rect 1674 9551 1730 9560
rect 1490 9480 1546 9489
rect 1490 9415 1546 9424
rect 1688 9382 1716 9551
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1688 4622 1716 9318
rect 1872 7342 1900 11086
rect 2240 10742 2268 13398
rect 2424 13326 2452 13874
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 2228 10736 2280 10742
rect 2228 10678 2280 10684
rect 2240 9722 2268 10678
rect 2332 10674 2360 13262
rect 2424 12918 2452 13262
rect 2412 12912 2464 12918
rect 2412 12854 2464 12860
rect 2424 12442 2452 12854
rect 2516 12832 2544 15030
rect 2608 12986 2636 21898
rect 3240 21888 3292 21894
rect 3240 21830 3292 21836
rect 2688 20800 2740 20806
rect 2688 20742 2740 20748
rect 2700 14346 2728 20742
rect 2964 19780 3016 19786
rect 2964 19722 3016 19728
rect 2976 15162 3004 19722
rect 3056 18216 3108 18222
rect 3056 18158 3108 18164
rect 3068 17202 3096 18158
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 3068 16522 3096 17138
rect 3056 16516 3108 16522
rect 3056 16458 3108 16464
rect 3068 15910 3096 16458
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 3068 14958 3096 15846
rect 3056 14952 3108 14958
rect 3056 14894 3108 14900
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2688 14340 2740 14346
rect 2688 14282 2740 14288
rect 2884 14074 2912 14350
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2688 12844 2740 12850
rect 2516 12804 2688 12832
rect 2688 12786 2740 12792
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2700 12594 2728 12786
rect 2792 12714 2820 13670
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2412 12436 2464 12442
rect 2412 12378 2464 12384
rect 2516 10742 2544 12582
rect 2608 12442 2636 12582
rect 2700 12566 2820 12594
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 2504 10736 2556 10742
rect 2504 10678 2556 10684
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2332 9994 2360 10610
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2320 9988 2372 9994
rect 2320 9930 2372 9936
rect 2228 9716 2280 9722
rect 2228 9658 2280 9664
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2148 8974 2176 9522
rect 2240 9042 2268 9658
rect 2332 9586 2360 9930
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2424 9042 2452 10542
rect 2516 10198 2544 10678
rect 2608 10470 2636 12378
rect 2792 12170 2820 12566
rect 2780 12164 2832 12170
rect 2780 12106 2832 12112
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2792 11150 2820 11630
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2504 10192 2556 10198
rect 2504 10134 2556 10140
rect 2608 9586 2636 10406
rect 2792 10130 2820 11086
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 2044 8288 2096 8294
rect 2044 8230 2096 8236
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1872 2922 1900 7278
rect 2056 5574 2084 8230
rect 2148 7546 2176 8910
rect 2504 8900 2556 8906
rect 2504 8842 2556 8848
rect 2516 8430 2544 8842
rect 2608 8650 2636 9522
rect 2608 8622 2728 8650
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 2516 7886 2544 8366
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 2320 7472 2372 7478
rect 2320 7414 2372 7420
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2148 6186 2176 6734
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2136 6180 2188 6186
rect 2136 6122 2188 6128
rect 2148 5914 2176 6122
rect 2240 5914 2268 6258
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2228 5908 2280 5914
rect 2228 5850 2280 5856
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 2148 4706 2176 5850
rect 2332 5794 2360 7414
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2424 6322 2452 7142
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2240 5766 2360 5794
rect 2240 5642 2268 5766
rect 2516 5710 2544 7822
rect 2608 7818 2636 8434
rect 2700 8362 2728 8622
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2792 8090 2820 9862
rect 2884 8974 2912 14010
rect 3068 14006 3096 14894
rect 3056 14000 3108 14006
rect 3056 13942 3108 13948
rect 3252 13326 3280 21830
rect 4540 21622 4568 21966
rect 7484 21962 7512 24200
rect 9471 22332 9779 22341
rect 9471 22330 9477 22332
rect 9533 22330 9557 22332
rect 9613 22330 9637 22332
rect 9693 22330 9717 22332
rect 9773 22330 9779 22332
rect 9533 22278 9535 22330
rect 9715 22278 9717 22330
rect 9471 22276 9477 22278
rect 9533 22276 9557 22278
rect 9613 22276 9637 22278
rect 9693 22276 9717 22278
rect 9773 22276 9779 22278
rect 9471 22267 9779 22276
rect 12452 22114 12480 24200
rect 15152 22332 15460 22341
rect 15152 22330 15158 22332
rect 15214 22330 15238 22332
rect 15294 22330 15318 22332
rect 15374 22330 15398 22332
rect 15454 22330 15460 22332
rect 15214 22278 15216 22330
rect 15396 22278 15398 22330
rect 15152 22276 15158 22278
rect 15214 22276 15238 22278
rect 15294 22276 15318 22278
rect 15374 22276 15398 22278
rect 15454 22276 15460 22278
rect 15152 22267 15460 22276
rect 12716 22160 12768 22166
rect 12072 22092 12124 22098
rect 12452 22086 12572 22114
rect 12716 22102 12768 22108
rect 12072 22034 12124 22040
rect 11980 22024 12032 22030
rect 11980 21966 12032 21972
rect 7472 21956 7524 21962
rect 7472 21898 7524 21904
rect 6092 21888 6144 21894
rect 6092 21830 6144 21836
rect 7380 21888 7432 21894
rect 7380 21830 7432 21836
rect 3700 21616 3752 21622
rect 3700 21558 3752 21564
rect 4528 21616 4580 21622
rect 4528 21558 4580 21564
rect 3332 18692 3384 18698
rect 3332 18634 3384 18640
rect 3344 14618 3372 18634
rect 3516 18352 3568 18358
rect 3516 18294 3568 18300
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3240 13320 3292 13326
rect 3068 13280 3240 13308
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2976 12646 3004 12786
rect 3068 12714 3096 13280
rect 3436 13274 3464 16390
rect 3240 13262 3292 13268
rect 3344 13246 3464 13274
rect 3344 12968 3372 13246
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3160 12940 3372 12968
rect 3160 12782 3188 12940
rect 3436 12850 3464 13126
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 3056 12708 3108 12714
rect 3056 12650 3108 12656
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 2964 12164 3016 12170
rect 2964 12106 3016 12112
rect 2976 10810 3004 12106
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2962 10704 3018 10713
rect 3160 10674 3188 12718
rect 3252 12102 3280 12786
rect 3424 12708 3476 12714
rect 3424 12650 3476 12656
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 2962 10639 2964 10648
rect 3016 10639 3018 10648
rect 3148 10668 3200 10674
rect 2964 10610 3016 10616
rect 3148 10610 3200 10616
rect 3252 10198 3280 12038
rect 3240 10192 3292 10198
rect 3240 10134 3292 10140
rect 3252 9586 3280 10134
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2976 8498 3004 9318
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 3068 8294 3096 8774
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 2596 7812 2648 7818
rect 2596 7754 2648 7760
rect 2780 7812 2832 7818
rect 2780 7754 2832 7760
rect 2608 6202 2636 7754
rect 2792 7410 2820 7754
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2792 7002 2820 7346
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 6322 2728 6598
rect 3068 6322 3096 8026
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 3160 6662 3188 7278
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 2608 6174 2728 6202
rect 2700 5846 2728 6174
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2228 5636 2280 5642
rect 2228 5578 2280 5584
rect 2240 5234 2268 5578
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 1964 4678 2176 4706
rect 1964 4146 1992 4678
rect 2136 4548 2188 4554
rect 2136 4490 2188 4496
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 2056 4010 2084 4082
rect 2044 4004 2096 4010
rect 2044 3946 2096 3952
rect 1860 2916 1912 2922
rect 1860 2858 1912 2864
rect 1492 1012 1544 1018
rect 1492 954 1544 960
rect 1504 800 1532 954
rect 2148 800 2176 4490
rect 2240 4282 2268 5170
rect 2228 4276 2280 4282
rect 2228 4218 2280 4224
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2240 3058 2268 3334
rect 2332 3058 2360 3878
rect 2424 3516 2452 5510
rect 2516 5302 2544 5646
rect 2504 5296 2556 5302
rect 2504 5238 2556 5244
rect 2700 5166 2728 5782
rect 2872 5636 2924 5642
rect 2872 5578 2924 5584
rect 2884 5166 2912 5578
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2780 4548 2832 4554
rect 2780 4490 2832 4496
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2516 3738 2544 4082
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2608 3602 2636 4014
rect 2596 3596 2648 3602
rect 2596 3538 2648 3544
rect 2504 3528 2556 3534
rect 2424 3488 2504 3516
rect 2504 3470 2556 3476
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 2516 2972 2544 3470
rect 2608 3126 2636 3538
rect 2596 3120 2648 3126
rect 2596 3062 2648 3068
rect 2688 3120 2740 3126
rect 2688 3062 2740 3068
rect 2596 2984 2648 2990
rect 2516 2944 2596 2972
rect 2596 2926 2648 2932
rect 2700 2922 2728 3062
rect 2688 2916 2740 2922
rect 2688 2858 2740 2864
rect 2792 800 2820 4490
rect 2884 4010 2912 5102
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 2884 3670 2912 3946
rect 2976 3670 3004 6258
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 3068 5846 3096 6122
rect 3056 5840 3108 5846
rect 3056 5782 3108 5788
rect 3056 5704 3108 5710
rect 3054 5672 3056 5681
rect 3108 5672 3110 5681
rect 3054 5607 3110 5616
rect 3160 5234 3188 6598
rect 3252 5574 3280 8366
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3344 5114 3372 9318
rect 3436 7886 3464 12650
rect 3528 11830 3556 18294
rect 3608 16516 3660 16522
rect 3608 16458 3660 16464
rect 3516 11824 3568 11830
rect 3516 11766 3568 11772
rect 3620 9654 3648 16458
rect 3712 13462 3740 21558
rect 6104 21554 6132 21830
rect 6630 21788 6938 21797
rect 6630 21786 6636 21788
rect 6692 21786 6716 21788
rect 6772 21786 6796 21788
rect 6852 21786 6876 21788
rect 6932 21786 6938 21788
rect 6692 21734 6694 21786
rect 6874 21734 6876 21786
rect 6630 21732 6636 21734
rect 6692 21732 6716 21734
rect 6772 21732 6796 21734
rect 6852 21732 6876 21734
rect 6932 21732 6938 21734
rect 6630 21723 6938 21732
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 5724 21548 5776 21554
rect 5724 21490 5776 21496
rect 6092 21548 6144 21554
rect 6092 21490 6144 21496
rect 3790 21244 4098 21253
rect 3790 21242 3796 21244
rect 3852 21242 3876 21244
rect 3932 21242 3956 21244
rect 4012 21242 4036 21244
rect 4092 21242 4098 21244
rect 3852 21190 3854 21242
rect 4034 21190 4036 21242
rect 3790 21188 3796 21190
rect 3852 21188 3876 21190
rect 3932 21188 3956 21190
rect 4012 21188 4036 21190
rect 4092 21188 4098 21190
rect 3790 21179 4098 21188
rect 4172 20602 4200 21490
rect 4436 21344 4488 21350
rect 4436 21286 4488 21292
rect 4620 21344 4672 21350
rect 4620 21286 4672 21292
rect 4160 20596 4212 20602
rect 4160 20538 4212 20544
rect 3790 20156 4098 20165
rect 3790 20154 3796 20156
rect 3852 20154 3876 20156
rect 3932 20154 3956 20156
rect 4012 20154 4036 20156
rect 4092 20154 4098 20156
rect 3852 20102 3854 20154
rect 4034 20102 4036 20154
rect 3790 20100 3796 20102
rect 3852 20100 3876 20102
rect 3932 20100 3956 20102
rect 4012 20100 4036 20102
rect 4092 20100 4098 20102
rect 3790 20091 4098 20100
rect 4172 19922 4200 20538
rect 4344 20460 4396 20466
rect 4344 20402 4396 20408
rect 4160 19916 4212 19922
rect 4160 19858 4212 19864
rect 4172 19378 4200 19858
rect 4356 19378 4384 20402
rect 4160 19372 4212 19378
rect 4160 19314 4212 19320
rect 4344 19372 4396 19378
rect 4344 19314 4396 19320
rect 3790 19068 4098 19077
rect 3790 19066 3796 19068
rect 3852 19066 3876 19068
rect 3932 19066 3956 19068
rect 4012 19066 4036 19068
rect 4092 19066 4098 19068
rect 3852 19014 3854 19066
rect 4034 19014 4036 19066
rect 3790 19012 3796 19014
rect 3852 19012 3876 19014
rect 3932 19012 3956 19014
rect 4012 19012 4036 19014
rect 4092 19012 4098 19014
rect 3790 19003 4098 19012
rect 3790 17980 4098 17989
rect 3790 17978 3796 17980
rect 3852 17978 3876 17980
rect 3932 17978 3956 17980
rect 4012 17978 4036 17980
rect 4092 17978 4098 17980
rect 3852 17926 3854 17978
rect 4034 17926 4036 17978
rect 3790 17924 3796 17926
rect 3852 17924 3876 17926
rect 3932 17924 3956 17926
rect 4012 17924 4036 17926
rect 4092 17924 4098 17926
rect 3790 17915 4098 17924
rect 3790 16892 4098 16901
rect 3790 16890 3796 16892
rect 3852 16890 3876 16892
rect 3932 16890 3956 16892
rect 4012 16890 4036 16892
rect 4092 16890 4098 16892
rect 3852 16838 3854 16890
rect 4034 16838 4036 16890
rect 3790 16836 3796 16838
rect 3852 16836 3876 16838
rect 3932 16836 3956 16838
rect 4012 16836 4036 16838
rect 4092 16836 4098 16838
rect 3790 16827 4098 16836
rect 4356 16182 4384 19314
rect 4344 16176 4396 16182
rect 4344 16118 4396 16124
rect 3790 15804 4098 15813
rect 3790 15802 3796 15804
rect 3852 15802 3876 15804
rect 3932 15802 3956 15804
rect 4012 15802 4036 15804
rect 4092 15802 4098 15804
rect 3852 15750 3854 15802
rect 4034 15750 4036 15802
rect 3790 15748 3796 15750
rect 3852 15748 3876 15750
rect 3932 15748 3956 15750
rect 4012 15748 4036 15750
rect 4092 15748 4098 15750
rect 3790 15739 4098 15748
rect 3790 14716 4098 14725
rect 3790 14714 3796 14716
rect 3852 14714 3876 14716
rect 3932 14714 3956 14716
rect 4012 14714 4036 14716
rect 4092 14714 4098 14716
rect 3852 14662 3854 14714
rect 4034 14662 4036 14714
rect 3790 14660 3796 14662
rect 3852 14660 3876 14662
rect 3932 14660 3956 14662
rect 4012 14660 4036 14662
rect 4092 14660 4098 14662
rect 3790 14651 4098 14660
rect 4344 14340 4396 14346
rect 4344 14282 4396 14288
rect 3976 14272 4028 14278
rect 3976 14214 4028 14220
rect 3988 13938 4016 14214
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 3790 13628 4098 13637
rect 3790 13626 3796 13628
rect 3852 13626 3876 13628
rect 3932 13626 3956 13628
rect 4012 13626 4036 13628
rect 4092 13626 4098 13628
rect 3852 13574 3854 13626
rect 4034 13574 4036 13626
rect 3790 13572 3796 13574
rect 3852 13572 3876 13574
rect 3932 13572 3956 13574
rect 4012 13572 4036 13574
rect 4092 13572 4098 13574
rect 3790 13563 4098 13572
rect 3700 13456 3752 13462
rect 3700 13398 3752 13404
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 3790 12540 4098 12549
rect 3790 12538 3796 12540
rect 3852 12538 3876 12540
rect 3932 12538 3956 12540
rect 4012 12538 4036 12540
rect 4092 12538 4098 12540
rect 3852 12486 3854 12538
rect 4034 12486 4036 12538
rect 3790 12484 3796 12486
rect 3852 12484 3876 12486
rect 3932 12484 3956 12486
rect 4012 12484 4036 12486
rect 4092 12484 4098 12486
rect 3790 12475 4098 12484
rect 3700 12232 3752 12238
rect 3700 12174 3752 12180
rect 3712 11694 3740 12174
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3804 11694 3832 12038
rect 3700 11688 3752 11694
rect 3700 11630 3752 11636
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3712 11218 3740 11494
rect 3790 11452 4098 11461
rect 3790 11450 3796 11452
rect 3852 11450 3876 11452
rect 3932 11450 3956 11452
rect 4012 11450 4036 11452
rect 4092 11450 4098 11452
rect 3852 11398 3854 11450
rect 4034 11398 4036 11450
rect 3790 11396 3796 11398
rect 3852 11396 3876 11398
rect 3932 11396 3956 11398
rect 4012 11396 4036 11398
rect 4092 11396 4098 11398
rect 3790 11387 4098 11396
rect 4172 11286 4200 11630
rect 4160 11280 4212 11286
rect 4160 11222 4212 11228
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3712 10470 3740 11154
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3608 9648 3660 9654
rect 3608 9590 3660 9596
rect 3712 8838 3740 10406
rect 3790 10364 4098 10373
rect 3790 10362 3796 10364
rect 3852 10362 3876 10364
rect 3932 10362 3956 10364
rect 4012 10362 4036 10364
rect 4092 10362 4098 10364
rect 3852 10310 3854 10362
rect 4034 10310 4036 10362
rect 3790 10308 3796 10310
rect 3852 10308 3876 10310
rect 3932 10308 3956 10310
rect 4012 10308 4036 10310
rect 4092 10308 4098 10310
rect 3790 10299 4098 10308
rect 4172 10062 4200 10542
rect 4264 10266 4292 13262
rect 4356 11898 4384 14282
rect 4448 14074 4476 21286
rect 4632 20777 4660 21286
rect 5632 20800 5684 20806
rect 4618 20768 4674 20777
rect 5632 20742 5684 20748
rect 4618 20703 4674 20712
rect 5356 19712 5408 19718
rect 5356 19654 5408 19660
rect 4620 19440 4672 19446
rect 5368 19417 5396 19654
rect 4620 19382 4672 19388
rect 5354 19408 5410 19417
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4540 15502 4568 16934
rect 4528 15496 4580 15502
rect 4528 15438 4580 15444
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4540 12306 4568 14214
rect 4632 13802 4660 19382
rect 5354 19343 5410 19352
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4620 13796 4672 13802
rect 4620 13738 4672 13744
rect 4816 13462 4844 14010
rect 4804 13456 4856 13462
rect 4804 13398 4856 13404
rect 4816 12442 4844 13398
rect 4896 13320 4948 13326
rect 4894 13288 4896 13297
rect 4948 13288 4950 13297
rect 4894 13223 4950 13232
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 4528 12300 4580 12306
rect 4528 12242 4580 12248
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 4448 11218 4476 12174
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 4448 10742 4476 11154
rect 4540 11150 4568 12242
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4436 10736 4488 10742
rect 4436 10678 4488 10684
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4448 10130 4476 10678
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4080 9722 4108 9998
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 4172 9450 4200 9998
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 3790 9276 4098 9285
rect 3790 9274 3796 9276
rect 3852 9274 3876 9276
rect 3932 9274 3956 9276
rect 4012 9274 4036 9276
rect 4092 9274 4098 9276
rect 3852 9222 3854 9274
rect 4034 9222 4036 9274
rect 3790 9220 3796 9222
rect 3852 9220 3876 9222
rect 3932 9220 3956 9222
rect 4012 9220 4036 9222
rect 4092 9220 4098 9222
rect 3790 9211 4098 9220
rect 4172 8906 4200 9386
rect 4540 9110 4568 11086
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4632 9674 4660 9998
rect 4632 9646 4752 9674
rect 4724 9586 4752 9646
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4528 9104 4580 9110
rect 4528 9046 4580 9052
rect 4160 8900 4212 8906
rect 4160 8842 4212 8848
rect 4252 8900 4304 8906
rect 4252 8842 4304 8848
rect 3700 8832 3752 8838
rect 3700 8774 3752 8780
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 4080 8566 4108 8774
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 4172 8294 4200 8842
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3606 5672 3662 5681
rect 3606 5607 3608 5616
rect 3660 5607 3662 5616
rect 3608 5578 3660 5584
rect 3712 5302 3740 8230
rect 3790 8188 4098 8197
rect 3790 8186 3796 8188
rect 3852 8186 3876 8188
rect 3932 8186 3956 8188
rect 4012 8186 4036 8188
rect 4092 8186 4098 8188
rect 3852 8134 3854 8186
rect 4034 8134 4036 8186
rect 3790 8132 3796 8134
rect 3852 8132 3876 8134
rect 3932 8132 3956 8134
rect 4012 8132 4036 8134
rect 4092 8132 4098 8134
rect 3790 8123 4098 8132
rect 4264 8090 4292 8842
rect 4724 8362 4752 9522
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 4172 7410 4200 7958
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 3790 7100 4098 7109
rect 3790 7098 3796 7100
rect 3852 7098 3876 7100
rect 3932 7098 3956 7100
rect 4012 7098 4036 7100
rect 4092 7098 4098 7100
rect 3852 7046 3854 7098
rect 4034 7046 4036 7098
rect 3790 7044 3796 7046
rect 3852 7044 3876 7046
rect 3932 7044 3956 7046
rect 4012 7044 4036 7046
rect 4092 7044 4098 7046
rect 3790 7035 4098 7044
rect 4264 6746 4292 8026
rect 4540 7886 4568 8298
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4540 7546 4568 7822
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4172 6718 4292 6746
rect 4172 6186 4200 6718
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4160 6180 4212 6186
rect 4160 6122 4212 6128
rect 3790 6012 4098 6021
rect 3790 6010 3796 6012
rect 3852 6010 3876 6012
rect 3932 6010 3956 6012
rect 4012 6010 4036 6012
rect 4092 6010 4098 6012
rect 3852 5958 3854 6010
rect 4034 5958 4036 6010
rect 3790 5956 3796 5958
rect 3852 5956 3876 5958
rect 3932 5956 3956 5958
rect 4012 5956 4036 5958
rect 4092 5956 4098 5958
rect 3790 5947 4098 5956
rect 4172 5710 4200 6122
rect 4264 6118 4292 6598
rect 4344 6384 4396 6390
rect 4344 6326 4396 6332
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 5302 4108 5510
rect 3700 5296 3752 5302
rect 3620 5256 3700 5284
rect 3160 5086 3372 5114
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 2964 3664 3016 3670
rect 2964 3606 3016 3612
rect 2976 3194 3004 3606
rect 3068 3534 3096 4218
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 2962 2952 3018 2961
rect 2962 2887 2964 2896
rect 3016 2887 3018 2896
rect 2964 2858 3016 2864
rect 3160 2514 3188 5086
rect 3528 4554 3556 5102
rect 3516 4548 3568 4554
rect 3516 4490 3568 4496
rect 3620 4128 3648 5256
rect 3700 5238 3752 5244
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 3790 4924 4098 4933
rect 3790 4922 3796 4924
rect 3852 4922 3876 4924
rect 3932 4922 3956 4924
rect 4012 4922 4036 4924
rect 4092 4922 4098 4924
rect 3852 4870 3854 4922
rect 4034 4870 4036 4922
rect 3790 4868 3796 4870
rect 3852 4868 3876 4870
rect 3932 4868 3956 4870
rect 4012 4868 4036 4870
rect 4092 4868 4098 4870
rect 3790 4859 4098 4868
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3712 4214 3740 4558
rect 4068 4548 4120 4554
rect 4068 4490 4120 4496
rect 4080 4214 4108 4490
rect 3700 4208 3752 4214
rect 3700 4150 3752 4156
rect 4068 4208 4120 4214
rect 4068 4150 4120 4156
rect 3528 4100 3648 4128
rect 3884 4140 3936 4146
rect 3528 3602 3556 4100
rect 3884 4082 3936 4088
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 3620 3482 3648 3946
rect 3252 3466 3648 3482
rect 3240 3460 3648 3466
rect 3292 3454 3648 3460
rect 3240 3402 3292 3408
rect 3712 3126 3740 4014
rect 3896 4010 3924 4082
rect 4172 4078 4200 5646
rect 4264 4622 4292 6054
rect 4356 5846 4384 6326
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4448 6118 4476 6258
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4344 5840 4396 5846
rect 4344 5782 4396 5788
rect 4356 4622 4384 5782
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4448 4554 4476 5646
rect 4540 5234 4568 6802
rect 4632 6322 4660 6802
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4632 5370 4660 6258
rect 4724 5710 4752 8298
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4632 4622 4660 5306
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4436 4548 4488 4554
rect 4436 4490 4488 4496
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 3884 4004 3936 4010
rect 3884 3946 3936 3952
rect 4264 3942 4292 4218
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 3790 3836 4098 3845
rect 3790 3834 3796 3836
rect 3852 3834 3876 3836
rect 3932 3834 3956 3836
rect 4012 3834 4036 3836
rect 4092 3834 4098 3836
rect 3852 3782 3854 3834
rect 4034 3782 4036 3834
rect 3790 3780 3796 3782
rect 3852 3780 3876 3782
rect 3932 3780 3956 3782
rect 4012 3780 4036 3782
rect 4092 3780 4098 3782
rect 3790 3771 4098 3780
rect 4448 3738 4476 4490
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4540 4146 4568 4422
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 4252 3460 4304 3466
rect 4252 3402 4304 3408
rect 3700 3120 3752 3126
rect 3700 3062 3752 3068
rect 3422 2544 3478 2553
rect 3148 2508 3200 2514
rect 3422 2479 3478 2488
rect 3148 2450 3200 2456
rect 3436 2446 3464 2479
rect 3712 2446 3740 3062
rect 4080 2904 4108 3402
rect 4160 3052 4212 3058
rect 4264 3040 4292 3402
rect 4632 3398 4660 3946
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4632 3058 4660 3334
rect 4212 3012 4292 3040
rect 4620 3052 4672 3058
rect 4160 2994 4212 3000
rect 4620 2994 4672 3000
rect 4528 2916 4580 2922
rect 4080 2876 4200 2904
rect 3790 2748 4098 2757
rect 3790 2746 3796 2748
rect 3852 2746 3876 2748
rect 3932 2746 3956 2748
rect 4012 2746 4036 2748
rect 4092 2746 4098 2748
rect 3852 2694 3854 2746
rect 4034 2694 4036 2746
rect 3790 2692 3796 2694
rect 3852 2692 3876 2694
rect 3932 2692 3956 2694
rect 4012 2692 4036 2694
rect 4092 2692 4098 2694
rect 3790 2683 4098 2692
rect 4172 2530 4200 2876
rect 4528 2858 4580 2864
rect 4540 2582 4568 2858
rect 4632 2582 4660 2994
rect 4724 2990 4752 3538
rect 4816 3534 4844 11834
rect 5000 10062 5028 15438
rect 5092 11898 5120 18022
rect 5172 15428 5224 15434
rect 5172 15370 5224 15376
rect 5184 14482 5212 15370
rect 5172 14476 5224 14482
rect 5172 14418 5224 14424
rect 5184 13190 5212 14418
rect 5276 14074 5304 19246
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 5460 15094 5488 18566
rect 5448 15088 5500 15094
rect 5448 15030 5500 15036
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5368 14414 5396 14758
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 5184 12918 5212 13126
rect 5172 12912 5224 12918
rect 5172 12854 5224 12860
rect 5264 12640 5316 12646
rect 5368 12628 5396 14350
rect 5448 14340 5500 14346
rect 5448 14282 5500 14288
rect 5460 13530 5488 14282
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5552 13410 5580 13738
rect 5460 13382 5580 13410
rect 5460 12782 5488 13382
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5552 12850 5580 13262
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5316 12600 5396 12628
rect 5264 12582 5316 12588
rect 5644 12442 5672 20742
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 5172 11620 5224 11626
rect 5172 11562 5224 11568
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 4894 9616 4950 9625
rect 4894 9551 4950 9560
rect 4988 9580 5040 9586
rect 4908 9382 4936 9551
rect 4988 9522 5040 9528
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4908 6186 4936 7346
rect 5000 6186 5028 9522
rect 5092 8906 5120 10746
rect 5184 10062 5212 11562
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5184 9178 5212 9998
rect 5276 9674 5304 12378
rect 5448 12096 5500 12102
rect 5446 12064 5448 12073
rect 5500 12064 5502 12073
rect 5446 11999 5502 12008
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5368 10810 5396 11698
rect 5460 11354 5488 11698
rect 5552 11626 5580 11698
rect 5540 11620 5592 11626
rect 5540 11562 5592 11568
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5276 9646 5396 9674
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5080 8900 5132 8906
rect 5080 8842 5132 8848
rect 5092 7886 5120 8842
rect 5184 8566 5212 8978
rect 5276 8906 5304 9522
rect 5368 9382 5396 9646
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 5368 9178 5396 9318
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5460 9024 5488 11086
rect 5552 9654 5580 11562
rect 5632 11280 5684 11286
rect 5632 11222 5684 11228
rect 5644 10674 5672 11222
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5736 10470 5764 21490
rect 7196 21344 7248 21350
rect 7196 21286 7248 21292
rect 7208 20942 7236 21286
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 7196 20936 7248 20942
rect 7196 20878 7248 20884
rect 5828 18970 5856 20878
rect 7104 20868 7156 20874
rect 7104 20810 7156 20816
rect 6630 20700 6938 20709
rect 6630 20698 6636 20700
rect 6692 20698 6716 20700
rect 6772 20698 6796 20700
rect 6852 20698 6876 20700
rect 6932 20698 6938 20700
rect 6692 20646 6694 20698
rect 6874 20646 6876 20698
rect 6630 20644 6636 20646
rect 6692 20644 6716 20646
rect 6772 20644 6796 20646
rect 6852 20644 6876 20646
rect 6932 20644 6938 20646
rect 6630 20635 6938 20644
rect 6184 19780 6236 19786
rect 6184 19722 6236 19728
rect 5816 18964 5868 18970
rect 5816 18906 5868 18912
rect 5828 18766 5856 18906
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 6104 16697 6132 17478
rect 6090 16688 6146 16697
rect 6090 16623 6146 16632
rect 6000 15020 6052 15026
rect 6000 14962 6052 14968
rect 5908 14884 5960 14890
rect 5908 14826 5960 14832
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 5828 14006 5856 14350
rect 5816 14000 5868 14006
rect 5816 13942 5868 13948
rect 5828 13190 5856 13942
rect 5920 13734 5948 14826
rect 5908 13728 5960 13734
rect 5908 13670 5960 13676
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5828 11694 5856 11834
rect 5920 11830 5948 13466
rect 6012 13297 6040 14962
rect 6092 14952 6144 14958
rect 6092 14894 6144 14900
rect 6104 14618 6132 14894
rect 6092 14612 6144 14618
rect 6092 14554 6144 14560
rect 5998 13288 6054 13297
rect 5998 13223 6054 13232
rect 6012 12714 6040 13223
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6104 12986 6132 13126
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6092 12844 6144 12850
rect 6092 12786 6144 12792
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 5908 11824 5960 11830
rect 5908 11766 5960 11772
rect 5816 11688 5868 11694
rect 5816 11630 5868 11636
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5368 8996 5488 9024
rect 5264 8900 5316 8906
rect 5264 8842 5316 8848
rect 5172 8560 5224 8566
rect 5172 8502 5224 8508
rect 5184 8022 5212 8502
rect 5368 8498 5396 8996
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5172 8016 5224 8022
rect 5172 7958 5224 7964
rect 5368 7886 5396 8434
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5368 7478 5396 7686
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5276 6866 5304 7142
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5460 6730 5488 8842
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 5460 6322 5488 6666
rect 5540 6656 5592 6662
rect 5644 6644 5672 10202
rect 5828 10130 5856 10542
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5920 9586 5948 11630
rect 6104 11150 6132 12786
rect 6196 11898 6224 19722
rect 6630 19612 6938 19621
rect 6630 19610 6636 19612
rect 6692 19610 6716 19612
rect 6772 19610 6796 19612
rect 6852 19610 6876 19612
rect 6932 19610 6938 19612
rect 6692 19558 6694 19610
rect 6874 19558 6876 19610
rect 6630 19556 6636 19558
rect 6692 19556 6716 19558
rect 6772 19556 6796 19558
rect 6852 19556 6876 19558
rect 6932 19556 6938 19558
rect 6630 19547 6938 19556
rect 6630 18524 6938 18533
rect 6630 18522 6636 18524
rect 6692 18522 6716 18524
rect 6772 18522 6796 18524
rect 6852 18522 6876 18524
rect 6932 18522 6938 18524
rect 6692 18470 6694 18522
rect 6874 18470 6876 18522
rect 6630 18468 6636 18470
rect 6692 18468 6716 18470
rect 6772 18468 6796 18470
rect 6852 18468 6876 18470
rect 6932 18468 6938 18470
rect 6630 18459 6938 18468
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6564 17134 6592 17614
rect 6630 17436 6938 17445
rect 6630 17434 6636 17436
rect 6692 17434 6716 17436
rect 6772 17434 6796 17436
rect 6852 17434 6876 17436
rect 6932 17434 6938 17436
rect 6692 17382 6694 17434
rect 6874 17382 6876 17434
rect 6630 17380 6636 17382
rect 6692 17380 6716 17382
rect 6772 17380 6796 17382
rect 6852 17380 6876 17382
rect 6932 17380 6938 17382
rect 6630 17371 6938 17380
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6564 16658 6592 17070
rect 6552 16652 6604 16658
rect 7116 16640 7144 20810
rect 7208 19854 7236 20878
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 7116 16612 7236 16640
rect 6552 16594 6604 16600
rect 6276 16516 6328 16522
rect 6276 16458 6328 16464
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6288 11014 6316 16458
rect 6564 15570 6592 16594
rect 6630 16348 6938 16357
rect 6630 16346 6636 16348
rect 6692 16346 6716 16348
rect 6772 16346 6796 16348
rect 6852 16346 6876 16348
rect 6932 16346 6938 16348
rect 6692 16294 6694 16346
rect 6874 16294 6876 16346
rect 6630 16292 6636 16294
rect 6692 16292 6716 16294
rect 6772 16292 6796 16294
rect 6852 16292 6876 16294
rect 6932 16292 6938 16294
rect 6630 16283 6938 16292
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 6630 15260 6938 15269
rect 6630 15258 6636 15260
rect 6692 15258 6716 15260
rect 6772 15258 6796 15260
rect 6852 15258 6876 15260
rect 6932 15258 6938 15260
rect 6692 15206 6694 15258
rect 6874 15206 6876 15258
rect 6630 15204 6636 15206
rect 6692 15204 6716 15206
rect 6772 15204 6796 15206
rect 6852 15204 6876 15206
rect 6932 15204 6938 15206
rect 6630 15195 6938 15204
rect 7012 15088 7064 15094
rect 7012 15030 7064 15036
rect 6644 14884 6696 14890
rect 6644 14826 6696 14832
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6368 14340 6420 14346
rect 6368 14282 6420 14288
rect 6460 14340 6512 14346
rect 6460 14282 6512 14288
rect 6380 11082 6408 14282
rect 6472 14074 6500 14282
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 6460 13728 6512 13734
rect 6460 13670 6512 13676
rect 6472 12850 6500 13670
rect 6564 13326 6592 14758
rect 6656 14414 6684 14826
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6630 14172 6938 14181
rect 6630 14170 6636 14172
rect 6692 14170 6716 14172
rect 6772 14170 6796 14172
rect 6852 14170 6876 14172
rect 6932 14170 6938 14172
rect 6692 14118 6694 14170
rect 6874 14118 6876 14170
rect 6630 14116 6636 14118
rect 6692 14116 6716 14118
rect 6772 14116 6796 14118
rect 6852 14116 6876 14118
rect 6932 14116 6938 14118
rect 6630 14107 6938 14116
rect 7024 13530 7052 15030
rect 7104 14272 7156 14278
rect 7104 14214 7156 14220
rect 7116 13802 7144 14214
rect 7104 13796 7156 13802
rect 7104 13738 7156 13744
rect 7012 13524 7064 13530
rect 7064 13484 7144 13512
rect 7012 13466 7064 13472
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 6630 13084 6938 13093
rect 6630 13082 6636 13084
rect 6692 13082 6716 13084
rect 6772 13082 6796 13084
rect 6852 13082 6876 13084
rect 6932 13082 6938 13084
rect 6692 13030 6694 13082
rect 6874 13030 6876 13082
rect 6630 13028 6636 13030
rect 6692 13028 6716 13030
rect 6772 13028 6796 13030
rect 6852 13028 6876 13030
rect 6932 13028 6938 13030
rect 6630 13019 6938 13028
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6460 12708 6512 12714
rect 6460 12650 6512 12656
rect 6472 12434 6500 12650
rect 6472 12406 6592 12434
rect 6460 11824 6512 11830
rect 6564 11812 6592 12406
rect 6932 12238 6960 12854
rect 7024 12374 7052 13262
rect 7116 12918 7144 13484
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6630 11996 6938 12005
rect 6630 11994 6636 11996
rect 6692 11994 6716 11996
rect 6772 11994 6796 11996
rect 6852 11994 6876 11996
rect 6932 11994 6938 11996
rect 6692 11942 6694 11994
rect 6874 11942 6876 11994
rect 6630 11940 6636 11942
rect 6692 11940 6716 11942
rect 6772 11940 6796 11942
rect 6852 11940 6876 11942
rect 6932 11940 6938 11942
rect 6630 11931 6938 11940
rect 6564 11784 6684 11812
rect 6460 11766 6512 11772
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 6276 11008 6328 11014
rect 6276 10950 6328 10956
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 5724 9512 5776 9518
rect 5722 9480 5724 9489
rect 5776 9480 5778 9489
rect 5722 9415 5778 9424
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5920 7818 5948 8230
rect 5908 7812 5960 7818
rect 5908 7754 5960 7760
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5828 6798 5856 7142
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5736 6662 5764 6734
rect 5592 6616 5672 6644
rect 5724 6656 5776 6662
rect 5540 6598 5592 6604
rect 5920 6610 5948 7754
rect 5724 6598 5776 6604
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 4896 6180 4948 6186
rect 4896 6122 4948 6128
rect 4988 6180 5040 6186
rect 4988 6122 5040 6128
rect 4908 4078 4936 6122
rect 5552 5914 5580 6598
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 5000 5166 5028 5646
rect 5540 5636 5592 5642
rect 5540 5578 5592 5584
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 5000 4486 5028 5102
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4080 2502 4200 2530
rect 4528 2576 4580 2582
rect 4528 2518 4580 2524
rect 4620 2576 4672 2582
rect 4620 2518 4672 2524
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 3700 2440 3752 2446
rect 3700 2382 3752 2388
rect 3148 2372 3200 2378
rect 3148 2314 3200 2320
rect 3160 950 3188 2314
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3148 944 3200 950
rect 3148 886 3200 892
rect 3436 800 3464 2246
rect 4080 800 4108 2502
rect 4724 2446 4752 2926
rect 4908 2854 4936 4014
rect 5092 3466 5120 5170
rect 5552 4622 5580 5578
rect 5736 5574 5764 6598
rect 5828 6582 5948 6610
rect 5828 6118 5856 6582
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5644 4758 5672 5510
rect 5828 5234 5856 6054
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5264 4548 5316 4554
rect 5264 4490 5316 4496
rect 5276 4282 5304 4490
rect 5264 4276 5316 4282
rect 5264 4218 5316 4224
rect 5552 4214 5580 4558
rect 5540 4208 5592 4214
rect 5540 4150 5592 4156
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5276 3534 5304 4082
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5446 3496 5502 3505
rect 5080 3460 5132 3466
rect 5080 3402 5132 3408
rect 4896 2848 4948 2854
rect 4896 2790 4948 2796
rect 5276 2514 5304 3470
rect 5446 3431 5502 3440
rect 5460 3194 5488 3431
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5448 3052 5500 3058
rect 5552 3040 5580 4150
rect 5644 3398 5672 4694
rect 5736 3602 5764 5102
rect 5828 5001 5856 5170
rect 5814 4992 5870 5001
rect 5814 4927 5870 4936
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 5736 3194 5764 3538
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5500 3012 5580 3040
rect 5724 3052 5776 3058
rect 5448 2994 5500 3000
rect 5724 2994 5776 3000
rect 5736 2650 5764 2994
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 5540 2372 5592 2378
rect 5540 2314 5592 2320
rect 4712 944 4764 950
rect 5552 898 5580 2314
rect 5828 1018 5856 3538
rect 5920 3126 5948 6258
rect 5908 3120 5960 3126
rect 5908 3062 5960 3068
rect 6012 2774 6040 10950
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6196 9722 6224 10610
rect 6380 10010 6408 11018
rect 6288 9982 6408 10010
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6196 7818 6224 8978
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6288 7206 6316 9982
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6380 9058 6408 9862
rect 6472 9330 6500 11766
rect 6656 11286 6684 11784
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6748 11098 6776 11698
rect 6932 11626 6960 11698
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6564 11070 6776 11098
rect 6564 10810 6592 11070
rect 6630 10908 6938 10917
rect 6630 10906 6636 10908
rect 6692 10906 6716 10908
rect 6772 10906 6796 10908
rect 6852 10906 6876 10908
rect 6932 10906 6938 10908
rect 6692 10854 6694 10906
rect 6874 10854 6876 10906
rect 6630 10852 6636 10854
rect 6692 10852 6716 10854
rect 6772 10852 6796 10854
rect 6852 10852 6876 10854
rect 6932 10852 6938 10854
rect 6630 10843 6938 10852
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 7024 10742 7052 12310
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 7116 11778 7144 12106
rect 7208 11898 7236 16612
rect 7392 15026 7420 21830
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 8208 21480 8260 21486
rect 8208 21422 8260 21428
rect 8116 21344 8168 21350
rect 8116 21286 8168 21292
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7668 18970 7696 19314
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7668 18290 7696 18906
rect 7656 18284 7708 18290
rect 7656 18226 7708 18232
rect 7472 17604 7524 17610
rect 7472 17546 7524 17552
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7300 13258 7328 14350
rect 7392 14006 7420 14962
rect 7380 14000 7432 14006
rect 7380 13942 7432 13948
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7116 11750 7236 11778
rect 7208 11694 7236 11750
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7300 11626 7328 12378
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 7012 10736 7064 10742
rect 7012 10678 7064 10684
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6564 9625 6592 10066
rect 6630 9820 6938 9829
rect 6630 9818 6636 9820
rect 6692 9818 6716 9820
rect 6772 9818 6796 9820
rect 6852 9818 6876 9820
rect 6932 9818 6938 9820
rect 6692 9766 6694 9818
rect 6874 9766 6876 9818
rect 6630 9764 6636 9766
rect 6692 9764 6716 9766
rect 6772 9764 6796 9766
rect 6852 9764 6876 9766
rect 6932 9764 6938 9766
rect 6630 9755 6938 9764
rect 7024 9722 7052 10542
rect 7116 10062 7144 10610
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 6550 9616 6606 9625
rect 6550 9551 6606 9560
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 6472 9302 6868 9330
rect 6840 9178 6868 9302
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6380 9042 6868 9058
rect 6380 9036 6880 9042
rect 6380 9030 6828 9036
rect 6828 8978 6880 8984
rect 7024 8974 7052 9386
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 6472 8566 6500 8910
rect 6630 8732 6938 8741
rect 6630 8730 6636 8732
rect 6692 8730 6716 8732
rect 6772 8730 6796 8732
rect 6852 8730 6876 8732
rect 6932 8730 6938 8732
rect 6692 8678 6694 8730
rect 6874 8678 6876 8730
rect 6630 8676 6636 8678
rect 6692 8676 6716 8678
rect 6772 8676 6796 8678
rect 6852 8676 6876 8678
rect 6932 8676 6938 8678
rect 6630 8667 6938 8676
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6380 5846 6408 6054
rect 6368 5840 6420 5846
rect 6368 5782 6420 5788
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 6104 5166 6132 5714
rect 6380 5370 6408 5782
rect 6472 5574 6500 8502
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 6564 7410 6592 8366
rect 6828 8356 6880 8362
rect 6880 8316 6960 8344
rect 6828 8298 6880 8304
rect 6932 8022 6960 8316
rect 6920 8016 6972 8022
rect 6920 7958 6972 7964
rect 6932 7886 6960 7958
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6630 7644 6938 7653
rect 6630 7642 6636 7644
rect 6692 7642 6716 7644
rect 6772 7642 6796 7644
rect 6852 7642 6876 7644
rect 6932 7642 6938 7644
rect 6692 7590 6694 7642
rect 6874 7590 6876 7642
rect 6630 7588 6636 7590
rect 6692 7588 6716 7590
rect 6772 7588 6796 7590
rect 6852 7588 6876 7590
rect 6932 7588 6938 7590
rect 6630 7579 6938 7588
rect 7024 7410 7052 8910
rect 7116 8634 7144 9522
rect 7208 9178 7236 10542
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 6564 7206 6592 7346
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6564 5710 6592 7142
rect 6826 6760 6882 6769
rect 6826 6695 6828 6704
rect 6880 6695 6882 6704
rect 6828 6666 6880 6672
rect 6630 6556 6938 6565
rect 6630 6554 6636 6556
rect 6692 6554 6716 6556
rect 6772 6554 6796 6556
rect 6852 6554 6876 6556
rect 6932 6554 6938 6556
rect 6692 6502 6694 6554
rect 6874 6502 6876 6554
rect 6630 6500 6636 6502
rect 6692 6500 6716 6502
rect 6772 6500 6796 6502
rect 6852 6500 6876 6502
rect 6932 6500 6938 6502
rect 6630 6491 6938 6500
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6656 5642 6684 6258
rect 6644 5636 6696 5642
rect 6644 5578 6696 5584
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6828 5568 6880 5574
rect 6880 5528 7052 5556
rect 6828 5510 6880 5516
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 6104 4282 6132 5102
rect 6276 4548 6328 4554
rect 6276 4490 6328 4496
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 6288 3534 6316 4490
rect 6472 4146 6500 5510
rect 6630 5468 6938 5477
rect 6630 5466 6636 5468
rect 6692 5466 6716 5468
rect 6772 5466 6796 5468
rect 6852 5466 6876 5468
rect 6932 5466 6938 5468
rect 6692 5414 6694 5466
rect 6874 5414 6876 5466
rect 6630 5412 6636 5414
rect 6692 5412 6716 5414
rect 6772 5412 6796 5414
rect 6852 5412 6876 5414
rect 6932 5412 6938 5414
rect 6630 5403 6938 5412
rect 7024 5234 7052 5528
rect 7104 5296 7156 5302
rect 7104 5238 7156 5244
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 6642 5128 6698 5137
rect 6642 5063 6698 5072
rect 6920 5092 6972 5098
rect 6656 5030 6684 5063
rect 6920 5034 6972 5040
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6932 4622 6960 5034
rect 7116 4758 7144 5238
rect 7104 4752 7156 4758
rect 7104 4694 7156 4700
rect 6920 4616 6972 4622
rect 6972 4576 7052 4604
rect 6920 4558 6972 4564
rect 6630 4380 6938 4389
rect 6630 4378 6636 4380
rect 6692 4378 6716 4380
rect 6772 4378 6796 4380
rect 6852 4378 6876 4380
rect 6932 4378 6938 4380
rect 6692 4326 6694 4378
rect 6874 4326 6876 4378
rect 6630 4324 6636 4326
rect 6692 4324 6716 4326
rect 6772 4324 6796 4326
rect 6852 4324 6876 4326
rect 6932 4324 6938 4326
rect 6630 4315 6938 4324
rect 7024 4214 7052 4576
rect 7116 4282 7144 4694
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7208 4486 7236 4626
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7012 4208 7064 4214
rect 7300 4162 7328 11562
rect 7392 10266 7420 12174
rect 7484 10538 7512 17546
rect 7668 16182 7696 18226
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7656 16176 7708 16182
rect 7656 16118 7708 16124
rect 7760 14618 7788 16526
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7840 14408 7892 14414
rect 7840 14350 7892 14356
rect 7564 14340 7616 14346
rect 7564 14282 7616 14288
rect 7576 14074 7604 14282
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 7748 14000 7800 14006
rect 7748 13942 7800 13948
rect 7576 13394 7696 13410
rect 7576 13388 7708 13394
rect 7576 13382 7656 13388
rect 7576 12442 7604 13382
rect 7656 13330 7708 13336
rect 7760 13274 7788 13942
rect 7668 13246 7788 13274
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7576 9994 7604 12174
rect 7668 10674 7696 13246
rect 7852 11642 7880 14350
rect 7944 13462 7972 17138
rect 8036 16794 8064 17478
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8036 16590 8064 16730
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 7932 13456 7984 13462
rect 7932 13398 7984 13404
rect 7932 13252 7984 13258
rect 7932 13194 7984 13200
rect 7944 12238 7972 13194
rect 8036 12714 8064 14350
rect 8024 12708 8076 12714
rect 8024 12650 8076 12656
rect 8128 12442 8156 21286
rect 8220 20398 8248 21422
rect 9864 21344 9916 21350
rect 9864 21286 9916 21292
rect 9471 21244 9779 21253
rect 9471 21242 9477 21244
rect 9533 21242 9557 21244
rect 9613 21242 9637 21244
rect 9693 21242 9717 21244
rect 9773 21242 9779 21244
rect 9533 21190 9535 21242
rect 9715 21190 9717 21242
rect 9471 21188 9477 21190
rect 9533 21188 9557 21190
rect 9613 21188 9637 21190
rect 9693 21188 9717 21190
rect 9773 21188 9779 21190
rect 9471 21179 9779 21188
rect 8392 21072 8444 21078
rect 8392 21014 8444 21020
rect 8208 20392 8260 20398
rect 8208 20334 8260 20340
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 8220 19378 8248 19790
rect 8208 19372 8260 19378
rect 8208 19314 8260 19320
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8208 14544 8260 14550
rect 8208 14486 8260 14492
rect 8220 14074 8248 14486
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8220 13326 8248 14010
rect 8312 13938 8340 15438
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8116 12436 8168 12442
rect 8116 12378 8168 12384
rect 8220 12374 8248 13262
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8404 12238 8432 21014
rect 9128 20936 9180 20942
rect 9128 20878 9180 20884
rect 8484 20800 8536 20806
rect 8484 20742 8536 20748
rect 8496 19786 8524 20742
rect 9140 20262 9168 20878
rect 9128 20256 9180 20262
rect 9128 20198 9180 20204
rect 9140 19854 9168 20198
rect 9471 20156 9779 20165
rect 9471 20154 9477 20156
rect 9533 20154 9557 20156
rect 9613 20154 9637 20156
rect 9693 20154 9717 20156
rect 9773 20154 9779 20156
rect 9533 20102 9535 20154
rect 9715 20102 9717 20154
rect 9471 20100 9477 20102
rect 9533 20100 9557 20102
rect 9613 20100 9637 20102
rect 9693 20100 9717 20102
rect 9773 20100 9779 20102
rect 9471 20091 9779 20100
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 8484 19780 8536 19786
rect 8484 19722 8536 19728
rect 9140 18766 9168 19790
rect 9220 19712 9272 19718
rect 9220 19654 9272 19660
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9140 18426 9168 18702
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 8496 16658 8524 17070
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8668 14544 8720 14550
rect 8668 14486 8720 14492
rect 8484 14340 8536 14346
rect 8484 14282 8536 14288
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8496 12170 8524 14282
rect 8680 14278 8708 14486
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 7852 11614 8064 11642
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7564 9988 7616 9994
rect 7564 9930 7616 9936
rect 7380 9580 7432 9586
rect 7432 9540 7512 9568
rect 7380 9522 7432 9528
rect 7484 9500 7512 9540
rect 7656 9512 7708 9518
rect 7484 9472 7656 9500
rect 7656 9454 7708 9460
rect 7668 9042 7696 9454
rect 7944 9382 7972 11290
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7760 8634 7788 9318
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7668 8294 7696 8434
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7392 7818 7420 8026
rect 7760 7886 7788 8230
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7380 7812 7432 7818
rect 7380 7754 7432 7760
rect 7392 6322 7420 7754
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7760 6254 7788 7346
rect 7852 6798 7880 8978
rect 8036 8906 8064 11614
rect 8496 10713 8524 12106
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8482 10704 8538 10713
rect 8482 10639 8538 10648
rect 8496 9722 8524 10639
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 8116 9444 8168 9450
rect 8116 9386 8168 9392
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 8128 8090 8156 9386
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8116 8084 8168 8090
rect 8116 8026 8168 8032
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8128 7410 8156 7890
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7378 4992 7434 5001
rect 7378 4927 7434 4936
rect 7392 4690 7420 4927
rect 7760 4826 7788 6190
rect 7944 5846 7972 7278
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8128 6798 8156 7142
rect 8220 6866 8248 8502
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8312 7274 8340 8434
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8404 7546 8432 7754
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8496 7478 8524 8230
rect 8484 7472 8536 7478
rect 8484 7414 8536 7420
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 8392 6928 8444 6934
rect 8392 6870 8444 6876
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8220 6322 8248 6802
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 8220 5778 8248 6258
rect 8312 5846 8340 6734
rect 8404 5914 8432 6870
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8300 5840 8352 5846
rect 8300 5782 8352 5788
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8300 5704 8352 5710
rect 8404 5692 8432 5850
rect 8496 5846 8524 7414
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 8352 5664 8432 5692
rect 8300 5646 8352 5652
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7472 4616 7524 4622
rect 8036 4604 8064 5034
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 8116 4616 8168 4622
rect 8036 4576 8116 4604
rect 7472 4558 7524 4564
rect 8116 4558 8168 4564
rect 7012 4150 7064 4156
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 7116 4134 7328 4162
rect 6550 4040 6606 4049
rect 6550 3975 6606 3984
rect 6564 3534 6592 3975
rect 7116 3942 7144 4134
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6184 3460 6236 3466
rect 6184 3402 6236 3408
rect 6196 3058 6224 3402
rect 6288 3126 6316 3470
rect 7116 3369 7144 3878
rect 7208 3641 7236 4014
rect 7484 4010 7512 4558
rect 8128 4282 8156 4558
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 7472 4004 7524 4010
rect 7472 3946 7524 3952
rect 7194 3632 7250 3641
rect 7194 3567 7250 3576
rect 7102 3360 7158 3369
rect 6630 3292 6938 3301
rect 7102 3295 7158 3304
rect 6630 3290 6636 3292
rect 6692 3290 6716 3292
rect 6772 3290 6796 3292
rect 6852 3290 6876 3292
rect 6932 3290 6938 3292
rect 6692 3238 6694 3290
rect 6874 3238 6876 3290
rect 6630 3236 6636 3238
rect 6692 3236 6716 3238
rect 6772 3236 6796 3238
rect 6852 3236 6876 3238
rect 6932 3236 6938 3238
rect 6630 3227 6938 3236
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6276 3120 6328 3126
rect 6276 3062 6328 3068
rect 6564 3058 6592 3130
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6552 2916 6604 2922
rect 6552 2858 6604 2864
rect 5920 2746 6040 2774
rect 5920 2446 5948 2746
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 6000 2372 6052 2378
rect 6000 2314 6052 2320
rect 5816 1012 5868 1018
rect 5816 954 5868 960
rect 4712 886 4764 892
rect 4724 800 4752 886
rect 5368 870 5580 898
rect 5368 800 5396 870
rect 6012 800 6040 2314
rect 6564 1442 6592 2858
rect 7116 2446 7144 3295
rect 7484 2990 7512 3946
rect 7852 3534 7880 4082
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7944 3058 7972 4014
rect 8128 3534 8156 4218
rect 8220 3670 8248 4694
rect 8312 4146 8340 5170
rect 8588 5166 8616 12038
rect 8680 10674 8708 14214
rect 8864 13326 8892 16934
rect 9140 16658 9168 17614
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 9140 16250 9168 16594
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9140 15570 9168 16186
rect 9128 15564 9180 15570
rect 9128 15506 9180 15512
rect 9140 15026 9168 15506
rect 9128 15020 9180 15026
rect 9128 14962 9180 14968
rect 9232 14618 9260 19654
rect 9471 19068 9779 19077
rect 9471 19066 9477 19068
rect 9533 19066 9557 19068
rect 9613 19066 9637 19068
rect 9693 19066 9717 19068
rect 9773 19066 9779 19068
rect 9533 19014 9535 19066
rect 9715 19014 9717 19066
rect 9471 19012 9477 19014
rect 9533 19012 9557 19014
rect 9613 19012 9637 19014
rect 9693 19012 9717 19014
rect 9773 19012 9779 19014
rect 9471 19003 9779 19012
rect 9471 17980 9779 17989
rect 9471 17978 9477 17980
rect 9533 17978 9557 17980
rect 9613 17978 9637 17980
rect 9693 17978 9717 17980
rect 9773 17978 9779 17980
rect 9533 17926 9535 17978
rect 9715 17926 9717 17978
rect 9471 17924 9477 17926
rect 9533 17924 9557 17926
rect 9613 17924 9637 17926
rect 9693 17924 9717 17926
rect 9773 17924 9779 17926
rect 9471 17915 9779 17924
rect 9471 16892 9779 16901
rect 9471 16890 9477 16892
rect 9533 16890 9557 16892
rect 9613 16890 9637 16892
rect 9693 16890 9717 16892
rect 9773 16890 9779 16892
rect 9533 16838 9535 16890
rect 9715 16838 9717 16890
rect 9471 16836 9477 16838
rect 9533 16836 9557 16838
rect 9613 16836 9637 16838
rect 9693 16836 9717 16838
rect 9773 16836 9779 16838
rect 9471 16827 9779 16836
rect 9471 15804 9779 15813
rect 9471 15802 9477 15804
rect 9533 15802 9557 15804
rect 9613 15802 9637 15804
rect 9693 15802 9717 15804
rect 9773 15802 9779 15804
rect 9533 15750 9535 15802
rect 9715 15750 9717 15802
rect 9471 15748 9477 15750
rect 9533 15748 9557 15750
rect 9613 15748 9637 15750
rect 9693 15748 9717 15750
rect 9773 15748 9779 15750
rect 9471 15739 9779 15748
rect 9471 14716 9779 14725
rect 9471 14714 9477 14716
rect 9533 14714 9557 14716
rect 9613 14714 9637 14716
rect 9693 14714 9717 14716
rect 9773 14714 9779 14716
rect 9533 14662 9535 14714
rect 9715 14662 9717 14714
rect 9471 14660 9477 14662
rect 9533 14660 9557 14662
rect 9613 14660 9637 14662
rect 9693 14660 9717 14662
rect 9773 14660 9779 14662
rect 9471 14651 9779 14660
rect 9220 14612 9272 14618
rect 9220 14554 9272 14560
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9232 13530 9260 14214
rect 9471 13628 9779 13637
rect 9471 13626 9477 13628
rect 9533 13626 9557 13628
rect 9613 13626 9637 13628
rect 9693 13626 9717 13628
rect 9773 13626 9779 13628
rect 9533 13574 9535 13626
rect 9715 13574 9717 13626
rect 9471 13572 9477 13574
rect 9533 13572 9557 13574
rect 9613 13572 9637 13574
rect 9693 13572 9717 13574
rect 9773 13572 9779 13574
rect 9471 13563 9779 13572
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 8864 12918 8892 13262
rect 8852 12912 8904 12918
rect 8852 12854 8904 12860
rect 9036 12844 9088 12850
rect 9220 12844 9272 12850
rect 9088 12804 9168 12832
rect 9036 12786 9088 12792
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8772 10810 8800 11698
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8864 9450 8892 11698
rect 8944 11688 8996 11694
rect 8944 11630 8996 11636
rect 8956 11218 8984 11630
rect 9140 11558 9168 12804
rect 9220 12786 9272 12792
rect 9232 12374 9260 12786
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9220 12368 9272 12374
rect 9220 12310 9272 12316
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 9048 10554 9076 11086
rect 9140 10674 9168 11494
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9048 10526 9168 10554
rect 9140 10062 9168 10526
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 8956 9926 8984 9998
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 8956 9450 8984 9862
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8944 9444 8996 9450
rect 8944 9386 8996 9392
rect 9140 8974 9168 9998
rect 9232 9178 9260 12038
rect 9324 11132 9352 12582
rect 9471 12540 9779 12549
rect 9471 12538 9477 12540
rect 9533 12538 9557 12540
rect 9613 12538 9637 12540
rect 9693 12538 9717 12540
rect 9773 12538 9779 12540
rect 9533 12486 9535 12538
rect 9715 12486 9717 12538
rect 9471 12484 9477 12486
rect 9533 12484 9557 12486
rect 9613 12484 9637 12486
rect 9693 12484 9717 12486
rect 9773 12484 9779 12486
rect 9471 12475 9779 12484
rect 9876 12238 9904 21286
rect 9968 12850 9996 21490
rect 11992 21418 12020 21966
rect 11980 21412 12032 21418
rect 11980 21354 12032 21360
rect 10966 20904 11022 20913
rect 10966 20839 10968 20848
rect 11020 20839 11022 20848
rect 10968 20810 11020 20816
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 11072 20602 11100 20742
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11428 20460 11480 20466
rect 11428 20402 11480 20408
rect 11244 20324 11296 20330
rect 11244 20266 11296 20272
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 10152 14414 10180 15302
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9600 11558 9628 12174
rect 10060 11762 10088 13126
rect 10244 12850 10272 16934
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10336 12374 10364 19654
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10612 15638 10640 17138
rect 10600 15632 10652 15638
rect 10600 15574 10652 15580
rect 10416 15360 10468 15366
rect 10416 15302 10468 15308
rect 10324 12368 10376 12374
rect 10324 12310 10376 12316
rect 10232 12164 10284 12170
rect 10232 12106 10284 12112
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9471 11452 9779 11461
rect 9471 11450 9477 11452
rect 9533 11450 9557 11452
rect 9613 11450 9637 11452
rect 9693 11450 9717 11452
rect 9773 11450 9779 11452
rect 9533 11398 9535 11450
rect 9715 11398 9717 11450
rect 9471 11396 9477 11398
rect 9533 11396 9557 11398
rect 9613 11396 9637 11398
rect 9693 11396 9717 11398
rect 9773 11396 9779 11398
rect 9471 11387 9779 11396
rect 9404 11144 9456 11150
rect 9324 11104 9404 11132
rect 9404 11086 9456 11092
rect 9312 10804 9364 10810
rect 9312 10746 9364 10752
rect 9324 9586 9352 10746
rect 9416 10418 9444 11086
rect 10152 11082 10180 11698
rect 10244 11694 10272 12106
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 9407 10390 9444 10418
rect 9407 10282 9435 10390
rect 9471 10364 9779 10373
rect 9471 10362 9477 10364
rect 9533 10362 9557 10364
rect 9613 10362 9637 10364
rect 9693 10362 9717 10364
rect 9773 10362 9779 10364
rect 9533 10310 9535 10362
rect 9715 10310 9717 10362
rect 9471 10308 9477 10310
rect 9533 10308 9557 10310
rect 9613 10308 9637 10310
rect 9693 10308 9717 10310
rect 9773 10308 9779 10310
rect 9471 10299 9779 10308
rect 9407 10254 9444 10282
rect 9416 9722 9444 10254
rect 9876 10130 9904 11018
rect 10152 10742 10180 11018
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 9770 9616 9826 9625
rect 9312 9580 9364 9586
rect 9770 9551 9826 9560
rect 9864 9580 9916 9586
rect 9312 9522 9364 9528
rect 9784 9518 9812 9551
rect 9864 9522 9916 9528
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8864 7410 8892 8230
rect 9140 8022 9168 8910
rect 9128 8016 9180 8022
rect 9128 7958 9180 7964
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8956 7342 8984 7686
rect 9140 7546 9168 7822
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8852 7268 8904 7274
rect 8852 7210 8904 7216
rect 8864 5234 8892 7210
rect 8956 6322 8984 7278
rect 9048 7002 9076 7346
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8852 5228 8904 5234
rect 8852 5170 8904 5176
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8116 3528 8168 3534
rect 8036 3476 8116 3482
rect 8036 3470 8168 3476
rect 8036 3454 8156 3470
rect 8312 3466 8340 4082
rect 8496 4010 8524 4626
rect 8772 4146 8800 4966
rect 9140 4826 9168 7346
rect 9324 6202 9352 9386
rect 9471 9276 9779 9285
rect 9471 9274 9477 9276
rect 9533 9274 9557 9276
rect 9613 9274 9637 9276
rect 9693 9274 9717 9276
rect 9773 9274 9779 9276
rect 9533 9222 9535 9274
rect 9715 9222 9717 9274
rect 9471 9220 9477 9222
rect 9533 9220 9557 9222
rect 9613 9220 9637 9222
rect 9693 9220 9717 9222
rect 9773 9220 9779 9222
rect 9471 9211 9779 9220
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9600 8294 9628 8842
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9471 8188 9779 8197
rect 9471 8186 9477 8188
rect 9533 8186 9557 8188
rect 9613 8186 9637 8188
rect 9693 8186 9717 8188
rect 9773 8186 9779 8188
rect 9533 8134 9535 8186
rect 9715 8134 9717 8186
rect 9471 8132 9477 8134
rect 9533 8132 9557 8134
rect 9613 8132 9637 8134
rect 9693 8132 9717 8134
rect 9773 8132 9779 8134
rect 9471 8123 9779 8132
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9784 7188 9812 8026
rect 9876 7546 9904 9522
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9784 7160 9904 7188
rect 9471 7100 9779 7109
rect 9471 7098 9477 7100
rect 9533 7098 9557 7100
rect 9613 7098 9637 7100
rect 9693 7098 9717 7100
rect 9773 7098 9779 7100
rect 9533 7046 9535 7098
rect 9715 7046 9717 7098
rect 9471 7044 9477 7046
rect 9533 7044 9557 7046
rect 9613 7044 9637 7046
rect 9693 7044 9717 7046
rect 9773 7044 9779 7046
rect 9471 7035 9779 7044
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 6458 9720 6598
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9232 6174 9444 6202
rect 9232 5914 9260 6174
rect 9416 6118 9444 6174
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9220 5296 9272 5302
rect 9220 5238 9272 5244
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8300 3460 8352 3466
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 8036 2514 8064 3454
rect 8300 3402 8352 3408
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 8128 3194 8156 3334
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8128 2990 8156 3130
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 8404 2922 8432 3878
rect 8496 3058 8524 3946
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 8588 2854 8616 3674
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 8128 2514 8156 2790
rect 8864 2650 8892 3878
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8956 3058 8984 3334
rect 9048 3058 9076 4422
rect 9232 4146 9260 5238
rect 9324 4690 9352 6054
rect 9471 6012 9779 6021
rect 9471 6010 9477 6012
rect 9533 6010 9557 6012
rect 9613 6010 9637 6012
rect 9693 6010 9717 6012
rect 9773 6010 9779 6012
rect 9533 5958 9535 6010
rect 9715 5958 9717 6010
rect 9471 5956 9477 5958
rect 9533 5956 9557 5958
rect 9613 5956 9637 5958
rect 9693 5956 9717 5958
rect 9773 5956 9779 5958
rect 9471 5947 9779 5956
rect 9588 5840 9640 5846
rect 9588 5782 9640 5788
rect 9600 5166 9628 5782
rect 9876 5234 9904 7160
rect 9968 6866 9996 10610
rect 10152 10266 10180 10678
rect 10244 10554 10272 11630
rect 10428 11218 10456 15302
rect 10704 13326 10732 19450
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10520 12986 10548 13126
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10704 12918 10732 13262
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10520 11830 10548 12038
rect 10508 11824 10560 11830
rect 10508 11766 10560 11772
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10336 10674 10364 11154
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 10600 10600 10652 10606
rect 10244 10526 10364 10554
rect 10600 10542 10652 10548
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 10060 8974 10088 10066
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 10152 8634 10180 10202
rect 10336 9518 10364 10526
rect 10612 10470 10640 10542
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10232 9376 10284 9382
rect 10230 9344 10232 9353
rect 10284 9344 10286 9353
rect 10230 9279 10286 9288
rect 10336 9042 10364 9454
rect 10520 9450 10548 10406
rect 10508 9444 10560 9450
rect 10508 9386 10560 9392
rect 10612 9042 10640 10406
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10612 8838 10640 8978
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 10060 8022 10088 8298
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 10060 6866 10088 7958
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10244 7546 10272 7890
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10336 7546 10364 7822
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10428 7410 10456 8366
rect 10612 8090 10640 8366
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10336 6866 10364 7142
rect 10428 7002 10456 7346
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10060 6458 10088 6802
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9471 4924 9779 4933
rect 9471 4922 9477 4924
rect 9533 4922 9557 4924
rect 9613 4922 9637 4924
rect 9693 4922 9717 4924
rect 9773 4922 9779 4924
rect 9533 4870 9535 4922
rect 9715 4870 9717 4922
rect 9471 4868 9477 4870
rect 9533 4868 9557 4870
rect 9613 4868 9637 4870
rect 9693 4868 9717 4870
rect 9773 4868 9779 4870
rect 9471 4859 9779 4868
rect 10152 4690 10180 6734
rect 10336 6662 10364 6802
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10612 5710 10640 6598
rect 10704 6089 10732 12718
rect 10796 8378 10824 14486
rect 10888 14346 10916 14758
rect 10876 14340 10928 14346
rect 10876 14282 10928 14288
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10888 10198 10916 10406
rect 10876 10192 10928 10198
rect 10876 10134 10928 10140
rect 10980 9586 11008 18566
rect 11072 15434 11100 20198
rect 11256 15910 11284 20266
rect 11440 20058 11468 20402
rect 12084 20058 12112 22034
rect 12544 22030 12572 22086
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12311 21788 12619 21797
rect 12311 21786 12317 21788
rect 12373 21786 12397 21788
rect 12453 21786 12477 21788
rect 12533 21786 12557 21788
rect 12613 21786 12619 21788
rect 12373 21734 12375 21786
rect 12555 21734 12557 21786
rect 12311 21732 12317 21734
rect 12373 21732 12397 21734
rect 12453 21732 12477 21734
rect 12533 21732 12557 21734
rect 12613 21732 12619 21734
rect 12311 21723 12619 21732
rect 12728 21554 12756 22102
rect 15660 22092 15712 22098
rect 15660 22034 15712 22040
rect 13174 21992 13230 22001
rect 13174 21927 13176 21936
rect 13228 21927 13230 21936
rect 13176 21898 13228 21904
rect 13084 21888 13136 21894
rect 13084 21830 13136 21836
rect 14740 21888 14792 21894
rect 14740 21830 14792 21836
rect 13096 21554 13124 21830
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12532 21548 12584 21554
rect 12532 21490 12584 21496
rect 12716 21548 12768 21554
rect 12716 21490 12768 21496
rect 13084 21548 13136 21554
rect 13084 21490 13136 21496
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 11428 20052 11480 20058
rect 11428 19994 11480 20000
rect 12072 20052 12124 20058
rect 12072 19994 12124 20000
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11336 19848 11388 19854
rect 11336 19790 11388 19796
rect 11348 19378 11376 19790
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11716 17882 11744 19314
rect 11704 17876 11756 17882
rect 11704 17818 11756 17824
rect 11612 17672 11664 17678
rect 11612 17614 11664 17620
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11348 16726 11376 17274
rect 11336 16720 11388 16726
rect 11336 16662 11388 16668
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 11072 13258 11100 14962
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 11164 13870 11192 14282
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 11256 13410 11284 15846
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11164 13382 11284 13410
rect 11164 13258 11192 13382
rect 11348 13326 11376 15438
rect 11440 15366 11468 16390
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11440 13682 11468 15302
rect 11532 13802 11560 17478
rect 11624 14618 11652 17614
rect 11900 17270 11928 17614
rect 11888 17264 11940 17270
rect 11888 17206 11940 17212
rect 11704 16516 11756 16522
rect 11704 16458 11756 16464
rect 11716 16182 11744 16458
rect 11704 16176 11756 16182
rect 11704 16118 11756 16124
rect 11716 15502 11744 16118
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11716 13938 11744 14350
rect 11808 14074 11836 14350
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11900 13938 11928 14418
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11520 13796 11572 13802
rect 11520 13738 11572 13744
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11440 13654 11560 13682
rect 11336 13320 11388 13326
rect 11242 13288 11298 13297
rect 11060 13252 11112 13258
rect 11060 13194 11112 13200
rect 11152 13252 11204 13258
rect 11336 13262 11388 13268
rect 11242 13223 11298 13232
rect 11152 13194 11204 13200
rect 11072 9654 11100 13194
rect 11164 12646 11192 13194
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11256 11558 11284 13223
rect 11348 13190 11376 13262
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11256 9722 11284 10950
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10876 9376 10928 9382
rect 10874 9344 10876 9353
rect 10928 9344 10930 9353
rect 10874 9279 10930 9288
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 10796 8350 10916 8378
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10796 7886 10824 8230
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10888 6798 10916 8350
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 10980 6798 11008 7414
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10690 6080 10746 6089
rect 10690 6015 10746 6024
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10520 5234 10548 5646
rect 10704 5234 10732 6015
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10876 5228 10928 5234
rect 10980 5216 11008 6734
rect 11072 6254 11100 8230
rect 11164 7478 11192 8434
rect 11348 7818 11376 8774
rect 11440 8498 11468 11834
rect 11532 11268 11560 13654
rect 11716 13410 11744 13738
rect 11624 13382 11744 13410
rect 11624 12306 11652 13382
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11716 12918 11744 13262
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 11900 12714 11928 13874
rect 11992 13297 12020 19858
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 12084 18426 12112 18634
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 12084 15706 12112 18158
rect 12176 16454 12204 21490
rect 12452 21010 12480 21490
rect 12544 21457 12572 21490
rect 12530 21448 12586 21457
rect 12530 21383 12586 21392
rect 12440 21004 12492 21010
rect 12440 20946 12492 20952
rect 12716 20936 12768 20942
rect 12716 20878 12768 20884
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 12311 20700 12619 20709
rect 12311 20698 12317 20700
rect 12373 20698 12397 20700
rect 12453 20698 12477 20700
rect 12533 20698 12557 20700
rect 12613 20698 12619 20700
rect 12373 20646 12375 20698
rect 12555 20646 12557 20698
rect 12311 20644 12317 20646
rect 12373 20644 12397 20646
rect 12453 20644 12477 20646
rect 12533 20644 12557 20646
rect 12613 20644 12619 20646
rect 12311 20635 12619 20644
rect 12311 19612 12619 19621
rect 12311 19610 12317 19612
rect 12373 19610 12397 19612
rect 12453 19610 12477 19612
rect 12533 19610 12557 19612
rect 12613 19610 12619 19612
rect 12373 19558 12375 19610
rect 12555 19558 12557 19610
rect 12311 19556 12317 19558
rect 12373 19556 12397 19558
rect 12453 19556 12477 19558
rect 12533 19556 12557 19558
rect 12613 19556 12619 19558
rect 12311 19547 12619 19556
rect 12440 19440 12492 19446
rect 12440 19382 12492 19388
rect 12452 19310 12480 19382
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12544 18630 12572 19246
rect 12636 18834 12664 19314
rect 12728 18902 12756 20878
rect 12912 19514 12940 20878
rect 13096 20534 13124 21490
rect 13820 21480 13872 21486
rect 13820 21422 13872 21428
rect 14096 21480 14148 21486
rect 14096 21422 14148 21428
rect 13268 21344 13320 21350
rect 13268 21286 13320 21292
rect 13280 20942 13308 21286
rect 13268 20936 13320 20942
rect 13268 20878 13320 20884
rect 13832 20618 13860 21422
rect 13636 20596 13688 20602
rect 13636 20538 13688 20544
rect 13740 20590 13860 20618
rect 13084 20528 13136 20534
rect 13084 20470 13136 20476
rect 13096 20398 13124 20470
rect 13084 20392 13136 20398
rect 13084 20334 13136 20340
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 12716 18896 12768 18902
rect 12716 18838 12768 18844
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12311 18524 12619 18533
rect 12311 18522 12317 18524
rect 12373 18522 12397 18524
rect 12453 18522 12477 18524
rect 12533 18522 12557 18524
rect 12613 18522 12619 18524
rect 12373 18470 12375 18522
rect 12555 18470 12557 18522
rect 12311 18468 12317 18470
rect 12373 18468 12397 18470
rect 12453 18468 12477 18470
rect 12533 18468 12557 18470
rect 12613 18468 12619 18470
rect 12311 18459 12619 18468
rect 12728 18290 12756 18838
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12311 17436 12619 17445
rect 12311 17434 12317 17436
rect 12373 17434 12397 17436
rect 12453 17434 12477 17436
rect 12533 17434 12557 17436
rect 12613 17434 12619 17436
rect 12373 17382 12375 17434
rect 12555 17382 12557 17434
rect 12311 17380 12317 17382
rect 12373 17380 12397 17382
rect 12453 17380 12477 17382
rect 12533 17380 12557 17382
rect 12613 17380 12619 17382
rect 12311 17371 12619 17380
rect 12728 17338 12756 17614
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 12820 17134 12848 18702
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12544 16658 12572 16934
rect 12912 16658 12940 19314
rect 12992 19236 13044 19242
rect 12992 19178 13044 19184
rect 13004 18834 13032 19178
rect 12992 18828 13044 18834
rect 12992 18770 13044 18776
rect 13084 18760 13136 18766
rect 13084 18702 13136 18708
rect 12992 18352 13044 18358
rect 12992 18294 13044 18300
rect 13004 17066 13032 18294
rect 13096 17338 13124 18702
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 13188 17882 13216 18566
rect 13280 18358 13308 18566
rect 13268 18352 13320 18358
rect 13268 18294 13320 18300
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 13268 17876 13320 17882
rect 13268 17818 13320 17824
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 13176 17196 13228 17202
rect 13096 17156 13176 17184
rect 12992 17060 13044 17066
rect 12992 17002 13044 17008
rect 13096 16946 13124 17156
rect 13280 17184 13308 17818
rect 13360 17672 13412 17678
rect 13358 17640 13360 17649
rect 13412 17640 13414 17649
rect 13358 17575 13414 17584
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13372 17202 13400 17274
rect 13228 17156 13308 17184
rect 13360 17196 13412 17202
rect 13176 17138 13228 17144
rect 13360 17138 13412 17144
rect 13176 17060 13228 17066
rect 13176 17002 13228 17008
rect 13004 16918 13124 16946
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12900 16652 12952 16658
rect 12900 16594 12952 16600
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 12311 16348 12619 16357
rect 12311 16346 12317 16348
rect 12373 16346 12397 16348
rect 12453 16346 12477 16348
rect 12533 16346 12557 16348
rect 12613 16346 12619 16348
rect 12373 16294 12375 16346
rect 12555 16294 12557 16346
rect 12311 16292 12317 16294
rect 12373 16292 12397 16294
rect 12453 16292 12477 16294
rect 12533 16292 12557 16294
rect 12613 16292 12619 16294
rect 12311 16283 12619 16292
rect 12164 16108 12216 16114
rect 12164 16050 12216 16056
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 12176 15570 12204 16050
rect 12624 15972 12676 15978
rect 12624 15914 12676 15920
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 12164 15564 12216 15570
rect 12360 15552 12388 15846
rect 12440 15564 12492 15570
rect 12360 15524 12440 15552
rect 12164 15506 12216 15512
rect 12440 15506 12492 15512
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 12084 13870 12112 14894
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 11978 13288 12034 13297
rect 11978 13223 12034 13232
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11992 12850 12020 13126
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11612 11280 11664 11286
rect 11532 11240 11612 11268
rect 11612 11222 11664 11228
rect 11624 11082 11652 11222
rect 11716 11150 11744 11494
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11612 11076 11664 11082
rect 11612 11018 11664 11024
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11716 10062 11744 10746
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11808 9994 11836 11018
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11428 8492 11480 8498
rect 11428 8434 11480 8440
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 11152 7472 11204 7478
rect 11204 7432 11284 7460
rect 11152 7414 11204 7420
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 11072 5710 11100 6190
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 10928 5188 11008 5216
rect 10876 5170 10928 5176
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 9140 3194 9168 4014
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8956 2774 8984 2994
rect 8956 2746 9168 2774
rect 9140 2650 9168 2746
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 8116 2508 8168 2514
rect 8116 2450 8168 2456
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 6630 2204 6938 2213
rect 6630 2202 6636 2204
rect 6692 2202 6716 2204
rect 6772 2202 6796 2204
rect 6852 2202 6876 2204
rect 6932 2202 6938 2204
rect 6692 2150 6694 2202
rect 6874 2150 6876 2202
rect 6630 2148 6636 2150
rect 6692 2148 6716 2150
rect 6772 2148 6796 2150
rect 6852 2148 6876 2150
rect 6932 2148 6938 2150
rect 6630 2139 6938 2148
rect 6564 1414 6684 1442
rect 6656 800 6684 1414
rect 7288 1080 7340 1086
rect 7288 1022 7340 1028
rect 7300 800 7328 1022
rect 7932 1012 7984 1018
rect 7932 954 7984 960
rect 7944 800 7972 954
rect 8576 944 8628 950
rect 8576 886 8628 892
rect 8588 800 8616 886
rect 9232 800 9260 3470
rect 9324 2854 9352 4626
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9471 3836 9779 3845
rect 9471 3834 9477 3836
rect 9533 3834 9557 3836
rect 9613 3834 9637 3836
rect 9693 3834 9717 3836
rect 9773 3834 9779 3836
rect 9533 3782 9535 3834
rect 9715 3782 9717 3834
rect 9471 3780 9477 3782
rect 9533 3780 9557 3782
rect 9613 3780 9637 3782
rect 9693 3780 9717 3782
rect 9773 3780 9779 3782
rect 9471 3771 9779 3780
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 9471 2748 9779 2757
rect 9471 2746 9477 2748
rect 9533 2746 9557 2748
rect 9613 2746 9637 2748
rect 9693 2746 9717 2748
rect 9773 2746 9779 2748
rect 9533 2694 9535 2746
rect 9715 2694 9717 2746
rect 9471 2692 9477 2694
rect 9533 2692 9557 2694
rect 9613 2692 9637 2694
rect 9693 2692 9717 2694
rect 9773 2692 9779 2694
rect 9471 2683 9779 2692
rect 9876 2530 9904 3878
rect 9968 3670 9996 4490
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9956 3528 10008 3534
rect 10060 3482 10088 4422
rect 10244 3534 10272 4558
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10008 3476 10088 3482
rect 9956 3470 10088 3476
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 9968 3454 10088 3470
rect 9968 3097 9996 3454
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10152 3126 10180 3334
rect 10140 3120 10192 3126
rect 9954 3088 10010 3097
rect 10140 3062 10192 3068
rect 9954 3023 10010 3032
rect 9784 2502 9904 2530
rect 9784 950 9812 2502
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 9772 944 9824 950
rect 9772 886 9824 892
rect 9876 800 9904 2382
rect 10336 1018 10364 3878
rect 10428 1086 10456 3878
rect 10508 3596 10560 3602
rect 10508 3538 10560 3544
rect 10520 3126 10548 3538
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 10416 1080 10468 1086
rect 10416 1022 10468 1028
rect 10324 1012 10376 1018
rect 10324 954 10376 960
rect 10520 800 10548 2790
rect 10704 2514 10732 5170
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10796 3738 10824 4422
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10796 2854 10824 3674
rect 11072 3534 11100 4422
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11072 2990 11100 3470
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 2990 11192 3402
rect 11256 3398 11284 7432
rect 11348 5846 11376 7754
rect 11440 7342 11468 7822
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 11336 5840 11388 5846
rect 11336 5782 11388 5788
rect 11440 5710 11468 7278
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 11348 5370 11376 5646
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11440 5273 11468 5646
rect 11426 5264 11482 5273
rect 11426 5199 11482 5208
rect 11532 4826 11560 9658
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 11624 6662 11652 8298
rect 11716 8090 11744 8910
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11808 7970 11836 8434
rect 11716 7942 11836 7970
rect 11716 6934 11744 7942
rect 11704 6928 11756 6934
rect 11704 6870 11756 6876
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11336 4548 11388 4554
rect 11336 4490 11388 4496
rect 11348 3398 11376 4490
rect 11624 4078 11652 6598
rect 11716 5642 11744 6870
rect 11900 5846 11928 12106
rect 11992 11778 12020 12786
rect 12084 12238 12112 13806
rect 12176 13326 12204 15506
rect 12636 15434 12664 15914
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12311 15260 12619 15269
rect 12311 15258 12317 15260
rect 12373 15258 12397 15260
rect 12453 15258 12477 15260
rect 12533 15258 12557 15260
rect 12613 15258 12619 15260
rect 12373 15206 12375 15258
rect 12555 15206 12557 15258
rect 12311 15204 12317 15206
rect 12373 15204 12397 15206
rect 12453 15204 12477 15206
rect 12533 15204 12557 15206
rect 12613 15204 12619 15206
rect 12311 15195 12619 15204
rect 12728 14958 12756 15302
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12311 14172 12619 14181
rect 12311 14170 12317 14172
rect 12373 14170 12397 14172
rect 12453 14170 12477 14172
rect 12533 14170 12557 14172
rect 12613 14170 12619 14172
rect 12373 14118 12375 14170
rect 12555 14118 12557 14170
rect 12311 14116 12317 14118
rect 12373 14116 12397 14118
rect 12453 14116 12477 14118
rect 12533 14116 12557 14118
rect 12613 14116 12619 14118
rect 12311 14107 12619 14116
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12544 13326 12572 14010
rect 12820 13530 12848 16594
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12912 13394 12940 14962
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12084 11898 12112 12174
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 12176 11830 12204 13262
rect 12311 13084 12619 13093
rect 12311 13082 12317 13084
rect 12373 13082 12397 13084
rect 12453 13082 12477 13084
rect 12533 13082 12557 13084
rect 12613 13082 12619 13084
rect 12373 13030 12375 13082
rect 12555 13030 12557 13082
rect 12311 13028 12317 13030
rect 12373 13028 12397 13030
rect 12453 13028 12477 13030
rect 12533 13028 12557 13030
rect 12613 13028 12619 13030
rect 12311 13019 12619 13028
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 12728 12238 12756 12854
rect 13004 12306 13032 16918
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 13096 14006 13124 16730
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 12311 11996 12619 12005
rect 12311 11994 12317 11996
rect 12373 11994 12397 11996
rect 12453 11994 12477 11996
rect 12533 11994 12557 11996
rect 12613 11994 12619 11996
rect 12373 11942 12375 11994
rect 12555 11942 12557 11994
rect 12311 11940 12317 11942
rect 12373 11940 12397 11942
rect 12453 11940 12477 11942
rect 12533 11940 12557 11942
rect 12613 11940 12619 11942
rect 12311 11931 12619 11940
rect 12164 11824 12216 11830
rect 11992 11762 12112 11778
rect 12164 11766 12216 11772
rect 12716 11824 12768 11830
rect 12716 11766 12768 11772
rect 11992 11756 12124 11762
rect 11992 11750 12072 11756
rect 12072 11698 12124 11704
rect 12084 11234 12112 11698
rect 11992 11206 12112 11234
rect 11992 10062 12020 11206
rect 12311 10908 12619 10917
rect 12311 10906 12317 10908
rect 12373 10906 12397 10908
rect 12453 10906 12477 10908
rect 12533 10906 12557 10908
rect 12613 10906 12619 10908
rect 12373 10854 12375 10906
rect 12555 10854 12557 10906
rect 12311 10852 12317 10854
rect 12373 10852 12397 10854
rect 12453 10852 12477 10854
rect 12533 10852 12557 10854
rect 12613 10852 12619 10854
rect 12311 10843 12619 10852
rect 12728 10810 12756 11766
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11992 5914 12020 8910
rect 12084 8090 12112 10610
rect 12268 9908 12296 10610
rect 12176 9880 12296 9908
rect 12176 9625 12204 9880
rect 12311 9820 12619 9829
rect 12311 9818 12317 9820
rect 12373 9818 12397 9820
rect 12453 9818 12477 9820
rect 12533 9818 12557 9820
rect 12613 9818 12619 9820
rect 12373 9766 12375 9818
rect 12555 9766 12557 9818
rect 12311 9764 12317 9766
rect 12373 9764 12397 9766
rect 12453 9764 12477 9766
rect 12533 9764 12557 9766
rect 12613 9764 12619 9766
rect 12311 9755 12619 9764
rect 12728 9654 12756 10746
rect 12716 9648 12768 9654
rect 12162 9616 12218 9625
rect 12716 9590 12768 9596
rect 12162 9551 12218 9560
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 12176 8566 12204 8978
rect 12544 8974 12572 9318
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12311 8732 12619 8741
rect 12311 8730 12317 8732
rect 12373 8730 12397 8732
rect 12453 8730 12477 8732
rect 12533 8730 12557 8732
rect 12613 8730 12619 8732
rect 12373 8678 12375 8730
rect 12555 8678 12557 8730
rect 12311 8676 12317 8678
rect 12373 8676 12397 8678
rect 12453 8676 12477 8678
rect 12533 8676 12557 8678
rect 12613 8676 12619 8678
rect 12311 8667 12619 8676
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12544 8498 12572 8570
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12820 7886 12848 8842
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12084 6798 12112 7346
rect 12176 6866 12204 7822
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12311 7644 12619 7653
rect 12311 7642 12317 7644
rect 12373 7642 12397 7644
rect 12453 7642 12477 7644
rect 12533 7642 12557 7644
rect 12613 7642 12619 7644
rect 12373 7590 12375 7642
rect 12555 7590 12557 7642
rect 12311 7588 12317 7590
rect 12373 7588 12397 7590
rect 12453 7588 12477 7590
rect 12533 7588 12557 7590
rect 12613 7588 12619 7590
rect 12311 7579 12619 7588
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 11888 5840 11940 5846
rect 11888 5782 11940 5788
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 11808 5574 11836 5782
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11808 5234 11836 5510
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 11426 3496 11482 3505
rect 11426 3431 11428 3440
rect 11480 3431 11482 3440
rect 11428 3402 11480 3408
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 11336 3392 11388 3398
rect 11336 3334 11388 3340
rect 11348 3058 11376 3334
rect 11336 3052 11388 3058
rect 11336 2994 11388 3000
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 10692 2508 10744 2514
rect 10692 2450 10744 2456
rect 11440 2446 11468 3402
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 11532 3194 11560 3334
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11624 3058 11652 4014
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11716 3369 11744 3878
rect 11702 3360 11758 3369
rect 11702 3295 11758 3304
rect 11808 3233 11836 3878
rect 11888 3664 11940 3670
rect 11888 3606 11940 3612
rect 11794 3224 11850 3233
rect 11900 3194 11928 3606
rect 11794 3159 11850 3168
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 10980 898 11008 2382
rect 10980 870 11192 898
rect 11164 800 11192 870
rect 11808 800 11836 2450
rect 11992 2446 12020 5170
rect 12084 4826 12112 6326
rect 12176 5914 12204 6802
rect 12268 6662 12296 7414
rect 12728 7206 12756 7754
rect 13004 7750 13032 12106
rect 13096 11354 13124 13942
rect 13188 13530 13216 17002
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 13280 14618 13308 16594
rect 13464 15706 13492 19790
rect 13542 19272 13598 19281
rect 13542 19207 13544 19216
rect 13596 19207 13598 19216
rect 13544 19178 13596 19184
rect 13544 18284 13596 18290
rect 13544 18226 13596 18232
rect 13556 17746 13584 18226
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13544 17060 13596 17066
rect 13544 17002 13596 17008
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13280 14074 13308 14554
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13176 13320 13228 13326
rect 13176 13262 13228 13268
rect 13188 12986 13216 13262
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13280 12646 13308 14010
rect 13372 13433 13400 15438
rect 13358 13424 13414 13433
rect 13358 13359 13414 13368
rect 13464 12714 13492 15642
rect 13556 15094 13584 17002
rect 13648 16046 13676 20538
rect 13740 20466 13768 20590
rect 14108 20534 14136 21422
rect 14200 21321 14228 21490
rect 14660 21418 14688 21490
rect 14648 21412 14700 21418
rect 14648 21354 14700 21360
rect 14186 21312 14242 21321
rect 14186 21247 14242 21256
rect 14200 21146 14228 21247
rect 14188 21140 14240 21146
rect 14188 21082 14240 21088
rect 14280 21072 14332 21078
rect 14280 21014 14332 21020
rect 14292 20806 14320 21014
rect 14752 20942 14780 21830
rect 15016 21616 15068 21622
rect 15016 21558 15068 21564
rect 14832 21412 14884 21418
rect 14832 21354 14884 21360
rect 14556 20936 14608 20942
rect 14556 20878 14608 20884
rect 14740 20936 14792 20942
rect 14740 20878 14792 20884
rect 14372 20868 14424 20874
rect 14372 20810 14424 20816
rect 14280 20800 14332 20806
rect 14280 20742 14332 20748
rect 14096 20528 14148 20534
rect 14096 20470 14148 20476
rect 14292 20466 14320 20742
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 13820 20460 13872 20466
rect 13820 20402 13872 20408
rect 14280 20460 14332 20466
rect 14280 20402 14332 20408
rect 13740 19446 13768 20402
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 13832 18970 13860 20402
rect 14292 20058 14320 20402
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14384 19854 14412 20810
rect 14568 19990 14596 20878
rect 14556 19984 14608 19990
rect 14556 19926 14608 19932
rect 14372 19848 14424 19854
rect 14372 19790 14424 19796
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 13912 19712 13964 19718
rect 13912 19654 13964 19660
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13924 18714 13952 19654
rect 14004 19236 14056 19242
rect 14004 19178 14056 19184
rect 13832 18686 13952 18714
rect 13832 17678 13860 18686
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13924 18426 13952 18566
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13728 17604 13780 17610
rect 13728 17546 13780 17552
rect 13636 16040 13688 16046
rect 13636 15982 13688 15988
rect 13648 15502 13676 15982
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 13544 15088 13596 15094
rect 13544 15030 13596 15036
rect 13556 13258 13584 15030
rect 13648 14482 13676 15438
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13544 13252 13596 13258
rect 13544 13194 13596 13200
rect 13452 12708 13504 12714
rect 13452 12650 13504 12656
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13280 11898 13308 12174
rect 13544 12164 13596 12170
rect 13544 12106 13596 12112
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 13280 11082 13308 11834
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 13280 10742 13308 11018
rect 13268 10736 13320 10742
rect 13268 10678 13320 10684
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 13188 10130 13216 10474
rect 13280 10198 13308 10542
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 13188 8956 13216 10066
rect 13280 9926 13308 10134
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 13280 9722 13308 9862
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13372 9518 13400 11630
rect 13556 11354 13584 12106
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13648 10266 13676 13466
rect 13740 12918 13768 17546
rect 13832 17338 13860 17614
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 13820 17196 13872 17202
rect 13924 17184 13952 18362
rect 14016 18086 14044 19178
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 14096 18216 14148 18222
rect 14096 18158 14148 18164
rect 14004 18080 14056 18086
rect 14004 18022 14056 18028
rect 14004 17196 14056 17202
rect 13924 17156 14004 17184
rect 13820 17138 13872 17144
rect 14004 17138 14056 17144
rect 13832 14278 13860 17138
rect 14016 16522 14044 17138
rect 14004 16516 14056 16522
rect 14004 16458 14056 16464
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13924 14346 13952 15846
rect 14108 15144 14136 18158
rect 14188 18148 14240 18154
rect 14188 18090 14240 18096
rect 14200 17746 14228 18090
rect 14188 17740 14240 17746
rect 14188 17682 14240 17688
rect 14292 17678 14320 18226
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14384 17202 14412 19790
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 14476 18766 14504 19654
rect 14568 19378 14596 19790
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14740 19304 14792 19310
rect 14740 19246 14792 19252
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14568 18970 14596 19110
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14752 18873 14780 19246
rect 14844 19174 14872 21354
rect 15028 21146 15056 21558
rect 15152 21244 15460 21253
rect 15152 21242 15158 21244
rect 15214 21242 15238 21244
rect 15294 21242 15318 21244
rect 15374 21242 15398 21244
rect 15454 21242 15460 21244
rect 15214 21190 15216 21242
rect 15396 21190 15398 21242
rect 15152 21188 15158 21190
rect 15214 21188 15238 21190
rect 15294 21188 15318 21190
rect 15374 21188 15398 21190
rect 15454 21188 15460 21190
rect 15152 21179 15460 21188
rect 15016 21140 15068 21146
rect 15016 21082 15068 21088
rect 15672 20942 15700 22034
rect 17420 21962 17448 24200
rect 20833 22332 21141 22341
rect 20833 22330 20839 22332
rect 20895 22330 20919 22332
rect 20975 22330 20999 22332
rect 21055 22330 21079 22332
rect 21135 22330 21141 22332
rect 20895 22278 20897 22330
rect 21077 22278 21079 22330
rect 20833 22276 20839 22278
rect 20895 22276 20919 22278
rect 20975 22276 20999 22278
rect 21055 22276 21079 22278
rect 21135 22276 21141 22278
rect 20833 22267 21141 22276
rect 20444 22024 20496 22030
rect 20442 21992 20444 22001
rect 20720 22024 20772 22030
rect 20496 21992 20498 22001
rect 17408 21956 17460 21962
rect 20720 21966 20772 21972
rect 20442 21927 20498 21936
rect 17408 21898 17460 21904
rect 15844 21888 15896 21894
rect 15844 21830 15896 21836
rect 18880 21888 18932 21894
rect 18880 21830 18932 21836
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 15856 21554 15884 21830
rect 17992 21788 18300 21797
rect 17992 21786 17998 21788
rect 18054 21786 18078 21788
rect 18134 21786 18158 21788
rect 18214 21786 18238 21788
rect 18294 21786 18300 21788
rect 18054 21734 18056 21786
rect 18236 21734 18238 21786
rect 17992 21732 17998 21734
rect 18054 21732 18078 21734
rect 18134 21732 18158 21734
rect 18214 21732 18238 21734
rect 18294 21732 18300 21734
rect 17992 21723 18300 21732
rect 15936 21616 15988 21622
rect 15936 21558 15988 21564
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15752 21344 15804 21350
rect 15752 21286 15804 21292
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 14924 20800 14976 20806
rect 14924 20742 14976 20748
rect 14936 20466 14964 20742
rect 15672 20534 15700 20878
rect 15200 20528 15252 20534
rect 15200 20470 15252 20476
rect 15660 20528 15712 20534
rect 15660 20470 15712 20476
rect 14924 20460 14976 20466
rect 14924 20402 14976 20408
rect 14924 20256 14976 20262
rect 15212 20244 15240 20470
rect 15764 20466 15792 21286
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15568 20392 15620 20398
rect 15568 20334 15620 20340
rect 15212 20216 15516 20244
rect 14924 20198 14976 20204
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14738 18864 14794 18873
rect 14738 18799 14794 18808
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14648 18692 14700 18698
rect 14648 18634 14700 18640
rect 14568 17814 14596 18634
rect 14556 17808 14608 17814
rect 14556 17750 14608 17756
rect 14660 17746 14688 18634
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14372 17196 14424 17202
rect 14016 15116 14136 15144
rect 14200 17156 14372 17184
rect 13912 14340 13964 14346
rect 13912 14282 13964 14288
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13924 13870 13952 14282
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13728 12912 13780 12918
rect 13728 12854 13780 12860
rect 13832 12850 13860 13330
rect 14016 13326 14044 15116
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14108 14414 14136 14962
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14108 13938 14136 14350
rect 14200 14074 14228 17156
rect 14372 17138 14424 17144
rect 14464 17128 14516 17134
rect 14462 17096 14464 17105
rect 14516 17096 14518 17105
rect 14462 17031 14518 17040
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 14372 16720 14424 16726
rect 14372 16662 14424 16668
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14292 15026 14320 15438
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 14280 14544 14332 14550
rect 14280 14486 14332 14492
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 13912 12980 13964 12986
rect 14016 12968 14044 13262
rect 13964 12940 14044 12968
rect 13912 12922 13964 12928
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13740 10810 13768 12174
rect 13832 11762 13860 12310
rect 14108 11830 14136 13874
rect 14292 13870 14320 14486
rect 14280 13864 14332 13870
rect 14280 13806 14332 13812
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14200 12850 14228 13466
rect 14384 12986 14412 16662
rect 14568 15094 14596 16934
rect 14556 15088 14608 15094
rect 14556 15030 14608 15036
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 14648 15020 14700 15026
rect 14648 14962 14700 14968
rect 14476 13841 14504 14962
rect 14556 14884 14608 14890
rect 14556 14826 14608 14832
rect 14568 14278 14596 14826
rect 14660 14618 14688 14962
rect 14752 14906 14780 18022
rect 14844 16561 14872 18226
rect 14936 17542 14964 20198
rect 15152 20156 15460 20165
rect 15152 20154 15158 20156
rect 15214 20154 15238 20156
rect 15294 20154 15318 20156
rect 15374 20154 15398 20156
rect 15454 20154 15460 20156
rect 15214 20102 15216 20154
rect 15396 20102 15398 20154
rect 15152 20100 15158 20102
rect 15214 20100 15238 20102
rect 15294 20100 15318 20102
rect 15374 20100 15398 20102
rect 15454 20100 15460 20102
rect 15152 20091 15460 20100
rect 15016 20052 15068 20058
rect 15016 19994 15068 20000
rect 15028 18306 15056 19994
rect 15108 19916 15160 19922
rect 15108 19858 15160 19864
rect 15120 19446 15148 19858
rect 15108 19440 15160 19446
rect 15108 19382 15160 19388
rect 15152 19068 15460 19077
rect 15152 19066 15158 19068
rect 15214 19066 15238 19068
rect 15294 19066 15318 19068
rect 15374 19066 15398 19068
rect 15454 19066 15460 19068
rect 15214 19014 15216 19066
rect 15396 19014 15398 19066
rect 15152 19012 15158 19014
rect 15214 19012 15238 19014
rect 15294 19012 15318 19014
rect 15374 19012 15398 19014
rect 15454 19012 15460 19014
rect 15152 19003 15460 19012
rect 15108 18692 15160 18698
rect 15108 18634 15160 18640
rect 15120 18426 15148 18634
rect 15488 18426 15516 20216
rect 15580 20058 15608 20334
rect 15752 20324 15804 20330
rect 15752 20266 15804 20272
rect 15568 20052 15620 20058
rect 15568 19994 15620 20000
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15108 18420 15160 18426
rect 15108 18362 15160 18368
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15028 18278 15148 18306
rect 15120 18222 15148 18278
rect 15476 18284 15528 18290
rect 15580 18272 15608 19110
rect 15528 18244 15608 18272
rect 15476 18226 15528 18232
rect 15016 18216 15068 18222
rect 15014 18184 15016 18193
rect 15108 18216 15160 18222
rect 15068 18184 15070 18193
rect 15108 18158 15160 18164
rect 15014 18119 15070 18128
rect 15120 18086 15148 18158
rect 15488 18086 15516 18226
rect 15108 18080 15160 18086
rect 15108 18022 15160 18028
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15152 17980 15460 17989
rect 15152 17978 15158 17980
rect 15214 17978 15238 17980
rect 15294 17978 15318 17980
rect 15374 17978 15398 17980
rect 15454 17978 15460 17980
rect 15214 17926 15216 17978
rect 15396 17926 15398 17978
rect 15152 17924 15158 17926
rect 15214 17924 15238 17926
rect 15294 17924 15318 17926
rect 15374 17924 15398 17926
rect 15454 17924 15460 17926
rect 15152 17915 15460 17924
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 15106 17640 15162 17649
rect 14924 17536 14976 17542
rect 14924 17478 14976 17484
rect 14924 17332 14976 17338
rect 14924 17274 14976 17280
rect 14830 16552 14886 16561
rect 14936 16522 14964 17274
rect 15028 16998 15056 17614
rect 15106 17575 15162 17584
rect 15120 17066 15148 17575
rect 15212 17202 15240 17682
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15108 17060 15160 17066
rect 15108 17002 15160 17008
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 15152 16892 15460 16901
rect 15152 16890 15158 16892
rect 15214 16890 15238 16892
rect 15294 16890 15318 16892
rect 15374 16890 15398 16892
rect 15454 16890 15460 16892
rect 15214 16838 15216 16890
rect 15396 16838 15398 16890
rect 15152 16836 15158 16838
rect 15214 16836 15238 16838
rect 15294 16836 15318 16838
rect 15374 16836 15398 16838
rect 15454 16836 15460 16838
rect 15152 16827 15460 16836
rect 14830 16487 14886 16496
rect 14924 16516 14976 16522
rect 14924 16458 14976 16464
rect 15384 16448 15436 16454
rect 15488 16436 15516 18022
rect 15672 17678 15700 19858
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15568 17604 15620 17610
rect 15568 17546 15620 17552
rect 15436 16408 15516 16436
rect 15384 16390 15436 16396
rect 15016 16040 15068 16046
rect 15014 16008 15016 16017
rect 15068 16008 15070 16017
rect 15396 15994 15424 16390
rect 15580 16114 15608 17546
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 15672 16114 15700 17478
rect 15764 16250 15792 20266
rect 15856 19281 15884 21490
rect 15842 19272 15898 19281
rect 15842 19207 15898 19216
rect 15856 16522 15884 19207
rect 15948 19174 15976 21558
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 17868 21548 17920 21554
rect 17868 21490 17920 21496
rect 18144 21548 18196 21554
rect 18144 21490 18196 21496
rect 17132 21412 17184 21418
rect 17132 21354 17184 21360
rect 16028 21344 16080 21350
rect 16028 21286 16080 21292
rect 16040 19242 16068 21286
rect 17144 21146 17172 21354
rect 17132 21140 17184 21146
rect 17132 21082 17184 21088
rect 17420 21078 17448 21490
rect 17880 21078 17908 21490
rect 18156 21146 18184 21490
rect 18892 21486 18920 21830
rect 19260 21690 19288 21830
rect 19248 21684 19300 21690
rect 19248 21626 19300 21632
rect 19432 21616 19484 21622
rect 19432 21558 19484 21564
rect 18880 21480 18932 21486
rect 18880 21422 18932 21428
rect 18144 21140 18196 21146
rect 18144 21082 18196 21088
rect 17408 21072 17460 21078
rect 17408 21014 17460 21020
rect 17868 21072 17920 21078
rect 17868 21014 17920 21020
rect 16304 21004 16356 21010
rect 16304 20946 16356 20952
rect 16212 20936 16264 20942
rect 16212 20878 16264 20884
rect 16120 20324 16172 20330
rect 16120 20266 16172 20272
rect 16132 19922 16160 20266
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 16224 19514 16252 20878
rect 16316 19786 16344 20946
rect 18156 20942 18184 21082
rect 18248 20998 18460 21026
rect 18892 21010 18920 21422
rect 19340 21072 19392 21078
rect 19340 21014 19392 21020
rect 17408 20936 17460 20942
rect 17408 20878 17460 20884
rect 17500 20936 17552 20942
rect 17500 20878 17552 20884
rect 18144 20936 18196 20942
rect 18144 20878 18196 20884
rect 16396 20528 16448 20534
rect 16396 20470 16448 20476
rect 16304 19780 16356 19786
rect 16304 19722 16356 19728
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 16028 19236 16080 19242
rect 16028 19178 16080 19184
rect 15936 19168 15988 19174
rect 15936 19110 15988 19116
rect 16040 18902 16068 19178
rect 16028 18896 16080 18902
rect 16028 18838 16080 18844
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 15936 17808 15988 17814
rect 15936 17750 15988 17756
rect 15844 16516 15896 16522
rect 15844 16458 15896 16464
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15396 15966 15792 15994
rect 15014 15943 15070 15952
rect 15028 15570 15056 15943
rect 15152 15804 15460 15813
rect 15152 15802 15158 15804
rect 15214 15802 15238 15804
rect 15294 15802 15318 15804
rect 15374 15802 15398 15804
rect 15454 15802 15460 15804
rect 15214 15750 15216 15802
rect 15396 15750 15398 15802
rect 15152 15748 15158 15750
rect 15214 15748 15238 15750
rect 15294 15748 15318 15750
rect 15374 15748 15398 15750
rect 15454 15748 15460 15750
rect 15152 15739 15460 15748
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 14924 15360 14976 15366
rect 14924 15302 14976 15308
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 14936 15162 14964 15302
rect 14924 15156 14976 15162
rect 14924 15098 14976 15104
rect 15212 14958 15240 15302
rect 15200 14952 15252 14958
rect 14752 14878 14872 14906
rect 15200 14894 15252 14900
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14752 14414 14780 14758
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 14462 13832 14518 13841
rect 14462 13767 14518 13776
rect 14464 13252 14516 13258
rect 14464 13194 14516 13200
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14476 12889 14504 13194
rect 14462 12880 14518 12889
rect 14188 12844 14240 12850
rect 14462 12815 14518 12824
rect 14188 12786 14240 12792
rect 14200 11830 14228 12786
rect 14476 12782 14504 12815
rect 14464 12776 14516 12782
rect 14384 12736 14464 12764
rect 14384 12238 14412 12736
rect 14464 12718 14516 12724
rect 14568 12306 14596 14214
rect 14844 14090 14872 14878
rect 15152 14716 15460 14725
rect 15152 14714 15158 14716
rect 15214 14714 15238 14716
rect 15294 14714 15318 14716
rect 15374 14714 15398 14716
rect 15454 14714 15460 14716
rect 15214 14662 15216 14714
rect 15396 14662 15398 14714
rect 15152 14660 15158 14662
rect 15214 14660 15238 14662
rect 15294 14660 15318 14662
rect 15374 14660 15398 14662
rect 15454 14660 15460 14662
rect 15152 14651 15460 14660
rect 15488 14618 15516 15438
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15108 14340 15160 14346
rect 15108 14282 15160 14288
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 14660 14062 14872 14090
rect 14660 13530 14688 14062
rect 14832 14000 14884 14006
rect 14832 13942 14884 13948
rect 14844 13530 14872 13942
rect 15120 13938 15148 14282
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 14936 13530 14964 13874
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 14648 13524 14700 13530
rect 14648 13466 14700 13472
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 14924 13524 14976 13530
rect 14924 13466 14976 13472
rect 14740 13456 14792 13462
rect 14740 13398 14792 13404
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14660 12442 14688 13126
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 13912 11824 13964 11830
rect 13912 11766 13964 11772
rect 14096 11824 14148 11830
rect 14096 11766 14148 11772
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13832 11082 13860 11698
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13740 9654 13768 10746
rect 13832 9654 13860 11018
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13372 9042 13400 9454
rect 13832 9058 13860 9590
rect 13924 9586 13952 11766
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 14016 10674 14044 11630
rect 14292 11626 14320 12038
rect 14476 11762 14504 12174
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14280 11620 14332 11626
rect 14280 11562 14332 11568
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13740 9030 13860 9058
rect 14004 9104 14056 9110
rect 14004 9046 14056 9052
rect 13268 8968 13320 8974
rect 13188 8928 13268 8956
rect 13268 8910 13320 8916
rect 13280 8498 13308 8910
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13084 7812 13136 7818
rect 13084 7754 13136 7760
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 12716 7200 12768 7206
rect 12716 7142 12768 7148
rect 13004 6934 13032 7686
rect 13096 7002 13124 7754
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 12992 6928 13044 6934
rect 12992 6870 13044 6876
rect 13188 6746 13216 8434
rect 13740 8090 13768 9030
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13832 8362 13860 8910
rect 14016 8498 14044 9046
rect 14108 8498 14136 11154
rect 14292 10674 14320 11562
rect 14568 11354 14596 11834
rect 14752 11354 14780 13398
rect 14936 13258 14964 13466
rect 14924 13252 14976 13258
rect 14924 13194 14976 13200
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14844 12850 14872 13126
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14924 12300 14976 12306
rect 14924 12242 14976 12248
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14936 11082 14964 12242
rect 15028 11762 15056 13806
rect 15152 13628 15460 13637
rect 15152 13626 15158 13628
rect 15214 13626 15238 13628
rect 15294 13626 15318 13628
rect 15374 13626 15398 13628
rect 15454 13626 15460 13628
rect 15214 13574 15216 13626
rect 15396 13574 15398 13626
rect 15152 13572 15158 13574
rect 15214 13572 15238 13574
rect 15294 13572 15318 13574
rect 15374 13572 15398 13574
rect 15454 13572 15460 13574
rect 15152 13563 15460 13572
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15304 12850 15332 13262
rect 15396 12918 15424 13466
rect 15488 12918 15516 13806
rect 15580 13326 15608 14282
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15384 12912 15436 12918
rect 15384 12854 15436 12860
rect 15476 12912 15528 12918
rect 15672 12866 15700 14962
rect 15764 13190 15792 15966
rect 15844 15428 15896 15434
rect 15844 15370 15896 15376
rect 15856 15162 15884 15370
rect 15844 15156 15896 15162
rect 15844 15098 15896 15104
rect 15948 15026 15976 17750
rect 16040 17746 16068 18226
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 16040 17542 16068 17682
rect 16224 17678 16252 19246
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 16132 17202 16160 17478
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 15936 14884 15988 14890
rect 15936 14826 15988 14832
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15476 12854 15528 12860
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15580 12838 15700 12866
rect 15752 12844 15804 12850
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15152 12540 15460 12549
rect 15152 12538 15158 12540
rect 15214 12538 15238 12540
rect 15294 12538 15318 12540
rect 15374 12538 15398 12540
rect 15454 12538 15460 12540
rect 15214 12486 15216 12538
rect 15396 12486 15398 12538
rect 15152 12484 15158 12486
rect 15214 12484 15238 12486
rect 15294 12484 15318 12486
rect 15374 12484 15398 12486
rect 15454 12484 15460 12486
rect 15152 12475 15460 12484
rect 15200 12368 15252 12374
rect 15200 12310 15252 12316
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 15212 11642 15240 12310
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15396 11801 15424 11834
rect 15382 11792 15438 11801
rect 15382 11727 15438 11736
rect 15028 11614 15240 11642
rect 15028 11268 15056 11614
rect 15152 11452 15460 11461
rect 15152 11450 15158 11452
rect 15214 11450 15238 11452
rect 15294 11450 15318 11452
rect 15374 11450 15398 11452
rect 15454 11450 15460 11452
rect 15214 11398 15216 11450
rect 15396 11398 15398 11450
rect 15152 11396 15158 11398
rect 15214 11396 15238 11398
rect 15294 11396 15318 11398
rect 15374 11396 15398 11398
rect 15454 11396 15460 11398
rect 15152 11387 15460 11396
rect 15028 11240 15240 11268
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 15212 10674 15240 11240
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15304 10810 15332 11086
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 14188 10532 14240 10538
rect 14188 10474 14240 10480
rect 14200 9722 14228 10474
rect 14292 10198 14320 10610
rect 15212 10577 15240 10610
rect 15198 10568 15254 10577
rect 15198 10503 15254 10512
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14280 10192 14332 10198
rect 14280 10134 14332 10140
rect 14384 10062 14412 10406
rect 15152 10364 15460 10373
rect 15152 10362 15158 10364
rect 15214 10362 15238 10364
rect 15294 10362 15318 10364
rect 15374 10362 15398 10364
rect 15454 10362 15460 10364
rect 15214 10310 15216 10362
rect 15396 10310 15398 10362
rect 15152 10308 15158 10310
rect 15214 10308 15238 10310
rect 15294 10308 15318 10310
rect 15374 10308 15398 10310
rect 15454 10308 15460 10310
rect 15152 10299 15460 10308
rect 15488 10062 15516 12582
rect 15580 12374 15608 12838
rect 15752 12786 15804 12792
rect 15568 12368 15620 12374
rect 15568 12310 15620 12316
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15580 10810 15608 12174
rect 15672 11286 15700 12174
rect 15660 11280 15712 11286
rect 15660 11222 15712 11228
rect 15764 11218 15792 12786
rect 15856 12374 15884 14554
rect 15948 14278 15976 14826
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 15844 12368 15896 12374
rect 15844 12310 15896 12316
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15856 11762 15884 12174
rect 15948 11898 15976 14214
rect 16040 13530 16068 14962
rect 16132 14618 16160 17138
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 16224 13938 16252 17614
rect 16316 17338 16344 19722
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 16408 16114 16436 20470
rect 17420 19854 17448 20878
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17512 19514 17540 20878
rect 18248 20806 18276 20998
rect 18328 20868 18380 20874
rect 18328 20810 18380 20816
rect 18236 20800 18288 20806
rect 18236 20742 18288 20748
rect 17992 20700 18300 20709
rect 17992 20698 17998 20700
rect 18054 20698 18078 20700
rect 18134 20698 18158 20700
rect 18214 20698 18238 20700
rect 18294 20698 18300 20700
rect 18054 20646 18056 20698
rect 18236 20646 18238 20698
rect 17992 20644 17998 20646
rect 18054 20644 18078 20646
rect 18134 20644 18158 20646
rect 18214 20644 18238 20646
rect 18294 20644 18300 20646
rect 17992 20635 18300 20644
rect 18340 20602 18368 20810
rect 18328 20596 18380 20602
rect 18328 20538 18380 20544
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 17992 19612 18300 19621
rect 17992 19610 17998 19612
rect 18054 19610 18078 19612
rect 18134 19610 18158 19612
rect 18214 19610 18238 19612
rect 18294 19610 18300 19612
rect 18054 19558 18056 19610
rect 18236 19558 18238 19610
rect 17992 19556 17998 19558
rect 18054 19556 18078 19558
rect 18134 19556 18158 19558
rect 18214 19556 18238 19558
rect 18294 19556 18300 19558
rect 17992 19547 18300 19556
rect 17500 19508 17552 19514
rect 17500 19450 17552 19456
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 17408 19304 17460 19310
rect 17408 19246 17460 19252
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16776 18426 16804 18702
rect 16764 18420 16816 18426
rect 16764 18362 16816 18368
rect 16580 17672 16632 17678
rect 16486 17640 16542 17649
rect 16580 17614 16632 17620
rect 16486 17575 16542 17584
rect 16500 16590 16528 17575
rect 16592 16946 16620 17614
rect 16672 17604 16724 17610
rect 16672 17546 16724 17552
rect 16684 17338 16712 17546
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16592 16918 16712 16946
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16408 15570 16436 16050
rect 16396 15564 16448 15570
rect 16448 15524 16528 15552
rect 16396 15506 16448 15512
rect 16304 15020 16356 15026
rect 16304 14962 16356 14968
rect 16316 14482 16344 14962
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 16040 12170 16068 12854
rect 16224 12764 16252 13126
rect 16316 12918 16344 14418
rect 16500 14074 16528 15524
rect 16684 15366 16712 16918
rect 16776 16658 16804 18362
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16868 17270 16896 17614
rect 16856 17264 16908 17270
rect 17144 17252 17172 19246
rect 17236 18834 17264 19246
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 17236 17610 17264 18770
rect 17316 18692 17368 18698
rect 17316 18634 17368 18640
rect 17328 17814 17356 18634
rect 17420 18358 17448 19246
rect 17972 18680 18000 19314
rect 18236 18760 18288 18766
rect 18340 18748 18368 19790
rect 18432 18766 18460 20998
rect 18880 21004 18932 21010
rect 18880 20946 18932 20952
rect 18788 19712 18840 19718
rect 18788 19654 18840 19660
rect 18800 19514 18828 19654
rect 18512 19508 18564 19514
rect 18512 19450 18564 19456
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 18524 19310 18552 19450
rect 18604 19440 18656 19446
rect 18604 19382 18656 19388
rect 18512 19304 18564 19310
rect 18512 19246 18564 19252
rect 18512 18828 18564 18834
rect 18512 18770 18564 18776
rect 18288 18720 18368 18748
rect 18236 18702 18288 18708
rect 17880 18652 18000 18680
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 17500 18420 17552 18426
rect 17500 18362 17552 18368
rect 17408 18352 17460 18358
rect 17408 18294 17460 18300
rect 17408 18080 17460 18086
rect 17408 18022 17460 18028
rect 17316 17808 17368 17814
rect 17316 17750 17368 17756
rect 17224 17604 17276 17610
rect 17224 17546 17276 17552
rect 17316 17264 17368 17270
rect 17144 17224 17316 17252
rect 16856 17206 16908 17212
rect 17316 17206 17368 17212
rect 17328 16658 17356 17206
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 16856 16584 16908 16590
rect 16776 16532 16856 16538
rect 16776 16526 16908 16532
rect 16776 16510 16896 16526
rect 16948 16516 17000 16522
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16670 15192 16726 15201
rect 16670 15127 16726 15136
rect 16684 15026 16712 15127
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16408 13326 16436 14010
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 16224 12736 16344 12764
rect 16316 12220 16344 12736
rect 16500 12238 16528 14010
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16592 13161 16620 13262
rect 16578 13152 16634 13161
rect 16578 13087 16634 13096
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16592 12306 16620 12582
rect 16684 12374 16712 13262
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 16224 12192 16344 12220
rect 16488 12232 16540 12238
rect 16028 12164 16080 12170
rect 16028 12106 16080 12112
rect 15936 11892 15988 11898
rect 15936 11834 15988 11840
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15844 10668 15896 10674
rect 15948 10656 15976 11834
rect 16224 11558 16252 12192
rect 16488 12174 16540 12180
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 15896 10628 15976 10656
rect 15844 10610 15896 10616
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 14200 8498 14228 9658
rect 14292 8974 14320 9998
rect 14832 9988 14884 9994
rect 14832 9930 14884 9936
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14464 9444 14516 9450
rect 14464 9386 14516 9392
rect 14372 9036 14424 9042
rect 14372 8978 14424 8984
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14384 8566 14412 8978
rect 14476 8974 14504 9386
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14372 8560 14424 8566
rect 14372 8502 14424 8508
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13188 6718 13308 6746
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 12311 6556 12619 6565
rect 12311 6554 12317 6556
rect 12373 6554 12397 6556
rect 12453 6554 12477 6556
rect 12533 6554 12557 6556
rect 12613 6554 12619 6556
rect 12373 6502 12375 6554
rect 12555 6502 12557 6554
rect 12311 6500 12317 6502
rect 12373 6500 12397 6502
rect 12453 6500 12477 6502
rect 12533 6500 12557 6502
rect 12613 6500 12619 6502
rect 12311 6491 12619 6500
rect 13188 6390 13216 6598
rect 13176 6384 13228 6390
rect 13176 6326 13228 6332
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12164 5908 12216 5914
rect 12164 5850 12216 5856
rect 12268 5778 12296 6190
rect 12256 5772 12308 5778
rect 12256 5714 12308 5720
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12311 5468 12619 5477
rect 12311 5466 12317 5468
rect 12373 5466 12397 5468
rect 12453 5466 12477 5468
rect 12533 5466 12557 5468
rect 12613 5466 12619 5468
rect 12373 5414 12375 5466
rect 12555 5414 12557 5466
rect 12311 5412 12317 5414
rect 12373 5412 12397 5414
rect 12453 5412 12477 5414
rect 12533 5412 12557 5414
rect 12613 5412 12619 5414
rect 12311 5403 12619 5412
rect 12728 5370 12756 5510
rect 13280 5370 13308 6718
rect 13372 5710 13400 7142
rect 13728 6928 13780 6934
rect 13728 6870 13780 6876
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13464 6322 13492 6734
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 13268 5364 13320 5370
rect 13268 5306 13320 5312
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 12254 5128 12310 5137
rect 12254 5063 12310 5072
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 12176 4486 12204 4762
rect 12268 4622 12296 5063
rect 12728 4826 12756 5170
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12311 4380 12619 4389
rect 12311 4378 12317 4380
rect 12373 4378 12397 4380
rect 12453 4378 12477 4380
rect 12533 4378 12557 4380
rect 12613 4378 12619 4380
rect 12373 4326 12375 4378
rect 12555 4326 12557 4378
rect 12311 4324 12317 4326
rect 12373 4324 12397 4326
rect 12453 4324 12477 4326
rect 12533 4324 12557 4326
rect 12613 4324 12619 4326
rect 12311 4315 12619 4324
rect 12164 4004 12216 4010
rect 12164 3946 12216 3952
rect 12176 2990 12204 3946
rect 12728 3602 12756 4558
rect 12820 3738 12848 5170
rect 12912 5098 12940 5170
rect 12900 5092 12952 5098
rect 12900 5034 12952 5040
rect 12912 4758 12940 5034
rect 13372 5030 13400 5646
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 12900 4752 12952 4758
rect 12900 4694 12952 4700
rect 13556 4282 13584 6054
rect 13648 5778 13676 6054
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13648 4758 13676 4966
rect 13636 4752 13688 4758
rect 13636 4694 13688 4700
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12311 3292 12619 3301
rect 12311 3290 12317 3292
rect 12373 3290 12397 3292
rect 12453 3290 12477 3292
rect 12533 3290 12557 3292
rect 12613 3290 12619 3292
rect 12373 3238 12375 3290
rect 12555 3238 12557 3290
rect 12311 3236 12317 3238
rect 12373 3236 12397 3238
rect 12453 3236 12477 3238
rect 12533 3236 12557 3238
rect 12613 3236 12619 3238
rect 12311 3227 12619 3236
rect 12728 3194 12756 3538
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 12164 2984 12216 2990
rect 12164 2926 12216 2932
rect 12912 2650 12940 3470
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13280 3058 13308 3334
rect 13464 3058 13492 4218
rect 13556 4185 13584 4218
rect 13542 4176 13598 4185
rect 13542 4111 13598 4120
rect 13740 4010 13768 6870
rect 13924 6866 13952 8434
rect 14108 7410 14136 8434
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 14292 6798 14320 7346
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14108 6254 14136 6734
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14004 6112 14056 6118
rect 14002 6080 14004 6089
rect 14056 6080 14058 6089
rect 14002 6015 14058 6024
rect 14016 5234 14044 6015
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 13924 4826 13952 4966
rect 13912 4820 13964 4826
rect 13912 4762 13964 4768
rect 14476 4468 14504 8570
rect 14568 8430 14596 8978
rect 14752 8974 14780 9522
rect 14844 9382 14872 9930
rect 14924 9648 14976 9654
rect 14924 9590 14976 9596
rect 14832 9376 14884 9382
rect 14832 9318 14884 9324
rect 14844 9042 14872 9318
rect 14832 9036 14884 9042
rect 14832 8978 14884 8984
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14752 8090 14780 8910
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 14660 7478 14688 7822
rect 14648 7472 14700 7478
rect 14648 7414 14700 7420
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 14568 4622 14596 6190
rect 14752 5710 14780 6190
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14556 4480 14608 4486
rect 14476 4440 14556 4468
rect 14556 4422 14608 4428
rect 14568 4146 14596 4422
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 13726 3088 13782 3097
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 13452 3052 13504 3058
rect 14292 3058 14320 3470
rect 13726 3023 13728 3032
rect 13452 2994 13504 3000
rect 13780 3023 13782 3032
rect 14280 3052 14332 3058
rect 13728 2994 13780 3000
rect 14280 2994 14332 3000
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 12311 2204 12619 2213
rect 12311 2202 12317 2204
rect 12373 2202 12397 2204
rect 12453 2202 12477 2204
rect 12533 2202 12557 2204
rect 12613 2202 12619 2204
rect 12373 2150 12375 2202
rect 12555 2150 12557 2202
rect 12311 2148 12317 2150
rect 12373 2148 12397 2150
rect 12453 2148 12477 2150
rect 12533 2148 12557 2150
rect 12613 2148 12619 2150
rect 12311 2139 12619 2148
rect 12452 870 12572 898
rect 12452 800 12480 870
rect 1490 0 1546 800
rect 2134 0 2190 800
rect 2778 0 2834 800
rect 3422 0 3478 800
rect 4066 0 4122 800
rect 4710 0 4766 800
rect 5354 0 5410 800
rect 5998 0 6054 800
rect 6642 0 6698 800
rect 7286 0 7342 800
rect 7930 0 7986 800
rect 8574 0 8630 800
rect 9218 0 9274 800
rect 9862 0 9918 800
rect 10506 0 10562 800
rect 11150 0 11206 800
rect 11794 0 11850 800
rect 12438 0 12494 800
rect 12544 762 12572 870
rect 12728 762 12756 2382
rect 13096 800 13124 2382
rect 13832 898 13860 2382
rect 13740 870 13860 898
rect 13740 800 13768 870
rect 14384 800 14412 3538
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14568 2961 14596 2994
rect 14554 2952 14610 2961
rect 14554 2887 14610 2896
rect 14660 2514 14688 5170
rect 14752 4622 14780 5306
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14752 4214 14780 4558
rect 14740 4208 14792 4214
rect 14740 4150 14792 4156
rect 14844 3738 14872 8978
rect 14936 8974 14964 9590
rect 15120 9586 15148 9998
rect 15580 9994 15608 10406
rect 15568 9988 15620 9994
rect 15568 9930 15620 9936
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 16040 9518 16068 11154
rect 16224 11082 16252 11494
rect 16316 11150 16344 11494
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 16212 11076 16264 11082
rect 16212 11018 16264 11024
rect 16224 10198 16252 11018
rect 16212 10192 16264 10198
rect 16212 10134 16264 10140
rect 16212 9988 16264 9994
rect 16212 9930 16264 9936
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 15152 9276 15460 9285
rect 15152 9274 15158 9276
rect 15214 9274 15238 9276
rect 15294 9274 15318 9276
rect 15374 9274 15398 9276
rect 15454 9274 15460 9276
rect 15214 9222 15216 9274
rect 15396 9222 15398 9274
rect 15152 9220 15158 9222
rect 15214 9220 15238 9222
rect 15294 9220 15318 9222
rect 15374 9220 15398 9222
rect 15454 9220 15460 9222
rect 15152 9211 15460 9220
rect 15568 9104 15620 9110
rect 15568 9046 15620 9052
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 15580 8634 15608 9046
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 15660 8832 15712 8838
rect 15660 8774 15712 8780
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15152 8188 15460 8197
rect 15152 8186 15158 8188
rect 15214 8186 15238 8188
rect 15294 8186 15318 8188
rect 15374 8186 15398 8188
rect 15454 8186 15460 8188
rect 15214 8134 15216 8186
rect 15396 8134 15398 8186
rect 15152 8132 15158 8134
rect 15214 8132 15238 8134
rect 15294 8132 15318 8134
rect 15374 8132 15398 8134
rect 15454 8132 15460 8134
rect 15152 8123 15460 8132
rect 15488 8090 15516 8570
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 15580 7886 15608 8570
rect 15672 8498 15700 8774
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15568 7880 15620 7886
rect 15568 7822 15620 7828
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 15028 7546 15056 7686
rect 15212 7546 15240 7822
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 15028 7206 15056 7482
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 15028 6254 15056 7142
rect 15152 7100 15460 7109
rect 15152 7098 15158 7100
rect 15214 7098 15238 7100
rect 15294 7098 15318 7100
rect 15374 7098 15398 7100
rect 15454 7098 15460 7100
rect 15214 7046 15216 7098
rect 15396 7046 15398 7098
rect 15152 7044 15158 7046
rect 15214 7044 15238 7046
rect 15294 7044 15318 7046
rect 15374 7044 15398 7046
rect 15454 7044 15460 7046
rect 15152 7035 15460 7044
rect 15580 6662 15608 7686
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15580 6322 15608 6598
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15016 6248 15068 6254
rect 15016 6190 15068 6196
rect 15568 6180 15620 6186
rect 15568 6122 15620 6128
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15152 6012 15460 6021
rect 15152 6010 15158 6012
rect 15214 6010 15238 6012
rect 15294 6010 15318 6012
rect 15374 6010 15398 6012
rect 15454 6010 15460 6012
rect 15214 5958 15216 6010
rect 15396 5958 15398 6010
rect 15152 5956 15158 5958
rect 15214 5956 15238 5958
rect 15294 5956 15318 5958
rect 15374 5956 15398 5958
rect 15454 5956 15460 5958
rect 15152 5947 15460 5956
rect 15108 5704 15160 5710
rect 15028 5664 15108 5692
rect 14924 5636 14976 5642
rect 14924 5578 14976 5584
rect 14936 5370 14964 5578
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 15028 4826 15056 5664
rect 15108 5646 15160 5652
rect 15488 5370 15516 6054
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15292 5296 15344 5302
rect 15292 5238 15344 5244
rect 15304 5030 15332 5238
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15488 5098 15516 5170
rect 15476 5092 15528 5098
rect 15476 5034 15528 5040
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 15152 4924 15460 4933
rect 15152 4922 15158 4924
rect 15214 4922 15238 4924
rect 15294 4922 15318 4924
rect 15374 4922 15398 4924
rect 15454 4922 15460 4924
rect 15214 4870 15216 4922
rect 15396 4870 15398 4922
rect 15152 4868 15158 4870
rect 15214 4868 15238 4870
rect 15294 4868 15318 4870
rect 15374 4868 15398 4870
rect 15454 4868 15460 4870
rect 15152 4859 15460 4868
rect 15016 4820 15068 4826
rect 15016 4762 15068 4768
rect 15488 4264 15516 5034
rect 15580 4826 15608 6122
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15488 4236 15608 4264
rect 15384 4208 15436 4214
rect 15436 4168 15516 4196
rect 15384 4150 15436 4156
rect 15152 3836 15460 3845
rect 15152 3834 15158 3836
rect 15214 3834 15238 3836
rect 15294 3834 15318 3836
rect 15374 3834 15398 3836
rect 15454 3834 15460 3836
rect 15214 3782 15216 3834
rect 15396 3782 15398 3834
rect 15152 3780 15158 3782
rect 15214 3780 15238 3782
rect 15294 3780 15318 3782
rect 15374 3780 15398 3782
rect 15454 3780 15460 3782
rect 15152 3771 15460 3780
rect 14832 3732 14884 3738
rect 14832 3674 14884 3680
rect 14922 3632 14978 3641
rect 14922 3567 14978 3576
rect 14936 3058 14964 3567
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14648 2508 14700 2514
rect 14648 2450 14700 2456
rect 15028 800 15056 3470
rect 15200 3460 15252 3466
rect 15200 3402 15252 3408
rect 15212 2990 15240 3402
rect 15488 3398 15516 4168
rect 15580 3398 15608 4236
rect 15672 3942 15700 7890
rect 15856 7410 15884 8026
rect 15936 7880 15988 7886
rect 15936 7822 15988 7828
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15568 3392 15620 3398
rect 15568 3334 15620 3340
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 15152 2748 15460 2757
rect 15152 2746 15158 2748
rect 15214 2746 15238 2748
rect 15294 2746 15318 2748
rect 15374 2746 15398 2748
rect 15454 2746 15460 2748
rect 15214 2694 15216 2746
rect 15396 2694 15398 2746
rect 15152 2692 15158 2694
rect 15214 2692 15238 2694
rect 15294 2692 15318 2694
rect 15374 2692 15398 2694
rect 15454 2692 15460 2694
rect 15152 2683 15460 2692
rect 15488 2582 15516 3334
rect 15568 3120 15620 3126
rect 15568 3062 15620 3068
rect 15580 2990 15608 3062
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15476 2576 15528 2582
rect 15476 2518 15528 2524
rect 15580 2446 15608 2926
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15672 800 15700 3470
rect 15764 2650 15792 6190
rect 15856 5642 15884 7346
rect 15948 6186 15976 7822
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 15948 5914 15976 6122
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 16040 5710 16068 8910
rect 16224 8634 16252 9930
rect 16316 9654 16344 11086
rect 16500 11082 16528 11290
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 16592 10742 16620 11766
rect 16684 11354 16712 12174
rect 16776 11694 16804 16510
rect 16948 16458 17000 16464
rect 17040 16516 17092 16522
rect 17040 16458 17092 16464
rect 16856 15428 16908 15434
rect 16856 15370 16908 15376
rect 16868 14890 16896 15370
rect 16856 14884 16908 14890
rect 16856 14826 16908 14832
rect 16868 14414 16896 14826
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16854 13832 16910 13841
rect 16854 13767 16856 13776
rect 16908 13767 16910 13776
rect 16856 13738 16908 13744
rect 16960 13682 16988 16458
rect 17052 16114 17080 16458
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 17224 16108 17276 16114
rect 17224 16050 17276 16056
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 17052 15706 17080 15846
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 17236 15026 17264 16050
rect 17328 15910 17356 16594
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17328 15162 17356 15846
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 16868 13654 16988 13682
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16868 11626 16896 13654
rect 17052 13530 17080 14894
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 17144 13938 17172 14418
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 17144 13410 17172 13874
rect 17144 13394 17356 13410
rect 17420 13394 17448 18022
rect 17512 17626 17540 18362
rect 17604 17746 17632 18566
rect 17880 18408 17908 18652
rect 17992 18524 18300 18533
rect 17992 18522 17998 18524
rect 18054 18522 18078 18524
rect 18134 18522 18158 18524
rect 18214 18522 18238 18524
rect 18294 18522 18300 18524
rect 18054 18470 18056 18522
rect 18236 18470 18238 18522
rect 17992 18468 17998 18470
rect 18054 18468 18078 18470
rect 18134 18468 18158 18470
rect 18214 18468 18238 18470
rect 18294 18468 18300 18470
rect 17992 18459 18300 18468
rect 18340 18426 18368 18720
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18432 18426 18460 18702
rect 18328 18420 18380 18426
rect 17880 18380 18000 18408
rect 17776 18284 17828 18290
rect 17776 18226 17828 18232
rect 17682 18184 17738 18193
rect 17682 18119 17738 18128
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 17512 17598 17632 17626
rect 17500 17128 17552 17134
rect 17500 17070 17552 17076
rect 17512 16590 17540 17070
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17512 15638 17540 16526
rect 17604 16114 17632 17598
rect 17696 17134 17724 18119
rect 17684 17128 17736 17134
rect 17684 17070 17736 17076
rect 17592 16108 17644 16114
rect 17592 16050 17644 16056
rect 17696 15994 17724 17070
rect 17788 16658 17816 18226
rect 17972 18154 18000 18380
rect 18328 18362 18380 18368
rect 18420 18420 18472 18426
rect 18420 18362 18472 18368
rect 17960 18148 18012 18154
rect 17960 18090 18012 18096
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 18328 18080 18380 18086
rect 18328 18022 18380 18028
rect 17776 16652 17828 16658
rect 17776 16594 17828 16600
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 17604 15966 17724 15994
rect 17500 15632 17552 15638
rect 17500 15574 17552 15580
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17132 13388 17356 13394
rect 17184 13382 17356 13388
rect 17132 13330 17184 13336
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17144 12850 17172 12922
rect 17222 12880 17278 12889
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 17132 12844 17184 12850
rect 17222 12815 17224 12824
rect 17132 12786 17184 12792
rect 17276 12815 17278 12824
rect 17224 12786 17276 12792
rect 16960 12442 16988 12786
rect 17040 12708 17092 12714
rect 17040 12650 17092 12656
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 17052 12374 17080 12650
rect 17040 12368 17092 12374
rect 17144 12345 17172 12786
rect 17040 12310 17092 12316
rect 17130 12336 17186 12345
rect 17052 11762 17080 12310
rect 17130 12271 17186 12280
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 17040 11144 17092 11150
rect 17038 11112 17040 11121
rect 17092 11112 17094 11121
rect 17038 11047 17094 11056
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16580 10736 16632 10742
rect 16580 10678 16632 10684
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16868 10062 16896 10610
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 16592 9926 16620 9998
rect 16960 9994 16988 10950
rect 17144 10810 17172 12271
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 16948 9988 17000 9994
rect 16948 9930 17000 9936
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16304 9648 16356 9654
rect 16304 9590 16356 9596
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16408 8566 16436 9454
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 15844 5636 15896 5642
rect 15844 5578 15896 5584
rect 15842 5264 15898 5273
rect 15842 5199 15844 5208
rect 15896 5199 15898 5208
rect 15844 5170 15896 5176
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 15948 4622 15976 4762
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 16028 4616 16080 4622
rect 16028 4558 16080 4564
rect 15948 4264 15976 4558
rect 15856 4236 15976 4264
rect 15856 4146 15884 4236
rect 15934 4176 15990 4185
rect 15844 4140 15896 4146
rect 15934 4111 15990 4120
rect 15844 4082 15896 4088
rect 15844 3392 15896 3398
rect 15844 3334 15896 3340
rect 15856 3058 15884 3334
rect 15948 3126 15976 4111
rect 16040 3466 16068 4558
rect 16132 4554 16160 6734
rect 16408 5914 16436 8502
rect 16500 7818 16528 8978
rect 16592 8634 16620 9862
rect 17236 9654 17264 12786
rect 17328 12102 17356 13382
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17408 13252 17460 13258
rect 17408 13194 17460 13200
rect 17420 12850 17448 13194
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 17512 12442 17540 15098
rect 17604 12986 17632 15966
rect 17684 15904 17736 15910
rect 17684 15846 17736 15852
rect 17696 15570 17724 15846
rect 17684 15564 17736 15570
rect 17684 15506 17736 15512
rect 17788 15502 17816 16390
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 17684 15156 17736 15162
rect 17684 15098 17736 15104
rect 17696 13161 17724 15098
rect 17880 15094 17908 18022
rect 17992 17436 18300 17445
rect 17992 17434 17998 17436
rect 18054 17434 18078 17436
rect 18134 17434 18158 17436
rect 18214 17434 18238 17436
rect 18294 17434 18300 17436
rect 18054 17382 18056 17434
rect 18236 17382 18238 17434
rect 17992 17380 17998 17382
rect 18054 17380 18078 17382
rect 18134 17380 18158 17382
rect 18214 17380 18238 17382
rect 18294 17380 18300 17382
rect 17992 17371 18300 17380
rect 17960 17332 18012 17338
rect 17960 17274 18012 17280
rect 17972 16726 18000 17274
rect 17960 16720 18012 16726
rect 17960 16662 18012 16668
rect 17992 16348 18300 16357
rect 17992 16346 17998 16348
rect 18054 16346 18078 16348
rect 18134 16346 18158 16348
rect 18214 16346 18238 16348
rect 18294 16346 18300 16348
rect 18054 16294 18056 16346
rect 18236 16294 18238 16346
rect 17992 16292 17998 16294
rect 18054 16292 18078 16294
rect 18134 16292 18158 16294
rect 18214 16292 18238 16294
rect 18294 16292 18300 16294
rect 17992 16283 18300 16292
rect 17992 15260 18300 15269
rect 17992 15258 17998 15260
rect 18054 15258 18078 15260
rect 18134 15258 18158 15260
rect 18214 15258 18238 15260
rect 18294 15258 18300 15260
rect 18054 15206 18056 15258
rect 18236 15206 18238 15258
rect 17992 15204 17998 15206
rect 18054 15204 18078 15206
rect 18134 15204 18158 15206
rect 18214 15204 18238 15206
rect 18294 15204 18300 15206
rect 17992 15195 18300 15204
rect 17868 15088 17920 15094
rect 17868 15030 17920 15036
rect 17776 14952 17828 14958
rect 17776 14894 17828 14900
rect 17682 13152 17738 13161
rect 17682 13087 17738 13096
rect 17592 12980 17644 12986
rect 17592 12922 17644 12928
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17328 11898 17356 12038
rect 17420 11898 17448 12174
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17512 11218 17540 12378
rect 17592 11756 17644 11762
rect 17592 11698 17644 11704
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16488 7812 16540 7818
rect 16488 7754 16540 7760
rect 16592 7342 16620 8570
rect 16776 8362 16804 9522
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 16868 9042 16896 9318
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16776 7750 16804 8298
rect 16868 8022 16896 8978
rect 16948 8832 17000 8838
rect 16948 8774 17000 8780
rect 16960 8634 16988 8774
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 16856 8016 16908 8022
rect 16856 7958 16908 7964
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16776 7410 16804 7686
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 16592 7002 16620 7278
rect 16580 6996 16632 7002
rect 16580 6938 16632 6944
rect 16488 6384 16540 6390
rect 16488 6326 16540 6332
rect 16396 5908 16448 5914
rect 16396 5850 16448 5856
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 16316 5370 16344 5646
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 16500 4690 16528 6326
rect 16592 5710 16620 6938
rect 16764 6248 16816 6254
rect 16764 6190 16816 6196
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 16592 4690 16620 4762
rect 16488 4684 16540 4690
rect 16488 4626 16540 4632
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 16120 4548 16172 4554
rect 16120 4490 16172 4496
rect 16500 4486 16528 4626
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 16302 4176 16358 4185
rect 16120 4143 16172 4149
rect 16302 4111 16304 4120
rect 16120 4085 16172 4091
rect 16356 4111 16358 4120
rect 16028 3460 16080 3466
rect 16028 3402 16080 3408
rect 16132 3194 16160 4085
rect 16304 4082 16356 4088
rect 16684 4060 16712 6054
rect 16776 4826 16804 6190
rect 16868 5370 16896 7822
rect 16960 5710 16988 8366
rect 17144 8090 17172 9318
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 17052 7410 17080 7958
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 17052 6866 17080 7346
rect 17144 7274 17172 8026
rect 17236 7886 17264 9318
rect 17328 7954 17356 10610
rect 17604 10198 17632 11698
rect 17592 10192 17644 10198
rect 17592 10134 17644 10140
rect 17696 10044 17724 13087
rect 17788 12306 17816 14894
rect 17992 14172 18300 14181
rect 17992 14170 17998 14172
rect 18054 14170 18078 14172
rect 18134 14170 18158 14172
rect 18214 14170 18238 14172
rect 18294 14170 18300 14172
rect 18054 14118 18056 14170
rect 18236 14118 18238 14170
rect 17992 14116 17998 14118
rect 18054 14116 18078 14118
rect 18134 14116 18158 14118
rect 18214 14116 18238 14118
rect 18294 14116 18300 14118
rect 17992 14107 18300 14116
rect 17992 13084 18300 13093
rect 17992 13082 17998 13084
rect 18054 13082 18078 13084
rect 18134 13082 18158 13084
rect 18214 13082 18238 13084
rect 18294 13082 18300 13084
rect 18054 13030 18056 13082
rect 18236 13030 18238 13082
rect 17992 13028 17998 13030
rect 18054 13028 18078 13030
rect 18134 13028 18158 13030
rect 18214 13028 18238 13030
rect 18294 13028 18300 13030
rect 17992 13019 18300 13028
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 17868 12640 17920 12646
rect 17868 12582 17920 12588
rect 17880 12306 17908 12582
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 17868 12300 17920 12306
rect 17868 12242 17920 12248
rect 17776 12096 17828 12102
rect 18248 12084 18276 12718
rect 18340 12442 18368 18022
rect 18432 13802 18460 18362
rect 18420 13796 18472 13802
rect 18420 13738 18472 13744
rect 18524 12986 18552 18770
rect 18616 17105 18644 19382
rect 18696 18896 18748 18902
rect 18696 18838 18748 18844
rect 18602 17096 18658 17105
rect 18602 17031 18658 17040
rect 18616 16590 18644 17031
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18708 16522 18736 18838
rect 18800 17184 18828 19450
rect 18880 19440 18932 19446
rect 18880 19382 18932 19388
rect 18892 18970 18920 19382
rect 18880 18964 18932 18970
rect 18880 18906 18932 18912
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18892 17338 18920 18702
rect 19352 18426 19380 21014
rect 19444 20058 19472 21558
rect 20456 21554 20484 21927
rect 20732 21622 20760 21966
rect 22388 21690 22416 24200
rect 22652 21956 22704 21962
rect 22652 21898 22704 21904
rect 22664 21690 22692 21898
rect 22836 21888 22888 21894
rect 22836 21830 22888 21836
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 22376 21684 22428 21690
rect 22376 21626 22428 21632
rect 22652 21684 22704 21690
rect 22652 21626 22704 21632
rect 20720 21616 20772 21622
rect 20720 21558 20772 21564
rect 19708 21548 19760 21554
rect 19708 21490 19760 21496
rect 20260 21548 20312 21554
rect 20260 21490 20312 21496
rect 20444 21548 20496 21554
rect 20444 21490 20496 21496
rect 19522 21448 19578 21457
rect 19522 21383 19578 21392
rect 19536 21146 19564 21383
rect 19524 21140 19576 21146
rect 19524 21082 19576 21088
rect 19524 20936 19576 20942
rect 19524 20878 19576 20884
rect 19616 20936 19668 20942
rect 19616 20878 19668 20884
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 19432 19236 19484 19242
rect 19432 19178 19484 19184
rect 19444 18970 19472 19178
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19536 18834 19564 20878
rect 19628 20777 19656 20878
rect 19614 20768 19670 20777
rect 19614 20703 19670 20712
rect 19720 20618 19748 21490
rect 19800 20936 19852 20942
rect 20168 20936 20220 20942
rect 19852 20884 20116 20890
rect 19800 20878 20116 20884
rect 20168 20878 20220 20884
rect 19628 20590 19748 20618
rect 19812 20874 20116 20878
rect 19812 20868 20128 20874
rect 19812 20862 20076 20868
rect 19628 19378 19656 20590
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 19708 19372 19760 19378
rect 19708 19314 19760 19320
rect 19524 18828 19576 18834
rect 19524 18770 19576 18776
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19156 18148 19208 18154
rect 19156 18090 19208 18096
rect 18880 17332 18932 17338
rect 18880 17274 18932 17280
rect 19168 17270 19196 18090
rect 19156 17264 19208 17270
rect 19156 17206 19208 17212
rect 18880 17196 18932 17202
rect 18800 17156 18880 17184
rect 18880 17138 18932 17144
rect 19248 17196 19300 17202
rect 19248 17138 19300 17144
rect 18788 16652 18840 16658
rect 18788 16594 18840 16600
rect 18696 16516 18748 16522
rect 18696 16458 18748 16464
rect 18708 16250 18736 16458
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 18800 15162 18828 16594
rect 18788 15156 18840 15162
rect 18788 15098 18840 15104
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18708 14278 18736 14894
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 18512 12776 18564 12782
rect 18512 12718 18564 12724
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18248 12056 18368 12084
rect 17776 12038 17828 12044
rect 17788 11150 17816 12038
rect 17992 11996 18300 12005
rect 17992 11994 17998 11996
rect 18054 11994 18078 11996
rect 18134 11994 18158 11996
rect 18214 11994 18238 11996
rect 18294 11994 18300 11996
rect 18054 11942 18056 11994
rect 18236 11942 18238 11994
rect 17992 11940 17998 11942
rect 18054 11940 18078 11942
rect 18134 11940 18158 11942
rect 18214 11940 18238 11942
rect 18294 11940 18300 11942
rect 17992 11931 18300 11940
rect 17866 11792 17922 11801
rect 17866 11727 17922 11736
rect 17880 11694 17908 11727
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17880 10996 17908 11630
rect 18340 11354 18368 12056
rect 18328 11348 18380 11354
rect 18328 11290 18380 11296
rect 18524 11218 18552 12718
rect 18616 12714 18644 13738
rect 18604 12708 18656 12714
rect 18604 12650 18656 12656
rect 18708 11558 18736 14214
rect 18800 13326 18828 14962
rect 18892 14550 18920 17138
rect 18972 16108 19024 16114
rect 18972 16050 19024 16056
rect 18880 14544 18932 14550
rect 18880 14486 18932 14492
rect 18788 13320 18840 13326
rect 18786 13288 18788 13297
rect 18840 13288 18842 13297
rect 18786 13223 18842 13232
rect 18800 12782 18828 13223
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18512 11212 18564 11218
rect 18432 11172 18512 11200
rect 18432 11082 18460 11172
rect 18512 11154 18564 11160
rect 18420 11076 18472 11082
rect 18420 11018 18472 11024
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18788 11076 18840 11082
rect 18788 11018 18840 11024
rect 17604 10016 17724 10044
rect 17788 10968 17908 10996
rect 17604 9674 17632 10016
rect 17788 9897 17816 10968
rect 17992 10908 18300 10917
rect 17992 10906 17998 10908
rect 18054 10906 18078 10908
rect 18134 10906 18158 10908
rect 18214 10906 18238 10908
rect 18294 10906 18300 10908
rect 18054 10854 18056 10906
rect 18236 10854 18238 10906
rect 17992 10852 17998 10854
rect 18054 10852 18078 10854
rect 18134 10852 18158 10854
rect 18214 10852 18238 10854
rect 18294 10852 18300 10854
rect 17992 10843 18300 10852
rect 18432 10810 18460 11018
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18064 10266 18092 10406
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 17774 9888 17830 9897
rect 17774 9823 17830 9832
rect 17604 9654 17724 9674
rect 17604 9648 17736 9654
rect 17604 9646 17684 9648
rect 17684 9590 17736 9596
rect 17880 9178 17908 10202
rect 18340 10062 18368 10406
rect 18524 10062 18552 11018
rect 18604 10668 18656 10674
rect 18604 10610 18656 10616
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18432 9908 18460 9998
rect 18340 9880 18460 9908
rect 17992 9820 18300 9829
rect 17992 9818 17998 9820
rect 18054 9818 18078 9820
rect 18134 9818 18158 9820
rect 18214 9818 18238 9820
rect 18294 9818 18300 9820
rect 18054 9766 18056 9818
rect 18236 9766 18238 9818
rect 17992 9764 17998 9766
rect 18054 9764 18078 9766
rect 18134 9764 18158 9766
rect 18214 9764 18238 9766
rect 18294 9764 18300 9766
rect 17992 9755 18300 9764
rect 17958 9688 18014 9697
rect 17958 9623 18014 9632
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17500 8492 17552 8498
rect 17420 8452 17500 8480
rect 17420 8022 17448 8452
rect 17500 8434 17552 8440
rect 17408 8016 17460 8022
rect 17408 7958 17460 7964
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17420 7886 17448 7958
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17420 7478 17448 7822
rect 17604 7478 17632 8978
rect 17972 8922 18000 9623
rect 18340 9518 18368 9880
rect 18420 9580 18472 9586
rect 18524 9568 18552 9998
rect 18472 9540 18552 9568
rect 18420 9522 18472 9528
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 17880 8894 18000 8922
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17880 8838 17908 8894
rect 18064 8838 18092 8910
rect 18328 8900 18380 8906
rect 18328 8842 18380 8848
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 17880 8616 17908 8774
rect 17992 8732 18300 8741
rect 17992 8730 17998 8732
rect 18054 8730 18078 8732
rect 18134 8730 18158 8732
rect 18214 8730 18238 8732
rect 18294 8730 18300 8732
rect 18054 8678 18056 8730
rect 18236 8678 18238 8730
rect 17992 8676 17998 8678
rect 18054 8676 18078 8678
rect 18134 8676 18158 8678
rect 18214 8676 18238 8678
rect 18294 8676 18300 8678
rect 17992 8667 18300 8676
rect 18340 8634 18368 8842
rect 18328 8628 18380 8634
rect 17880 8588 18000 8616
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17788 7886 17816 8366
rect 17972 8362 18000 8588
rect 18328 8570 18380 8576
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 18156 7818 18184 8434
rect 18432 8090 18460 9522
rect 18616 9382 18644 10610
rect 18708 10266 18736 10610
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18616 9110 18644 9318
rect 18604 9104 18656 9110
rect 18604 9046 18656 9052
rect 18708 8974 18736 10202
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 18708 7886 18736 8910
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18144 7812 18196 7818
rect 18196 7772 18368 7800
rect 18144 7754 18196 7760
rect 17992 7644 18300 7653
rect 17992 7642 17998 7644
rect 18054 7642 18078 7644
rect 18134 7642 18158 7644
rect 18214 7642 18238 7644
rect 18294 7642 18300 7644
rect 18054 7590 18056 7642
rect 18236 7590 18238 7642
rect 17992 7588 17998 7590
rect 18054 7588 18078 7590
rect 18134 7588 18158 7590
rect 18214 7588 18238 7590
rect 18294 7588 18300 7590
rect 17992 7579 18300 7588
rect 17408 7472 17460 7478
rect 17408 7414 17460 7420
rect 17592 7472 17644 7478
rect 17592 7414 17644 7420
rect 18340 7410 18368 7772
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 17132 7268 17184 7274
rect 17132 7210 17184 7216
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 18328 6860 18380 6866
rect 18328 6802 18380 6808
rect 17992 6556 18300 6565
rect 17992 6554 17998 6556
rect 18054 6554 18078 6556
rect 18134 6554 18158 6556
rect 18214 6554 18238 6556
rect 18294 6554 18300 6556
rect 18054 6502 18056 6554
rect 18236 6502 18238 6554
rect 17992 6500 17998 6502
rect 18054 6500 18078 6502
rect 18134 6500 18158 6502
rect 18214 6500 18238 6502
rect 18294 6500 18300 6502
rect 17992 6491 18300 6500
rect 18340 6458 18368 6802
rect 18694 6760 18750 6769
rect 18694 6695 18750 6704
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 17132 6316 17184 6322
rect 17408 6316 17460 6322
rect 17132 6258 17184 6264
rect 17328 6276 17408 6304
rect 17144 5778 17172 6258
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 17328 5710 17356 6276
rect 17408 6258 17460 6264
rect 18236 6248 18288 6254
rect 18236 6190 18288 6196
rect 17500 6180 17552 6186
rect 17500 6122 17552 6128
rect 17512 5778 17540 6122
rect 18248 5778 18276 6190
rect 17500 5772 17552 5778
rect 17500 5714 17552 5720
rect 18236 5772 18288 5778
rect 18236 5714 18288 5720
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16960 5302 16988 5646
rect 16948 5296 17000 5302
rect 16948 5238 17000 5244
rect 17328 5030 17356 5646
rect 17512 5302 17540 5714
rect 17992 5468 18300 5477
rect 17992 5466 17998 5468
rect 18054 5466 18078 5468
rect 18134 5466 18158 5468
rect 18214 5466 18238 5468
rect 18294 5466 18300 5468
rect 18054 5414 18056 5466
rect 18236 5414 18238 5466
rect 17992 5412 17998 5414
rect 18054 5412 18078 5414
rect 18134 5412 18158 5414
rect 18214 5412 18238 5414
rect 18294 5412 18300 5414
rect 17992 5403 18300 5412
rect 17500 5296 17552 5302
rect 17500 5238 17552 5244
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 18328 5228 18380 5234
rect 18328 5170 18380 5176
rect 18420 5228 18472 5234
rect 18420 5170 18472 5176
rect 17500 5092 17552 5098
rect 17500 5034 17552 5040
rect 17316 5024 17368 5030
rect 17316 4966 17368 4972
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 17224 4480 17276 4486
rect 17224 4422 17276 4428
rect 16684 4032 16804 4060
rect 16776 3398 16804 4032
rect 16764 3392 16816 3398
rect 16764 3334 16816 3340
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 15936 3120 15988 3126
rect 15936 3062 15988 3068
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 15752 2644 15804 2650
rect 15752 2586 15804 2592
rect 16580 2508 16632 2514
rect 16580 2450 16632 2456
rect 16592 898 16620 2450
rect 16776 2378 16804 3334
rect 17236 3058 17264 4422
rect 17328 4146 17356 4966
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17328 3058 17356 3878
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17420 3194 17448 3334
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 17052 2650 17080 2994
rect 17132 2916 17184 2922
rect 17132 2858 17184 2864
rect 17040 2644 17092 2650
rect 17040 2586 17092 2592
rect 17144 2446 17172 2858
rect 17420 2854 17448 3130
rect 17512 3058 17540 5034
rect 18156 4826 18184 5170
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 17592 3732 17644 3738
rect 17592 3674 17644 3680
rect 17776 3732 17828 3738
rect 17776 3674 17828 3680
rect 17604 3058 17632 3674
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17592 3052 17644 3058
rect 17592 2994 17644 3000
rect 17788 2854 17816 3674
rect 17880 3670 17908 4558
rect 17992 4380 18300 4389
rect 17992 4378 17998 4380
rect 18054 4378 18078 4380
rect 18134 4378 18158 4380
rect 18214 4378 18238 4380
rect 18294 4378 18300 4380
rect 18054 4326 18056 4378
rect 18236 4326 18238 4378
rect 17992 4324 17998 4326
rect 18054 4324 18078 4326
rect 18134 4324 18158 4326
rect 18214 4324 18238 4326
rect 18294 4324 18300 4326
rect 17992 4315 18300 4324
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 17972 4078 18000 4218
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 17972 3738 18000 4014
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 17868 3664 17920 3670
rect 17868 3606 17920 3612
rect 17880 2990 17908 3606
rect 18340 3505 18368 5170
rect 18432 5137 18460 5170
rect 18418 5128 18474 5137
rect 18418 5063 18474 5072
rect 18420 4752 18472 4758
rect 18420 4694 18472 4700
rect 18432 3534 18460 4694
rect 18708 4214 18736 6695
rect 18800 6458 18828 11018
rect 18892 9518 18920 14486
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18892 6662 18920 9454
rect 18984 8634 19012 16050
rect 19064 16040 19116 16046
rect 19062 16008 19064 16017
rect 19116 16008 19118 16017
rect 19062 15943 19118 15952
rect 19156 15972 19208 15978
rect 19156 15914 19208 15920
rect 19064 14476 19116 14482
rect 19064 14418 19116 14424
rect 19076 12850 19104 14418
rect 19168 12889 19196 15914
rect 19260 15570 19288 17138
rect 19430 16552 19486 16561
rect 19430 16487 19486 16496
rect 19444 15638 19472 16487
rect 19536 16454 19564 18770
rect 19720 17338 19748 19314
rect 19812 18630 19840 20862
rect 20076 20810 20128 20816
rect 20180 20330 20208 20878
rect 20272 20806 20300 21490
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20628 20936 20680 20942
rect 20732 20890 20760 21422
rect 20833 21244 21141 21253
rect 20833 21242 20839 21244
rect 20895 21242 20919 21244
rect 20975 21242 20999 21244
rect 21055 21242 21079 21244
rect 21135 21242 21141 21244
rect 20895 21190 20897 21242
rect 21077 21190 21079 21242
rect 20833 21188 20839 21190
rect 20895 21188 20919 21190
rect 20975 21188 20999 21190
rect 21055 21188 21079 21190
rect 21135 21188 21141 21190
rect 20833 21179 21141 21188
rect 20680 20884 20760 20890
rect 20628 20878 20760 20884
rect 20640 20862 20760 20878
rect 20260 20800 20312 20806
rect 20260 20742 20312 20748
rect 20272 20534 20300 20742
rect 20732 20602 20760 20862
rect 21914 20904 21970 20913
rect 21914 20839 21916 20848
rect 21968 20839 21970 20848
rect 21916 20810 21968 20816
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 20260 20528 20312 20534
rect 20260 20470 20312 20476
rect 20168 20324 20220 20330
rect 20168 20266 20220 20272
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 20088 19378 20116 19790
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19800 18624 19852 18630
rect 19800 18566 19852 18572
rect 19800 18352 19852 18358
rect 19800 18294 19852 18300
rect 19616 17332 19668 17338
rect 19616 17274 19668 17280
rect 19708 17332 19760 17338
rect 19708 17274 19760 17280
rect 19524 16448 19576 16454
rect 19524 16390 19576 16396
rect 19628 16266 19656 17274
rect 19812 17202 19840 18294
rect 19892 18284 19944 18290
rect 19892 18226 19944 18232
rect 19904 18057 19932 18226
rect 19890 18048 19946 18057
rect 19890 17983 19946 17992
rect 19800 17196 19852 17202
rect 19800 17138 19852 17144
rect 19892 16516 19944 16522
rect 19892 16458 19944 16464
rect 19536 16238 19656 16266
rect 19432 15632 19484 15638
rect 19432 15574 19484 15580
rect 19248 15564 19300 15570
rect 19300 15524 19380 15552
rect 19248 15506 19300 15512
rect 19352 14278 19380 15524
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19248 13864 19300 13870
rect 19248 13806 19300 13812
rect 19260 13530 19288 13806
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19248 13252 19300 13258
rect 19248 13194 19300 13200
rect 19154 12880 19210 12889
rect 19064 12844 19116 12850
rect 19154 12815 19210 12824
rect 19064 12786 19116 12792
rect 19076 12170 19104 12786
rect 19156 12708 19208 12714
rect 19156 12650 19208 12656
rect 19064 12164 19116 12170
rect 19064 12106 19116 12112
rect 19076 11082 19104 12106
rect 19064 11076 19116 11082
rect 19064 11018 19116 11024
rect 19168 10130 19196 12650
rect 19260 11014 19288 13194
rect 19352 12442 19380 13330
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19338 12336 19394 12345
rect 19338 12271 19340 12280
rect 19392 12271 19394 12280
rect 19340 12242 19392 12248
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 19444 10742 19472 14962
rect 19536 13462 19564 16238
rect 19904 15978 19932 16458
rect 19892 15972 19944 15978
rect 19892 15914 19944 15920
rect 19708 15156 19760 15162
rect 19708 15098 19760 15104
rect 19616 14272 19668 14278
rect 19616 14214 19668 14220
rect 19628 13462 19656 14214
rect 19524 13456 19576 13462
rect 19524 13398 19576 13404
rect 19616 13456 19668 13462
rect 19616 13398 19668 13404
rect 19524 12436 19576 12442
rect 19524 12378 19576 12384
rect 19536 11082 19564 12378
rect 19628 12374 19656 13398
rect 19720 12442 19748 15098
rect 19996 14618 20024 18702
rect 20088 18290 20116 19314
rect 20168 18624 20220 18630
rect 20168 18566 20220 18572
rect 20076 18284 20128 18290
rect 20076 18226 20128 18232
rect 20088 14958 20116 18226
rect 20180 15502 20208 18566
rect 20272 18358 20300 20470
rect 22296 20466 22324 21626
rect 22652 21004 22704 21010
rect 22652 20946 22704 20952
rect 22664 20602 22692 20946
rect 22652 20596 22704 20602
rect 22652 20538 22704 20544
rect 22848 20466 22876 21830
rect 23673 21788 23981 21797
rect 23673 21786 23679 21788
rect 23735 21786 23759 21788
rect 23815 21786 23839 21788
rect 23895 21786 23919 21788
rect 23975 21786 23981 21788
rect 23735 21734 23737 21786
rect 23917 21734 23919 21786
rect 23673 21732 23679 21734
rect 23735 21732 23759 21734
rect 23815 21732 23839 21734
rect 23895 21732 23919 21734
rect 23975 21732 23981 21734
rect 23673 21723 23981 21732
rect 23673 20700 23981 20709
rect 23673 20698 23679 20700
rect 23735 20698 23759 20700
rect 23815 20698 23839 20700
rect 23895 20698 23919 20700
rect 23975 20698 23981 20700
rect 23735 20646 23737 20698
rect 23917 20646 23919 20698
rect 23673 20644 23679 20646
rect 23735 20644 23759 20646
rect 23815 20644 23839 20646
rect 23895 20644 23919 20646
rect 23975 20644 23981 20646
rect 23673 20635 23981 20644
rect 22008 20460 22060 20466
rect 22008 20402 22060 20408
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 22836 20460 22888 20466
rect 22836 20402 22888 20408
rect 20536 20324 20588 20330
rect 20536 20266 20588 20272
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20260 18352 20312 18358
rect 20260 18294 20312 18300
rect 20456 17882 20484 18702
rect 20444 17876 20496 17882
rect 20444 17818 20496 17824
rect 20352 16720 20404 16726
rect 20352 16662 20404 16668
rect 20260 16108 20312 16114
rect 20260 16050 20312 16056
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19800 13932 19852 13938
rect 19800 13874 19852 13880
rect 19708 12436 19760 12442
rect 19708 12378 19760 12384
rect 19616 12368 19668 12374
rect 19616 12310 19668 12316
rect 19812 12306 19840 13874
rect 19800 12300 19852 12306
rect 19800 12242 19852 12248
rect 19800 11620 19852 11626
rect 19800 11562 19852 11568
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19524 11076 19576 11082
rect 19524 11018 19576 11024
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 19338 10568 19394 10577
rect 19338 10503 19394 10512
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 19168 9110 19196 10066
rect 19260 9518 19288 10406
rect 19352 9586 19380 10503
rect 19444 10062 19472 10678
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19156 9104 19208 9110
rect 19156 9046 19208 9052
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 18984 8401 19012 8570
rect 19064 8560 19116 8566
rect 19064 8502 19116 8508
rect 18970 8392 19026 8401
rect 18970 8327 19026 8336
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 18984 6866 19012 7346
rect 18972 6860 19024 6866
rect 18972 6802 19024 6808
rect 18880 6656 18932 6662
rect 18880 6598 18932 6604
rect 18788 6452 18840 6458
rect 18788 6394 18840 6400
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18800 5914 18828 6258
rect 18984 6186 19012 6802
rect 19076 6798 19104 8502
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 19168 7410 19196 8434
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 19168 6746 19196 7346
rect 19352 6798 19380 9522
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19444 8498 19472 9318
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 19536 8294 19564 11018
rect 19616 10464 19668 10470
rect 19616 10406 19668 10412
rect 19628 9110 19656 10406
rect 19616 9104 19668 9110
rect 19616 9046 19668 9052
rect 19628 8566 19656 9046
rect 19616 8560 19668 8566
rect 19616 8502 19668 8508
rect 19524 8288 19576 8294
rect 19524 8230 19576 8236
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 19432 7744 19484 7750
rect 19432 7686 19484 7692
rect 19444 6798 19472 7686
rect 19628 6798 19656 7822
rect 19720 7342 19748 11494
rect 19812 11150 19840 11562
rect 19800 11144 19852 11150
rect 19800 11086 19852 11092
rect 19800 8900 19852 8906
rect 19800 8842 19852 8848
rect 19708 7336 19760 7342
rect 19708 7278 19760 7284
rect 19340 6792 19392 6798
rect 19168 6730 19288 6746
rect 19340 6734 19392 6740
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19168 6724 19300 6730
rect 19168 6718 19248 6724
rect 19168 6254 19196 6718
rect 19248 6666 19300 6672
rect 19444 6254 19472 6734
rect 19628 6390 19656 6734
rect 19616 6384 19668 6390
rect 19616 6326 19668 6332
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 18972 6180 19024 6186
rect 18972 6122 19024 6128
rect 18788 5908 18840 5914
rect 18788 5850 18840 5856
rect 19628 5710 19656 6326
rect 19812 5778 19840 8842
rect 19904 8634 19932 14350
rect 20272 14074 20300 16050
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 19996 11898 20024 13874
rect 20088 12986 20116 13874
rect 20364 13190 20392 16662
rect 20456 16250 20484 17818
rect 20444 16244 20496 16250
rect 20444 16186 20496 16192
rect 20548 15910 20576 20266
rect 20833 20156 21141 20165
rect 20833 20154 20839 20156
rect 20895 20154 20919 20156
rect 20975 20154 20999 20156
rect 21055 20154 21079 20156
rect 21135 20154 21141 20156
rect 20895 20102 20897 20154
rect 21077 20102 21079 20154
rect 20833 20100 20839 20102
rect 20895 20100 20919 20102
rect 20975 20100 20999 20102
rect 21055 20100 21079 20102
rect 21135 20100 21141 20102
rect 20833 20091 21141 20100
rect 22020 19922 22048 20402
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22284 19984 22336 19990
rect 22284 19926 22336 19932
rect 22008 19916 22060 19922
rect 22008 19858 22060 19864
rect 22020 19514 22048 19858
rect 22008 19508 22060 19514
rect 22008 19450 22060 19456
rect 21180 19304 21232 19310
rect 21180 19246 21232 19252
rect 20833 19068 21141 19077
rect 20833 19066 20839 19068
rect 20895 19066 20919 19068
rect 20975 19066 20999 19068
rect 21055 19066 21079 19068
rect 21135 19066 21141 19068
rect 20895 19014 20897 19066
rect 21077 19014 21079 19066
rect 20833 19012 20839 19014
rect 20895 19012 20919 19014
rect 20975 19012 20999 19014
rect 21055 19012 21079 19014
rect 21135 19012 21141 19014
rect 20833 19003 21141 19012
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20732 16250 20760 18158
rect 20833 17980 21141 17989
rect 20833 17978 20839 17980
rect 20895 17978 20919 17980
rect 20975 17978 20999 17980
rect 21055 17978 21079 17980
rect 21135 17978 21141 17980
rect 20895 17926 20897 17978
rect 21077 17926 21079 17978
rect 20833 17924 20839 17926
rect 20895 17924 20919 17926
rect 20975 17924 20999 17926
rect 21055 17924 21079 17926
rect 21135 17924 21141 17926
rect 20833 17915 21141 17924
rect 21192 17066 21220 19246
rect 22296 19174 22324 19926
rect 22284 19168 22336 19174
rect 22284 19110 22336 19116
rect 22296 17678 22324 19110
rect 22572 17882 22600 20334
rect 23673 19612 23981 19621
rect 23673 19610 23679 19612
rect 23735 19610 23759 19612
rect 23815 19610 23839 19612
rect 23895 19610 23919 19612
rect 23975 19610 23981 19612
rect 23735 19558 23737 19610
rect 23917 19558 23919 19610
rect 23673 19556 23679 19558
rect 23735 19556 23759 19558
rect 23815 19556 23839 19558
rect 23895 19556 23919 19558
rect 23975 19556 23981 19558
rect 23673 19547 23981 19556
rect 23673 18524 23981 18533
rect 23673 18522 23679 18524
rect 23735 18522 23759 18524
rect 23815 18522 23839 18524
rect 23895 18522 23919 18524
rect 23975 18522 23981 18524
rect 23735 18470 23737 18522
rect 23917 18470 23919 18522
rect 23673 18468 23679 18470
rect 23735 18468 23759 18470
rect 23815 18468 23839 18470
rect 23895 18468 23919 18470
rect 23975 18468 23981 18470
rect 23673 18459 23981 18468
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22192 17672 22244 17678
rect 22192 17614 22244 17620
rect 22284 17672 22336 17678
rect 22284 17614 22336 17620
rect 22376 17672 22428 17678
rect 22376 17614 22428 17620
rect 21824 17128 21876 17134
rect 21824 17070 21876 17076
rect 21180 17060 21232 17066
rect 21180 17002 21232 17008
rect 21272 17060 21324 17066
rect 21272 17002 21324 17008
rect 20833 16892 21141 16901
rect 20833 16890 20839 16892
rect 20895 16890 20919 16892
rect 20975 16890 20999 16892
rect 21055 16890 21079 16892
rect 21135 16890 21141 16892
rect 20895 16838 20897 16890
rect 21077 16838 21079 16890
rect 20833 16836 20839 16838
rect 20895 16836 20919 16838
rect 20975 16836 20999 16838
rect 21055 16836 21079 16838
rect 21135 16836 21141 16838
rect 20833 16827 21141 16836
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20444 15088 20496 15094
rect 20444 15030 20496 15036
rect 20456 14550 20484 15030
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20444 14544 20496 14550
rect 20444 14486 20496 14492
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 20352 13184 20404 13190
rect 20352 13126 20404 13132
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 20364 12646 20392 13126
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 20352 12232 20404 12238
rect 20352 12174 20404 12180
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 20088 11354 20116 12174
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 20076 11348 20128 11354
rect 20076 11290 20128 11296
rect 20180 9926 20208 11630
rect 20260 11620 20312 11626
rect 20260 11562 20312 11568
rect 20272 10062 20300 11562
rect 20364 11354 20392 12174
rect 20456 11694 20484 14282
rect 20548 14074 20576 14894
rect 20536 14068 20588 14074
rect 20536 14010 20588 14016
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20548 11762 20576 12038
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20444 11688 20496 11694
rect 20444 11630 20496 11636
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20456 10577 20484 11494
rect 20442 10568 20498 10577
rect 20442 10503 20498 10512
rect 20260 10056 20312 10062
rect 20260 9998 20312 10004
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 19892 8424 19944 8430
rect 19892 8366 19944 8372
rect 19904 5914 19932 8366
rect 20180 7818 20208 9862
rect 20272 8498 20300 9998
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20260 8492 20312 8498
rect 20260 8434 20312 8440
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20272 7954 20300 8434
rect 20364 8294 20392 8434
rect 20352 8288 20404 8294
rect 20352 8230 20404 8236
rect 20456 7970 20484 9454
rect 20548 9110 20576 11698
rect 20640 10146 20668 16050
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20732 15434 20760 15846
rect 20833 15804 21141 15813
rect 20833 15802 20839 15804
rect 20895 15802 20919 15804
rect 20975 15802 20999 15804
rect 21055 15802 21079 15804
rect 21135 15802 21141 15804
rect 20895 15750 20897 15802
rect 21077 15750 21079 15802
rect 20833 15748 20839 15750
rect 20895 15748 20919 15750
rect 20975 15748 20999 15750
rect 21055 15748 21079 15750
rect 21135 15748 21141 15750
rect 20833 15739 21141 15748
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20732 14550 20760 15370
rect 21192 15162 21220 16594
rect 21284 15366 21312 17002
rect 21456 16448 21508 16454
rect 21456 16390 21508 16396
rect 21272 15360 21324 15366
rect 21272 15302 21324 15308
rect 21180 15156 21232 15162
rect 21180 15098 21232 15104
rect 21192 14822 21220 15098
rect 21180 14816 21232 14822
rect 21180 14758 21232 14764
rect 20833 14716 21141 14725
rect 20833 14714 20839 14716
rect 20895 14714 20919 14716
rect 20975 14714 20999 14716
rect 21055 14714 21079 14716
rect 21135 14714 21141 14716
rect 20895 14662 20897 14714
rect 21077 14662 21079 14714
rect 20833 14660 20839 14662
rect 20895 14660 20919 14662
rect 20975 14660 20999 14662
rect 21055 14660 21079 14662
rect 21135 14660 21141 14662
rect 20833 14651 21141 14660
rect 21192 14600 21220 14758
rect 21100 14572 21220 14600
rect 20720 14544 20772 14550
rect 20720 14486 20772 14492
rect 20732 13410 20760 14486
rect 20996 14476 21048 14482
rect 20996 14418 21048 14424
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20916 13802 20944 14214
rect 21008 13802 21036 14418
rect 21100 13818 21128 14572
rect 21284 13954 21312 15302
rect 21468 14346 21496 16390
rect 21836 15706 21864 17070
rect 21824 15700 21876 15706
rect 21824 15642 21876 15648
rect 22100 15496 22152 15502
rect 22100 15438 22152 15444
rect 21640 15428 21692 15434
rect 21640 15370 21692 15376
rect 21548 14884 21600 14890
rect 21548 14826 21600 14832
rect 21456 14340 21508 14346
rect 21456 14282 21508 14288
rect 21192 13938 21312 13954
rect 21180 13932 21312 13938
rect 21232 13926 21312 13932
rect 21180 13874 21232 13880
rect 20904 13796 20956 13802
rect 20904 13738 20956 13744
rect 20996 13796 21048 13802
rect 21100 13790 21220 13818
rect 20996 13738 21048 13744
rect 20833 13628 21141 13637
rect 20833 13626 20839 13628
rect 20895 13626 20919 13628
rect 20975 13626 20999 13628
rect 21055 13626 21079 13628
rect 21135 13626 21141 13628
rect 20895 13574 20897 13626
rect 21077 13574 21079 13626
rect 20833 13572 20839 13574
rect 20895 13572 20919 13574
rect 20975 13572 20999 13574
rect 21055 13572 21079 13574
rect 21135 13572 21141 13574
rect 20833 13563 21141 13572
rect 20732 13394 20852 13410
rect 20732 13388 20864 13394
rect 20732 13382 20812 13388
rect 20812 13330 20864 13336
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20732 12238 20760 13262
rect 20833 12540 21141 12549
rect 20833 12538 20839 12540
rect 20895 12538 20919 12540
rect 20975 12538 20999 12540
rect 21055 12538 21079 12540
rect 21135 12538 21141 12540
rect 20895 12486 20897 12538
rect 21077 12486 21079 12538
rect 20833 12484 20839 12486
rect 20895 12484 20919 12486
rect 20975 12484 20999 12486
rect 21055 12484 21079 12486
rect 21135 12484 21141 12486
rect 20833 12475 21141 12484
rect 21192 12424 21220 13790
rect 21272 13796 21324 13802
rect 21272 13738 21324 13744
rect 20824 12396 21220 12424
rect 21284 12434 21312 13738
rect 21284 12406 21404 12434
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 20824 11642 20852 12396
rect 21272 12368 21324 12374
rect 21086 12336 21142 12345
rect 21272 12310 21324 12316
rect 21086 12271 21088 12280
rect 21140 12271 21142 12280
rect 21088 12242 21140 12248
rect 21180 12232 21232 12238
rect 21180 12174 21232 12180
rect 20732 11614 20852 11642
rect 20732 10470 20760 11614
rect 20833 11452 21141 11461
rect 20833 11450 20839 11452
rect 20895 11450 20919 11452
rect 20975 11450 20999 11452
rect 21055 11450 21079 11452
rect 21135 11450 21141 11452
rect 20895 11398 20897 11450
rect 21077 11398 21079 11450
rect 20833 11396 20839 11398
rect 20895 11396 20919 11398
rect 20975 11396 20999 11398
rect 21055 11396 21079 11398
rect 21135 11396 21141 11398
rect 20833 11387 21141 11396
rect 21192 10674 21220 12174
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 20720 10464 20772 10470
rect 20720 10406 20772 10412
rect 20732 10248 20760 10406
rect 20833 10364 21141 10373
rect 20833 10362 20839 10364
rect 20895 10362 20919 10364
rect 20975 10362 20999 10364
rect 21055 10362 21079 10364
rect 21135 10362 21141 10364
rect 20895 10310 20897 10362
rect 21077 10310 21079 10362
rect 20833 10308 20839 10310
rect 20895 10308 20919 10310
rect 20975 10308 20999 10310
rect 21055 10308 21079 10310
rect 21135 10308 21141 10310
rect 20833 10299 21141 10308
rect 20732 10220 20852 10248
rect 20640 10118 20760 10146
rect 20824 10130 20852 10220
rect 20628 10056 20680 10062
rect 20628 9998 20680 10004
rect 20640 9586 20668 9998
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20536 9104 20588 9110
rect 20536 9046 20588 9052
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 20548 8090 20576 8910
rect 20640 8566 20668 9522
rect 20732 8634 20760 10118
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20824 9586 20852 10066
rect 21088 10056 21140 10062
rect 21088 9998 21140 10004
rect 21100 9722 21128 9998
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 21192 9654 21220 10610
rect 21284 10452 21312 12310
rect 21376 11762 21404 12406
rect 21468 12374 21496 14282
rect 21560 12434 21588 14826
rect 21652 14414 21680 15370
rect 21732 15020 21784 15026
rect 21732 14962 21784 14968
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21652 12850 21680 14350
rect 21640 12844 21692 12850
rect 21640 12786 21692 12792
rect 21560 12406 21680 12434
rect 21456 12368 21508 12374
rect 21456 12310 21508 12316
rect 21548 12368 21600 12374
rect 21548 12310 21600 12316
rect 21456 12232 21508 12238
rect 21560 12220 21588 12310
rect 21508 12192 21588 12220
rect 21456 12174 21508 12180
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21376 11626 21404 11698
rect 21364 11620 21416 11626
rect 21364 11562 21416 11568
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21376 10810 21404 11086
rect 21364 10804 21416 10810
rect 21364 10746 21416 10752
rect 21284 10424 21496 10452
rect 21364 10056 21416 10062
rect 21364 9998 21416 10004
rect 21180 9648 21232 9654
rect 21180 9590 21232 9596
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 21180 9512 21232 9518
rect 21180 9454 21232 9460
rect 20833 9276 21141 9285
rect 20833 9274 20839 9276
rect 20895 9274 20919 9276
rect 20975 9274 20999 9276
rect 21055 9274 21079 9276
rect 21135 9274 21141 9276
rect 20895 9222 20897 9274
rect 21077 9222 21079 9274
rect 20833 9220 20839 9222
rect 20895 9220 20919 9222
rect 20975 9220 20999 9222
rect 21055 9220 21079 9222
rect 21135 9220 21141 9222
rect 20833 9211 21141 9220
rect 20996 9172 21048 9178
rect 20996 9114 21048 9120
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 20720 8628 20772 8634
rect 20720 8570 20772 8576
rect 20628 8560 20680 8566
rect 20628 8502 20680 8508
rect 20536 8084 20588 8090
rect 20536 8026 20588 8032
rect 20260 7948 20312 7954
rect 20456 7942 20576 7970
rect 20260 7890 20312 7896
rect 19984 7812 20036 7818
rect 19984 7754 20036 7760
rect 20168 7812 20220 7818
rect 20168 7754 20220 7760
rect 19996 6322 20024 7754
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 20444 7336 20496 7342
rect 20444 7278 20496 7284
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 19892 5908 19944 5914
rect 19892 5850 19944 5856
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 19996 5370 20024 6258
rect 20168 6248 20220 6254
rect 20168 6190 20220 6196
rect 20180 5846 20208 6190
rect 20076 5840 20128 5846
rect 20076 5782 20128 5788
rect 20168 5840 20220 5846
rect 20168 5782 20220 5788
rect 19248 5364 19300 5370
rect 19248 5306 19300 5312
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 19260 5273 19288 5306
rect 19246 5264 19302 5273
rect 19246 5199 19302 5208
rect 19800 5092 19852 5098
rect 19800 5034 19852 5040
rect 18696 4208 18748 4214
rect 18696 4150 18748 4156
rect 19812 4146 19840 5034
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19800 4140 19852 4146
rect 19800 4082 19852 4088
rect 18880 4072 18932 4078
rect 18880 4014 18932 4020
rect 18420 3528 18472 3534
rect 18326 3496 18382 3505
rect 18420 3470 18472 3476
rect 18326 3431 18382 3440
rect 18892 3398 18920 4014
rect 18880 3392 18932 3398
rect 18880 3334 18932 3340
rect 17992 3292 18300 3301
rect 17992 3290 17998 3292
rect 18054 3290 18078 3292
rect 18134 3290 18158 3292
rect 18214 3290 18238 3292
rect 18294 3290 18300 3292
rect 18054 3238 18056 3290
rect 18236 3238 18238 3290
rect 17992 3236 17998 3238
rect 18054 3236 18078 3238
rect 18134 3236 18158 3238
rect 18214 3236 18238 3238
rect 18294 3236 18300 3238
rect 17992 3227 18300 3236
rect 18892 3058 18920 3334
rect 19260 3058 19288 4082
rect 19536 3126 19564 4082
rect 19524 3120 19576 3126
rect 19524 3062 19576 3068
rect 19812 3058 19840 4082
rect 20088 3602 20116 5782
rect 20272 5234 20300 7278
rect 20456 6390 20484 7278
rect 20548 6662 20576 7942
rect 20640 6798 20668 8502
rect 20824 8378 20852 8978
rect 21008 8566 21036 9114
rect 21088 9104 21140 9110
rect 21088 9046 21140 9052
rect 21100 8974 21128 9046
rect 21088 8968 21140 8974
rect 21088 8910 21140 8916
rect 21100 8566 21128 8910
rect 20996 8560 21048 8566
rect 20996 8502 21048 8508
rect 21088 8560 21140 8566
rect 21088 8502 21140 8508
rect 21192 8430 21220 9454
rect 21284 9042 21312 9590
rect 21272 9036 21324 9042
rect 21272 8978 21324 8984
rect 21376 8838 21404 9998
rect 21468 8974 21496 10424
rect 21560 9654 21588 12192
rect 21548 9648 21600 9654
rect 21548 9590 21600 9596
rect 21652 9382 21680 12406
rect 21744 11150 21772 14962
rect 22008 14952 22060 14958
rect 22008 14894 22060 14900
rect 21824 14612 21876 14618
rect 21824 14554 21876 14560
rect 21836 14074 21864 14554
rect 22020 14414 22048 14894
rect 22008 14408 22060 14414
rect 22008 14350 22060 14356
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 22112 13802 22140 15438
rect 22204 14618 22232 17614
rect 22388 17320 22416 17614
rect 23673 17436 23981 17445
rect 23673 17434 23679 17436
rect 23735 17434 23759 17436
rect 23815 17434 23839 17436
rect 23895 17434 23919 17436
rect 23975 17434 23981 17436
rect 23735 17382 23737 17434
rect 23917 17382 23919 17434
rect 23673 17380 23679 17382
rect 23735 17380 23759 17382
rect 23815 17380 23839 17382
rect 23895 17380 23919 17382
rect 23975 17380 23981 17382
rect 23673 17371 23981 17380
rect 22296 17292 22416 17320
rect 22296 17134 22324 17292
rect 22376 17196 22428 17202
rect 22376 17138 22428 17144
rect 22284 17128 22336 17134
rect 22284 17070 22336 17076
rect 22296 16794 22324 17070
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22388 16250 22416 17138
rect 23673 16348 23981 16357
rect 23673 16346 23679 16348
rect 23735 16346 23759 16348
rect 23815 16346 23839 16348
rect 23895 16346 23919 16348
rect 23975 16346 23981 16348
rect 23735 16294 23737 16346
rect 23917 16294 23919 16346
rect 23673 16292 23679 16294
rect 23735 16292 23759 16294
rect 23815 16292 23839 16294
rect 23895 16292 23919 16294
rect 23975 16292 23981 16294
rect 23673 16283 23981 16292
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 22388 15910 22416 16186
rect 22928 16108 22980 16114
rect 22928 16050 22980 16056
rect 22376 15904 22428 15910
rect 22376 15846 22428 15852
rect 22652 15564 22704 15570
rect 22652 15506 22704 15512
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 22192 14612 22244 14618
rect 22192 14554 22244 14560
rect 22296 14414 22324 15438
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22100 13796 22152 13802
rect 22100 13738 22152 13744
rect 21916 13728 21968 13734
rect 22192 13728 22244 13734
rect 21968 13688 22048 13716
rect 21916 13670 21968 13676
rect 21824 13388 21876 13394
rect 21824 13330 21876 13336
rect 21836 12918 21864 13330
rect 21824 12912 21876 12918
rect 21824 12854 21876 12860
rect 21836 12442 21864 12854
rect 21824 12436 21876 12442
rect 22020 12434 22048 13688
rect 22192 13670 22244 13676
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 21824 12378 21876 12384
rect 21928 12406 22048 12434
rect 21928 12306 21956 12406
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 21928 11218 21956 12242
rect 22008 12164 22060 12170
rect 22008 12106 22060 12112
rect 22020 11898 22048 12106
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 21916 11212 21968 11218
rect 21916 11154 21968 11160
rect 22112 11150 22140 12786
rect 21732 11144 21784 11150
rect 21732 11086 21784 11092
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 21744 10470 21772 11086
rect 22112 10606 22140 11086
rect 22100 10600 22152 10606
rect 22100 10542 22152 10548
rect 21732 10464 21784 10470
rect 21784 10424 21864 10452
rect 21732 10406 21784 10412
rect 21732 9580 21784 9586
rect 21732 9522 21784 9528
rect 21640 9376 21692 9382
rect 21640 9318 21692 9324
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21364 8832 21416 8838
rect 21364 8774 21416 8780
rect 20732 8350 20852 8378
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 20732 7886 20760 8350
rect 20833 8188 21141 8197
rect 20833 8186 20839 8188
rect 20895 8186 20919 8188
rect 20975 8186 20999 8188
rect 21055 8186 21079 8188
rect 21135 8186 21141 8188
rect 20895 8134 20897 8186
rect 21077 8134 21079 8186
rect 20833 8132 20839 8134
rect 20895 8132 20919 8134
rect 20975 8132 20999 8134
rect 21055 8132 21079 8134
rect 21135 8132 21141 8134
rect 20833 8123 21141 8132
rect 21192 7886 21220 8366
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 20833 7100 21141 7109
rect 20833 7098 20839 7100
rect 20895 7098 20919 7100
rect 20975 7098 20999 7100
rect 21055 7098 21079 7100
rect 21135 7098 21141 7100
rect 20895 7046 20897 7098
rect 21077 7046 21079 7098
rect 20833 7044 20839 7046
rect 20895 7044 20919 7046
rect 20975 7044 20999 7046
rect 21055 7044 21079 7046
rect 21135 7044 21141 7046
rect 20833 7035 21141 7044
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20444 6384 20496 6390
rect 20444 6326 20496 6332
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 20272 4826 20300 5170
rect 20444 5160 20496 5166
rect 20548 5148 20576 6598
rect 20640 5778 20668 6734
rect 21284 6322 21312 6734
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 20833 6012 21141 6021
rect 20833 6010 20839 6012
rect 20895 6010 20919 6012
rect 20975 6010 20999 6012
rect 21055 6010 21079 6012
rect 21135 6010 21141 6012
rect 20895 5958 20897 6010
rect 21077 5958 21079 6010
rect 20833 5956 20839 5958
rect 20895 5956 20919 5958
rect 20975 5956 20999 5958
rect 21055 5956 21079 5958
rect 21135 5956 21141 5958
rect 20833 5947 21141 5956
rect 21272 5908 21324 5914
rect 21272 5850 21324 5856
rect 20628 5772 20680 5778
rect 20628 5714 20680 5720
rect 21178 5672 21234 5681
rect 20628 5636 20680 5642
rect 21178 5607 21234 5616
rect 20628 5578 20680 5584
rect 20640 5234 20668 5578
rect 21192 5370 21220 5607
rect 21180 5364 21232 5370
rect 21180 5306 21232 5312
rect 21284 5234 21312 5850
rect 20628 5228 20680 5234
rect 20628 5170 20680 5176
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 20496 5120 20576 5148
rect 20444 5102 20496 5108
rect 20640 4826 20668 5170
rect 20833 4924 21141 4933
rect 20833 4922 20839 4924
rect 20895 4922 20919 4924
rect 20975 4922 20999 4924
rect 21055 4922 21079 4924
rect 21135 4922 21141 4924
rect 20895 4870 20897 4922
rect 21077 4870 21079 4922
rect 20833 4868 20839 4870
rect 20895 4868 20919 4870
rect 20975 4868 20999 4870
rect 21055 4868 21079 4870
rect 21135 4868 21141 4870
rect 20833 4859 21141 4868
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20628 4820 20680 4826
rect 20628 4762 20680 4768
rect 21468 4690 21496 8910
rect 21640 8832 21692 8838
rect 21640 8774 21692 8780
rect 21548 8492 21600 8498
rect 21548 8434 21600 8440
rect 21560 6798 21588 8434
rect 21548 6792 21600 6798
rect 21548 6734 21600 6740
rect 21652 6730 21680 8774
rect 21744 7546 21772 9522
rect 21836 9042 21864 10424
rect 22112 9722 22140 10542
rect 22100 9716 22152 9722
rect 22100 9658 22152 9664
rect 22020 9586 22140 9602
rect 22008 9580 22140 9586
rect 22060 9574 22140 9580
rect 22008 9522 22060 9528
rect 22112 9382 22140 9574
rect 22100 9376 22152 9382
rect 22100 9318 22152 9324
rect 22204 9178 22232 13670
rect 22296 11218 22324 14350
rect 22376 13728 22428 13734
rect 22376 13670 22428 13676
rect 22388 12102 22416 13670
rect 22480 12850 22508 15302
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22480 12374 22508 12786
rect 22468 12368 22520 12374
rect 22468 12310 22520 12316
rect 22480 12170 22508 12310
rect 22468 12164 22520 12170
rect 22468 12106 22520 12112
rect 22376 12096 22428 12102
rect 22376 12038 22428 12044
rect 22572 11830 22600 15098
rect 22664 12434 22692 15506
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22756 13433 22784 13670
rect 22742 13424 22798 13433
rect 22742 13359 22798 13368
rect 22848 13326 22876 14214
rect 22940 13530 22968 16050
rect 23673 15260 23981 15269
rect 23673 15258 23679 15260
rect 23735 15258 23759 15260
rect 23815 15258 23839 15260
rect 23895 15258 23919 15260
rect 23975 15258 23981 15260
rect 23735 15206 23737 15258
rect 23917 15206 23919 15258
rect 23673 15204 23679 15206
rect 23735 15204 23759 15206
rect 23815 15204 23839 15206
rect 23895 15204 23919 15206
rect 23975 15204 23981 15206
rect 23673 15195 23981 15204
rect 23204 14408 23256 14414
rect 23204 14350 23256 14356
rect 22928 13524 22980 13530
rect 22928 13466 22980 13472
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22928 12640 22980 12646
rect 22928 12582 22980 12588
rect 22664 12406 22876 12434
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22652 12164 22704 12170
rect 22652 12106 22704 12112
rect 22560 11824 22612 11830
rect 22560 11766 22612 11772
rect 22376 11280 22428 11286
rect 22376 11222 22428 11228
rect 22284 11212 22336 11218
rect 22284 11154 22336 11160
rect 22296 9926 22324 11154
rect 22388 10538 22416 11222
rect 22664 11150 22692 12106
rect 22756 11830 22784 12174
rect 22744 11824 22796 11830
rect 22744 11766 22796 11772
rect 22468 11144 22520 11150
rect 22468 11086 22520 11092
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 22376 10532 22428 10538
rect 22376 10474 22428 10480
rect 22480 10266 22508 11086
rect 22560 10464 22612 10470
rect 22560 10406 22612 10412
rect 22468 10260 22520 10266
rect 22468 10202 22520 10208
rect 22284 9920 22336 9926
rect 22284 9862 22336 9868
rect 22296 9568 22324 9862
rect 22296 9540 22416 9568
rect 22284 9444 22336 9450
rect 22284 9386 22336 9392
rect 22192 9172 22244 9178
rect 22192 9114 22244 9120
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 22296 8498 22324 9386
rect 22388 9382 22416 9540
rect 22376 9376 22428 9382
rect 22376 9318 22428 9324
rect 22468 8968 22520 8974
rect 22468 8910 22520 8916
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 22376 8424 22428 8430
rect 22006 8392 22062 8401
rect 22376 8366 22428 8372
rect 22006 8327 22062 8336
rect 21732 7540 21784 7546
rect 21732 7482 21784 7488
rect 21640 6724 21692 6730
rect 21640 6666 21692 6672
rect 22020 6322 22048 8327
rect 22284 8016 22336 8022
rect 22284 7958 22336 7964
rect 22190 6896 22246 6905
rect 22190 6831 22192 6840
rect 22244 6831 22246 6840
rect 22192 6802 22244 6808
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 22008 6316 22060 6322
rect 22008 6258 22060 6264
rect 22112 5710 22140 6598
rect 22296 5778 22324 7958
rect 22388 6458 22416 8366
rect 22480 7274 22508 8910
rect 22572 8498 22600 10406
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 22560 7744 22612 7750
rect 22560 7686 22612 7692
rect 22468 7268 22520 7274
rect 22468 7210 22520 7216
rect 22376 6452 22428 6458
rect 22376 6394 22428 6400
rect 22480 6390 22508 7210
rect 22468 6384 22520 6390
rect 22468 6326 22520 6332
rect 22480 5914 22508 6326
rect 22468 5908 22520 5914
rect 22468 5850 22520 5856
rect 22284 5772 22336 5778
rect 22284 5714 22336 5720
rect 22100 5704 22152 5710
rect 22100 5646 22152 5652
rect 22112 5302 22140 5646
rect 22100 5296 22152 5302
rect 22100 5238 22152 5244
rect 21456 4684 21508 4690
rect 21456 4626 21508 4632
rect 22296 4622 22324 5714
rect 22572 5710 22600 7686
rect 22664 6866 22692 9318
rect 22756 9110 22784 11766
rect 22848 9178 22876 12406
rect 22940 12306 22968 12582
rect 22928 12300 22980 12306
rect 22928 12242 22980 12248
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22744 9104 22796 9110
rect 22744 9046 22796 9052
rect 22756 8090 22784 9046
rect 22836 8900 22888 8906
rect 22836 8842 22888 8848
rect 22744 8084 22796 8090
rect 22744 8026 22796 8032
rect 22756 7546 22784 8026
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22848 7410 22876 8842
rect 22836 7404 22888 7410
rect 22836 7346 22888 7352
rect 22744 7200 22796 7206
rect 22744 7142 22796 7148
rect 22652 6860 22704 6866
rect 22652 6802 22704 6808
rect 22756 6798 22784 7142
rect 22744 6792 22796 6798
rect 22744 6734 22796 6740
rect 22848 6118 22876 7346
rect 22652 6112 22704 6118
rect 22652 6054 22704 6060
rect 22836 6112 22888 6118
rect 22836 6054 22888 6060
rect 22560 5704 22612 5710
rect 22560 5646 22612 5652
rect 22284 4616 22336 4622
rect 22284 4558 22336 4564
rect 22664 4282 22692 6054
rect 22940 5778 22968 12242
rect 23216 12238 23244 14350
rect 23673 14172 23981 14181
rect 23673 14170 23679 14172
rect 23735 14170 23759 14172
rect 23815 14170 23839 14172
rect 23895 14170 23919 14172
rect 23975 14170 23981 14172
rect 23735 14118 23737 14170
rect 23917 14118 23919 14170
rect 23673 14116 23679 14118
rect 23735 14116 23759 14118
rect 23815 14116 23839 14118
rect 23895 14116 23919 14118
rect 23975 14116 23981 14118
rect 23673 14107 23981 14116
rect 23673 13084 23981 13093
rect 23673 13082 23679 13084
rect 23735 13082 23759 13084
rect 23815 13082 23839 13084
rect 23895 13082 23919 13084
rect 23975 13082 23981 13084
rect 23735 13030 23737 13082
rect 23917 13030 23919 13082
rect 23673 13028 23679 13030
rect 23735 13028 23759 13030
rect 23815 13028 23839 13030
rect 23895 13028 23919 13030
rect 23975 13028 23981 13030
rect 23673 13019 23981 13028
rect 23020 12232 23072 12238
rect 23020 12174 23072 12180
rect 23204 12232 23256 12238
rect 23204 12174 23256 12180
rect 23032 11694 23060 12174
rect 23020 11688 23072 11694
rect 23020 11630 23072 11636
rect 23216 11286 23244 12174
rect 23673 11996 23981 12005
rect 23673 11994 23679 11996
rect 23735 11994 23759 11996
rect 23815 11994 23839 11996
rect 23895 11994 23919 11996
rect 23975 11994 23981 11996
rect 23735 11942 23737 11994
rect 23917 11942 23919 11994
rect 23673 11940 23679 11942
rect 23735 11940 23759 11942
rect 23815 11940 23839 11942
rect 23895 11940 23919 11942
rect 23975 11940 23981 11942
rect 23673 11931 23981 11940
rect 23204 11280 23256 11286
rect 23204 11222 23256 11228
rect 23216 8974 23244 11222
rect 23673 10908 23981 10917
rect 23673 10906 23679 10908
rect 23735 10906 23759 10908
rect 23815 10906 23839 10908
rect 23895 10906 23919 10908
rect 23975 10906 23981 10908
rect 23735 10854 23737 10906
rect 23917 10854 23919 10906
rect 23673 10852 23679 10854
rect 23735 10852 23759 10854
rect 23815 10852 23839 10854
rect 23895 10852 23919 10854
rect 23975 10852 23981 10854
rect 23673 10843 23981 10852
rect 23673 9820 23981 9829
rect 23673 9818 23679 9820
rect 23735 9818 23759 9820
rect 23815 9818 23839 9820
rect 23895 9818 23919 9820
rect 23975 9818 23981 9820
rect 23735 9766 23737 9818
rect 23917 9766 23919 9818
rect 23673 9764 23679 9766
rect 23735 9764 23759 9766
rect 23815 9764 23839 9766
rect 23895 9764 23919 9766
rect 23975 9764 23981 9766
rect 23673 9755 23981 9764
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 23020 8492 23072 8498
rect 23020 8434 23072 8440
rect 23032 6458 23060 8434
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 23216 6322 23244 8910
rect 23673 8732 23981 8741
rect 23673 8730 23679 8732
rect 23735 8730 23759 8732
rect 23815 8730 23839 8732
rect 23895 8730 23919 8732
rect 23975 8730 23981 8732
rect 23735 8678 23737 8730
rect 23917 8678 23919 8730
rect 23673 8676 23679 8678
rect 23735 8676 23759 8678
rect 23815 8676 23839 8678
rect 23895 8676 23919 8678
rect 23975 8676 23981 8678
rect 23673 8667 23981 8676
rect 23673 7644 23981 7653
rect 23673 7642 23679 7644
rect 23735 7642 23759 7644
rect 23815 7642 23839 7644
rect 23895 7642 23919 7644
rect 23975 7642 23981 7644
rect 23735 7590 23737 7642
rect 23917 7590 23919 7642
rect 23673 7588 23679 7590
rect 23735 7588 23759 7590
rect 23815 7588 23839 7590
rect 23895 7588 23919 7590
rect 23975 7588 23981 7590
rect 23673 7579 23981 7588
rect 23673 6556 23981 6565
rect 23673 6554 23679 6556
rect 23735 6554 23759 6556
rect 23815 6554 23839 6556
rect 23895 6554 23919 6556
rect 23975 6554 23981 6556
rect 23735 6502 23737 6554
rect 23917 6502 23919 6554
rect 23673 6500 23679 6502
rect 23735 6500 23759 6502
rect 23815 6500 23839 6502
rect 23895 6500 23919 6502
rect 23975 6500 23981 6502
rect 23673 6491 23981 6500
rect 23204 6316 23256 6322
rect 23204 6258 23256 6264
rect 23296 6248 23348 6254
rect 23296 6190 23348 6196
rect 22928 5772 22980 5778
rect 22928 5714 22980 5720
rect 22940 5386 22968 5714
rect 23308 5681 23336 6190
rect 23294 5672 23350 5681
rect 23294 5607 23350 5616
rect 23673 5468 23981 5477
rect 23673 5466 23679 5468
rect 23735 5466 23759 5468
rect 23815 5466 23839 5468
rect 23895 5466 23919 5468
rect 23975 5466 23981 5468
rect 23735 5414 23737 5466
rect 23917 5414 23919 5466
rect 23673 5412 23679 5414
rect 23735 5412 23759 5414
rect 23815 5412 23839 5414
rect 23895 5412 23919 5414
rect 23975 5412 23981 5414
rect 23673 5403 23981 5412
rect 22848 5370 22968 5386
rect 22836 5364 22968 5370
rect 22888 5358 22968 5364
rect 22836 5306 22888 5312
rect 22848 5234 22876 5306
rect 22928 5296 22980 5302
rect 22928 5238 22980 5244
rect 22836 5228 22888 5234
rect 22836 5170 22888 5176
rect 22940 4622 22968 5238
rect 22744 4616 22796 4622
rect 22744 4558 22796 4564
rect 22928 4616 22980 4622
rect 22928 4558 22980 4564
rect 22652 4276 22704 4282
rect 22652 4218 22704 4224
rect 22756 4146 22784 4558
rect 22940 4214 22968 4558
rect 23673 4380 23981 4389
rect 23673 4378 23679 4380
rect 23735 4378 23759 4380
rect 23815 4378 23839 4380
rect 23895 4378 23919 4380
rect 23975 4378 23981 4380
rect 23735 4326 23737 4378
rect 23917 4326 23919 4378
rect 23673 4324 23679 4326
rect 23735 4324 23759 4326
rect 23815 4324 23839 4326
rect 23895 4324 23919 4326
rect 23975 4324 23981 4326
rect 23673 4315 23981 4324
rect 22928 4208 22980 4214
rect 22928 4150 22980 4156
rect 22744 4140 22796 4146
rect 22744 4082 22796 4088
rect 20833 3836 21141 3845
rect 20833 3834 20839 3836
rect 20895 3834 20919 3836
rect 20975 3834 20999 3836
rect 21055 3834 21079 3836
rect 21135 3834 21141 3836
rect 20895 3782 20897 3834
rect 21077 3782 21079 3834
rect 20833 3780 20839 3782
rect 20895 3780 20919 3782
rect 20975 3780 20999 3782
rect 21055 3780 21079 3782
rect 21135 3780 21141 3782
rect 20833 3771 21141 3780
rect 20076 3596 20128 3602
rect 20076 3538 20128 3544
rect 23388 3596 23440 3602
rect 23388 3538 23440 3544
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 19996 3194 20024 3334
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 20640 3126 20668 3334
rect 20628 3120 20680 3126
rect 20628 3062 20680 3068
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 19248 3052 19300 3058
rect 19248 2994 19300 3000
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 17868 2984 17920 2990
rect 17868 2926 17920 2932
rect 19524 2916 19576 2922
rect 19524 2858 19576 2864
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17420 2446 17448 2790
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 16764 2372 16816 2378
rect 16764 2314 16816 2320
rect 17992 2204 18300 2213
rect 17992 2202 17998 2204
rect 18054 2202 18078 2204
rect 18134 2202 18158 2204
rect 18214 2202 18238 2204
rect 18294 2202 18300 2204
rect 18054 2150 18056 2202
rect 18236 2150 18238 2202
rect 17992 2148 17998 2150
rect 18054 2148 18078 2150
rect 18134 2148 18158 2150
rect 18214 2148 18238 2150
rect 18294 2148 18300 2150
rect 17992 2139 18300 2148
rect 18524 1086 18552 2382
rect 16948 1080 17000 1086
rect 16948 1022 17000 1028
rect 18512 1080 18564 1086
rect 18512 1022 18564 1028
rect 18880 1080 18932 1086
rect 18880 1022 18932 1028
rect 16316 870 16620 898
rect 16316 800 16344 870
rect 16960 800 16988 1022
rect 18236 1012 18288 1018
rect 18236 954 18288 960
rect 17592 944 17644 950
rect 17592 886 17644 892
rect 17604 800 17632 886
rect 18248 800 18276 954
rect 18892 800 18920 1022
rect 19444 950 19472 2382
rect 19432 944 19484 950
rect 19432 886 19484 892
rect 19536 800 19564 2858
rect 21456 2848 21508 2854
rect 21456 2790 21508 2796
rect 22100 2848 22152 2854
rect 22100 2790 22152 2796
rect 20833 2748 21141 2757
rect 20833 2746 20839 2748
rect 20895 2746 20919 2748
rect 20975 2746 20999 2748
rect 21055 2746 21079 2748
rect 21135 2746 21141 2748
rect 20895 2694 20897 2746
rect 21077 2694 21079 2746
rect 20833 2692 20839 2694
rect 20895 2692 20919 2694
rect 20975 2692 20999 2694
rect 21055 2692 21079 2694
rect 21135 2692 21141 2694
rect 20833 2683 21141 2692
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 20088 1018 20116 2382
rect 20732 1086 20760 2382
rect 20720 1080 20772 1086
rect 20720 1022 20772 1028
rect 20076 1012 20128 1018
rect 20076 954 20128 960
rect 20812 1012 20864 1018
rect 20812 954 20864 960
rect 20168 944 20220 950
rect 20168 886 20220 892
rect 20180 800 20208 886
rect 20824 800 20852 954
rect 21468 800 21496 2790
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 22020 950 22048 2382
rect 22008 944 22060 950
rect 22008 886 22060 892
rect 22112 800 22140 2790
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 22664 1018 22692 2382
rect 22652 1012 22704 1018
rect 22652 954 22704 960
rect 22756 800 22784 3470
rect 23400 800 23428 3538
rect 23673 3292 23981 3301
rect 23673 3290 23679 3292
rect 23735 3290 23759 3292
rect 23815 3290 23839 3292
rect 23895 3290 23919 3292
rect 23975 3290 23981 3292
rect 23735 3238 23737 3290
rect 23917 3238 23919 3290
rect 23673 3236 23679 3238
rect 23735 3236 23759 3238
rect 23815 3236 23839 3238
rect 23895 3236 23919 3238
rect 23975 3236 23981 3238
rect 23673 3227 23981 3236
rect 23673 2204 23981 2213
rect 23673 2202 23679 2204
rect 23735 2202 23759 2204
rect 23815 2202 23839 2204
rect 23895 2202 23919 2204
rect 23975 2202 23981 2204
rect 23735 2150 23737 2202
rect 23917 2150 23919 2202
rect 23673 2148 23679 2150
rect 23735 2148 23759 2150
rect 23815 2148 23839 2150
rect 23895 2148 23919 2150
rect 23975 2148 23981 2150
rect 23673 2139 23981 2148
rect 12544 734 12756 762
rect 13082 0 13138 800
rect 13726 0 13782 800
rect 14370 0 14426 800
rect 15014 0 15070 800
rect 15658 0 15714 800
rect 16302 0 16358 800
rect 16946 0 17002 800
rect 17590 0 17646 800
rect 18234 0 18290 800
rect 18878 0 18934 800
rect 19522 0 19578 800
rect 20166 0 20222 800
rect 20810 0 20866 800
rect 21454 0 21510 800
rect 22098 0 22154 800
rect 22742 0 22798 800
rect 23386 0 23442 800
<< via2 >>
rect 3796 22330 3852 22332
rect 3876 22330 3932 22332
rect 3956 22330 4012 22332
rect 4036 22330 4092 22332
rect 3796 22278 3842 22330
rect 3842 22278 3852 22330
rect 3876 22278 3906 22330
rect 3906 22278 3918 22330
rect 3918 22278 3932 22330
rect 3956 22278 3970 22330
rect 3970 22278 3982 22330
rect 3982 22278 4012 22330
rect 4036 22278 4046 22330
rect 4046 22278 4092 22330
rect 3796 22276 3852 22278
rect 3876 22276 3932 22278
rect 3956 22276 4012 22278
rect 4036 22276 4092 22278
rect 1674 9560 1730 9616
rect 1490 9424 1546 9480
rect 9477 22330 9533 22332
rect 9557 22330 9613 22332
rect 9637 22330 9693 22332
rect 9717 22330 9773 22332
rect 9477 22278 9523 22330
rect 9523 22278 9533 22330
rect 9557 22278 9587 22330
rect 9587 22278 9599 22330
rect 9599 22278 9613 22330
rect 9637 22278 9651 22330
rect 9651 22278 9663 22330
rect 9663 22278 9693 22330
rect 9717 22278 9727 22330
rect 9727 22278 9773 22330
rect 9477 22276 9533 22278
rect 9557 22276 9613 22278
rect 9637 22276 9693 22278
rect 9717 22276 9773 22278
rect 15158 22330 15214 22332
rect 15238 22330 15294 22332
rect 15318 22330 15374 22332
rect 15398 22330 15454 22332
rect 15158 22278 15204 22330
rect 15204 22278 15214 22330
rect 15238 22278 15268 22330
rect 15268 22278 15280 22330
rect 15280 22278 15294 22330
rect 15318 22278 15332 22330
rect 15332 22278 15344 22330
rect 15344 22278 15374 22330
rect 15398 22278 15408 22330
rect 15408 22278 15454 22330
rect 15158 22276 15214 22278
rect 15238 22276 15294 22278
rect 15318 22276 15374 22278
rect 15398 22276 15454 22278
rect 2962 10668 3018 10704
rect 2962 10648 2964 10668
rect 2964 10648 3016 10668
rect 3016 10648 3018 10668
rect 3054 5652 3056 5672
rect 3056 5652 3108 5672
rect 3108 5652 3110 5672
rect 3054 5616 3110 5652
rect 6636 21786 6692 21788
rect 6716 21786 6772 21788
rect 6796 21786 6852 21788
rect 6876 21786 6932 21788
rect 6636 21734 6682 21786
rect 6682 21734 6692 21786
rect 6716 21734 6746 21786
rect 6746 21734 6758 21786
rect 6758 21734 6772 21786
rect 6796 21734 6810 21786
rect 6810 21734 6822 21786
rect 6822 21734 6852 21786
rect 6876 21734 6886 21786
rect 6886 21734 6932 21786
rect 6636 21732 6692 21734
rect 6716 21732 6772 21734
rect 6796 21732 6852 21734
rect 6876 21732 6932 21734
rect 3796 21242 3852 21244
rect 3876 21242 3932 21244
rect 3956 21242 4012 21244
rect 4036 21242 4092 21244
rect 3796 21190 3842 21242
rect 3842 21190 3852 21242
rect 3876 21190 3906 21242
rect 3906 21190 3918 21242
rect 3918 21190 3932 21242
rect 3956 21190 3970 21242
rect 3970 21190 3982 21242
rect 3982 21190 4012 21242
rect 4036 21190 4046 21242
rect 4046 21190 4092 21242
rect 3796 21188 3852 21190
rect 3876 21188 3932 21190
rect 3956 21188 4012 21190
rect 4036 21188 4092 21190
rect 3796 20154 3852 20156
rect 3876 20154 3932 20156
rect 3956 20154 4012 20156
rect 4036 20154 4092 20156
rect 3796 20102 3842 20154
rect 3842 20102 3852 20154
rect 3876 20102 3906 20154
rect 3906 20102 3918 20154
rect 3918 20102 3932 20154
rect 3956 20102 3970 20154
rect 3970 20102 3982 20154
rect 3982 20102 4012 20154
rect 4036 20102 4046 20154
rect 4046 20102 4092 20154
rect 3796 20100 3852 20102
rect 3876 20100 3932 20102
rect 3956 20100 4012 20102
rect 4036 20100 4092 20102
rect 3796 19066 3852 19068
rect 3876 19066 3932 19068
rect 3956 19066 4012 19068
rect 4036 19066 4092 19068
rect 3796 19014 3842 19066
rect 3842 19014 3852 19066
rect 3876 19014 3906 19066
rect 3906 19014 3918 19066
rect 3918 19014 3932 19066
rect 3956 19014 3970 19066
rect 3970 19014 3982 19066
rect 3982 19014 4012 19066
rect 4036 19014 4046 19066
rect 4046 19014 4092 19066
rect 3796 19012 3852 19014
rect 3876 19012 3932 19014
rect 3956 19012 4012 19014
rect 4036 19012 4092 19014
rect 3796 17978 3852 17980
rect 3876 17978 3932 17980
rect 3956 17978 4012 17980
rect 4036 17978 4092 17980
rect 3796 17926 3842 17978
rect 3842 17926 3852 17978
rect 3876 17926 3906 17978
rect 3906 17926 3918 17978
rect 3918 17926 3932 17978
rect 3956 17926 3970 17978
rect 3970 17926 3982 17978
rect 3982 17926 4012 17978
rect 4036 17926 4046 17978
rect 4046 17926 4092 17978
rect 3796 17924 3852 17926
rect 3876 17924 3932 17926
rect 3956 17924 4012 17926
rect 4036 17924 4092 17926
rect 3796 16890 3852 16892
rect 3876 16890 3932 16892
rect 3956 16890 4012 16892
rect 4036 16890 4092 16892
rect 3796 16838 3842 16890
rect 3842 16838 3852 16890
rect 3876 16838 3906 16890
rect 3906 16838 3918 16890
rect 3918 16838 3932 16890
rect 3956 16838 3970 16890
rect 3970 16838 3982 16890
rect 3982 16838 4012 16890
rect 4036 16838 4046 16890
rect 4046 16838 4092 16890
rect 3796 16836 3852 16838
rect 3876 16836 3932 16838
rect 3956 16836 4012 16838
rect 4036 16836 4092 16838
rect 3796 15802 3852 15804
rect 3876 15802 3932 15804
rect 3956 15802 4012 15804
rect 4036 15802 4092 15804
rect 3796 15750 3842 15802
rect 3842 15750 3852 15802
rect 3876 15750 3906 15802
rect 3906 15750 3918 15802
rect 3918 15750 3932 15802
rect 3956 15750 3970 15802
rect 3970 15750 3982 15802
rect 3982 15750 4012 15802
rect 4036 15750 4046 15802
rect 4046 15750 4092 15802
rect 3796 15748 3852 15750
rect 3876 15748 3932 15750
rect 3956 15748 4012 15750
rect 4036 15748 4092 15750
rect 3796 14714 3852 14716
rect 3876 14714 3932 14716
rect 3956 14714 4012 14716
rect 4036 14714 4092 14716
rect 3796 14662 3842 14714
rect 3842 14662 3852 14714
rect 3876 14662 3906 14714
rect 3906 14662 3918 14714
rect 3918 14662 3932 14714
rect 3956 14662 3970 14714
rect 3970 14662 3982 14714
rect 3982 14662 4012 14714
rect 4036 14662 4046 14714
rect 4046 14662 4092 14714
rect 3796 14660 3852 14662
rect 3876 14660 3932 14662
rect 3956 14660 4012 14662
rect 4036 14660 4092 14662
rect 3796 13626 3852 13628
rect 3876 13626 3932 13628
rect 3956 13626 4012 13628
rect 4036 13626 4092 13628
rect 3796 13574 3842 13626
rect 3842 13574 3852 13626
rect 3876 13574 3906 13626
rect 3906 13574 3918 13626
rect 3918 13574 3932 13626
rect 3956 13574 3970 13626
rect 3970 13574 3982 13626
rect 3982 13574 4012 13626
rect 4036 13574 4046 13626
rect 4046 13574 4092 13626
rect 3796 13572 3852 13574
rect 3876 13572 3932 13574
rect 3956 13572 4012 13574
rect 4036 13572 4092 13574
rect 3796 12538 3852 12540
rect 3876 12538 3932 12540
rect 3956 12538 4012 12540
rect 4036 12538 4092 12540
rect 3796 12486 3842 12538
rect 3842 12486 3852 12538
rect 3876 12486 3906 12538
rect 3906 12486 3918 12538
rect 3918 12486 3932 12538
rect 3956 12486 3970 12538
rect 3970 12486 3982 12538
rect 3982 12486 4012 12538
rect 4036 12486 4046 12538
rect 4046 12486 4092 12538
rect 3796 12484 3852 12486
rect 3876 12484 3932 12486
rect 3956 12484 4012 12486
rect 4036 12484 4092 12486
rect 3796 11450 3852 11452
rect 3876 11450 3932 11452
rect 3956 11450 4012 11452
rect 4036 11450 4092 11452
rect 3796 11398 3842 11450
rect 3842 11398 3852 11450
rect 3876 11398 3906 11450
rect 3906 11398 3918 11450
rect 3918 11398 3932 11450
rect 3956 11398 3970 11450
rect 3970 11398 3982 11450
rect 3982 11398 4012 11450
rect 4036 11398 4046 11450
rect 4046 11398 4092 11450
rect 3796 11396 3852 11398
rect 3876 11396 3932 11398
rect 3956 11396 4012 11398
rect 4036 11396 4092 11398
rect 3796 10362 3852 10364
rect 3876 10362 3932 10364
rect 3956 10362 4012 10364
rect 4036 10362 4092 10364
rect 3796 10310 3842 10362
rect 3842 10310 3852 10362
rect 3876 10310 3906 10362
rect 3906 10310 3918 10362
rect 3918 10310 3932 10362
rect 3956 10310 3970 10362
rect 3970 10310 3982 10362
rect 3982 10310 4012 10362
rect 4036 10310 4046 10362
rect 4046 10310 4092 10362
rect 3796 10308 3852 10310
rect 3876 10308 3932 10310
rect 3956 10308 4012 10310
rect 4036 10308 4092 10310
rect 4618 20712 4674 20768
rect 5354 19352 5410 19408
rect 4894 13268 4896 13288
rect 4896 13268 4948 13288
rect 4948 13268 4950 13288
rect 4894 13232 4950 13268
rect 3796 9274 3852 9276
rect 3876 9274 3932 9276
rect 3956 9274 4012 9276
rect 4036 9274 4092 9276
rect 3796 9222 3842 9274
rect 3842 9222 3852 9274
rect 3876 9222 3906 9274
rect 3906 9222 3918 9274
rect 3918 9222 3932 9274
rect 3956 9222 3970 9274
rect 3970 9222 3982 9274
rect 3982 9222 4012 9274
rect 4036 9222 4046 9274
rect 4046 9222 4092 9274
rect 3796 9220 3852 9222
rect 3876 9220 3932 9222
rect 3956 9220 4012 9222
rect 4036 9220 4092 9222
rect 3606 5636 3662 5672
rect 3606 5616 3608 5636
rect 3608 5616 3660 5636
rect 3660 5616 3662 5636
rect 3796 8186 3852 8188
rect 3876 8186 3932 8188
rect 3956 8186 4012 8188
rect 4036 8186 4092 8188
rect 3796 8134 3842 8186
rect 3842 8134 3852 8186
rect 3876 8134 3906 8186
rect 3906 8134 3918 8186
rect 3918 8134 3932 8186
rect 3956 8134 3970 8186
rect 3970 8134 3982 8186
rect 3982 8134 4012 8186
rect 4036 8134 4046 8186
rect 4046 8134 4092 8186
rect 3796 8132 3852 8134
rect 3876 8132 3932 8134
rect 3956 8132 4012 8134
rect 4036 8132 4092 8134
rect 3796 7098 3852 7100
rect 3876 7098 3932 7100
rect 3956 7098 4012 7100
rect 4036 7098 4092 7100
rect 3796 7046 3842 7098
rect 3842 7046 3852 7098
rect 3876 7046 3906 7098
rect 3906 7046 3918 7098
rect 3918 7046 3932 7098
rect 3956 7046 3970 7098
rect 3970 7046 3982 7098
rect 3982 7046 4012 7098
rect 4036 7046 4046 7098
rect 4046 7046 4092 7098
rect 3796 7044 3852 7046
rect 3876 7044 3932 7046
rect 3956 7044 4012 7046
rect 4036 7044 4092 7046
rect 3796 6010 3852 6012
rect 3876 6010 3932 6012
rect 3956 6010 4012 6012
rect 4036 6010 4092 6012
rect 3796 5958 3842 6010
rect 3842 5958 3852 6010
rect 3876 5958 3906 6010
rect 3906 5958 3918 6010
rect 3918 5958 3932 6010
rect 3956 5958 3970 6010
rect 3970 5958 3982 6010
rect 3982 5958 4012 6010
rect 4036 5958 4046 6010
rect 4046 5958 4092 6010
rect 3796 5956 3852 5958
rect 3876 5956 3932 5958
rect 3956 5956 4012 5958
rect 4036 5956 4092 5958
rect 2962 2916 3018 2952
rect 2962 2896 2964 2916
rect 2964 2896 3016 2916
rect 3016 2896 3018 2916
rect 3796 4922 3852 4924
rect 3876 4922 3932 4924
rect 3956 4922 4012 4924
rect 4036 4922 4092 4924
rect 3796 4870 3842 4922
rect 3842 4870 3852 4922
rect 3876 4870 3906 4922
rect 3906 4870 3918 4922
rect 3918 4870 3932 4922
rect 3956 4870 3970 4922
rect 3970 4870 3982 4922
rect 3982 4870 4012 4922
rect 4036 4870 4046 4922
rect 4046 4870 4092 4922
rect 3796 4868 3852 4870
rect 3876 4868 3932 4870
rect 3956 4868 4012 4870
rect 4036 4868 4092 4870
rect 3796 3834 3852 3836
rect 3876 3834 3932 3836
rect 3956 3834 4012 3836
rect 4036 3834 4092 3836
rect 3796 3782 3842 3834
rect 3842 3782 3852 3834
rect 3876 3782 3906 3834
rect 3906 3782 3918 3834
rect 3918 3782 3932 3834
rect 3956 3782 3970 3834
rect 3970 3782 3982 3834
rect 3982 3782 4012 3834
rect 4036 3782 4046 3834
rect 4046 3782 4092 3834
rect 3796 3780 3852 3782
rect 3876 3780 3932 3782
rect 3956 3780 4012 3782
rect 4036 3780 4092 3782
rect 3422 2488 3478 2544
rect 3796 2746 3852 2748
rect 3876 2746 3932 2748
rect 3956 2746 4012 2748
rect 4036 2746 4092 2748
rect 3796 2694 3842 2746
rect 3842 2694 3852 2746
rect 3876 2694 3906 2746
rect 3906 2694 3918 2746
rect 3918 2694 3932 2746
rect 3956 2694 3970 2746
rect 3970 2694 3982 2746
rect 3982 2694 4012 2746
rect 4036 2694 4046 2746
rect 4046 2694 4092 2746
rect 3796 2692 3852 2694
rect 3876 2692 3932 2694
rect 3956 2692 4012 2694
rect 4036 2692 4092 2694
rect 4894 9560 4950 9616
rect 5446 12044 5448 12064
rect 5448 12044 5500 12064
rect 5500 12044 5502 12064
rect 5446 12008 5502 12044
rect 6636 20698 6692 20700
rect 6716 20698 6772 20700
rect 6796 20698 6852 20700
rect 6876 20698 6932 20700
rect 6636 20646 6682 20698
rect 6682 20646 6692 20698
rect 6716 20646 6746 20698
rect 6746 20646 6758 20698
rect 6758 20646 6772 20698
rect 6796 20646 6810 20698
rect 6810 20646 6822 20698
rect 6822 20646 6852 20698
rect 6876 20646 6886 20698
rect 6886 20646 6932 20698
rect 6636 20644 6692 20646
rect 6716 20644 6772 20646
rect 6796 20644 6852 20646
rect 6876 20644 6932 20646
rect 6090 16632 6146 16688
rect 5998 13232 6054 13288
rect 6636 19610 6692 19612
rect 6716 19610 6772 19612
rect 6796 19610 6852 19612
rect 6876 19610 6932 19612
rect 6636 19558 6682 19610
rect 6682 19558 6692 19610
rect 6716 19558 6746 19610
rect 6746 19558 6758 19610
rect 6758 19558 6772 19610
rect 6796 19558 6810 19610
rect 6810 19558 6822 19610
rect 6822 19558 6852 19610
rect 6876 19558 6886 19610
rect 6886 19558 6932 19610
rect 6636 19556 6692 19558
rect 6716 19556 6772 19558
rect 6796 19556 6852 19558
rect 6876 19556 6932 19558
rect 6636 18522 6692 18524
rect 6716 18522 6772 18524
rect 6796 18522 6852 18524
rect 6876 18522 6932 18524
rect 6636 18470 6682 18522
rect 6682 18470 6692 18522
rect 6716 18470 6746 18522
rect 6746 18470 6758 18522
rect 6758 18470 6772 18522
rect 6796 18470 6810 18522
rect 6810 18470 6822 18522
rect 6822 18470 6852 18522
rect 6876 18470 6886 18522
rect 6886 18470 6932 18522
rect 6636 18468 6692 18470
rect 6716 18468 6772 18470
rect 6796 18468 6852 18470
rect 6876 18468 6932 18470
rect 6636 17434 6692 17436
rect 6716 17434 6772 17436
rect 6796 17434 6852 17436
rect 6876 17434 6932 17436
rect 6636 17382 6682 17434
rect 6682 17382 6692 17434
rect 6716 17382 6746 17434
rect 6746 17382 6758 17434
rect 6758 17382 6772 17434
rect 6796 17382 6810 17434
rect 6810 17382 6822 17434
rect 6822 17382 6852 17434
rect 6876 17382 6886 17434
rect 6886 17382 6932 17434
rect 6636 17380 6692 17382
rect 6716 17380 6772 17382
rect 6796 17380 6852 17382
rect 6876 17380 6932 17382
rect 6636 16346 6692 16348
rect 6716 16346 6772 16348
rect 6796 16346 6852 16348
rect 6876 16346 6932 16348
rect 6636 16294 6682 16346
rect 6682 16294 6692 16346
rect 6716 16294 6746 16346
rect 6746 16294 6758 16346
rect 6758 16294 6772 16346
rect 6796 16294 6810 16346
rect 6810 16294 6822 16346
rect 6822 16294 6852 16346
rect 6876 16294 6886 16346
rect 6886 16294 6932 16346
rect 6636 16292 6692 16294
rect 6716 16292 6772 16294
rect 6796 16292 6852 16294
rect 6876 16292 6932 16294
rect 6636 15258 6692 15260
rect 6716 15258 6772 15260
rect 6796 15258 6852 15260
rect 6876 15258 6932 15260
rect 6636 15206 6682 15258
rect 6682 15206 6692 15258
rect 6716 15206 6746 15258
rect 6746 15206 6758 15258
rect 6758 15206 6772 15258
rect 6796 15206 6810 15258
rect 6810 15206 6822 15258
rect 6822 15206 6852 15258
rect 6876 15206 6886 15258
rect 6886 15206 6932 15258
rect 6636 15204 6692 15206
rect 6716 15204 6772 15206
rect 6796 15204 6852 15206
rect 6876 15204 6932 15206
rect 6636 14170 6692 14172
rect 6716 14170 6772 14172
rect 6796 14170 6852 14172
rect 6876 14170 6932 14172
rect 6636 14118 6682 14170
rect 6682 14118 6692 14170
rect 6716 14118 6746 14170
rect 6746 14118 6758 14170
rect 6758 14118 6772 14170
rect 6796 14118 6810 14170
rect 6810 14118 6822 14170
rect 6822 14118 6852 14170
rect 6876 14118 6886 14170
rect 6886 14118 6932 14170
rect 6636 14116 6692 14118
rect 6716 14116 6772 14118
rect 6796 14116 6852 14118
rect 6876 14116 6932 14118
rect 6636 13082 6692 13084
rect 6716 13082 6772 13084
rect 6796 13082 6852 13084
rect 6876 13082 6932 13084
rect 6636 13030 6682 13082
rect 6682 13030 6692 13082
rect 6716 13030 6746 13082
rect 6746 13030 6758 13082
rect 6758 13030 6772 13082
rect 6796 13030 6810 13082
rect 6810 13030 6822 13082
rect 6822 13030 6852 13082
rect 6876 13030 6886 13082
rect 6886 13030 6932 13082
rect 6636 13028 6692 13030
rect 6716 13028 6772 13030
rect 6796 13028 6852 13030
rect 6876 13028 6932 13030
rect 6636 11994 6692 11996
rect 6716 11994 6772 11996
rect 6796 11994 6852 11996
rect 6876 11994 6932 11996
rect 6636 11942 6682 11994
rect 6682 11942 6692 11994
rect 6716 11942 6746 11994
rect 6746 11942 6758 11994
rect 6758 11942 6772 11994
rect 6796 11942 6810 11994
rect 6810 11942 6822 11994
rect 6822 11942 6852 11994
rect 6876 11942 6886 11994
rect 6886 11942 6932 11994
rect 6636 11940 6692 11942
rect 6716 11940 6772 11942
rect 6796 11940 6852 11942
rect 6876 11940 6932 11942
rect 5722 9460 5724 9480
rect 5724 9460 5776 9480
rect 5776 9460 5778 9480
rect 5722 9424 5778 9460
rect 5446 3440 5502 3496
rect 5814 4936 5870 4992
rect 6636 10906 6692 10908
rect 6716 10906 6772 10908
rect 6796 10906 6852 10908
rect 6876 10906 6932 10908
rect 6636 10854 6682 10906
rect 6682 10854 6692 10906
rect 6716 10854 6746 10906
rect 6746 10854 6758 10906
rect 6758 10854 6772 10906
rect 6796 10854 6810 10906
rect 6810 10854 6822 10906
rect 6822 10854 6852 10906
rect 6876 10854 6886 10906
rect 6886 10854 6932 10906
rect 6636 10852 6692 10854
rect 6716 10852 6772 10854
rect 6796 10852 6852 10854
rect 6876 10852 6932 10854
rect 6636 9818 6692 9820
rect 6716 9818 6772 9820
rect 6796 9818 6852 9820
rect 6876 9818 6932 9820
rect 6636 9766 6682 9818
rect 6682 9766 6692 9818
rect 6716 9766 6746 9818
rect 6746 9766 6758 9818
rect 6758 9766 6772 9818
rect 6796 9766 6810 9818
rect 6810 9766 6822 9818
rect 6822 9766 6852 9818
rect 6876 9766 6886 9818
rect 6886 9766 6932 9818
rect 6636 9764 6692 9766
rect 6716 9764 6772 9766
rect 6796 9764 6852 9766
rect 6876 9764 6932 9766
rect 6550 9560 6606 9616
rect 6636 8730 6692 8732
rect 6716 8730 6772 8732
rect 6796 8730 6852 8732
rect 6876 8730 6932 8732
rect 6636 8678 6682 8730
rect 6682 8678 6692 8730
rect 6716 8678 6746 8730
rect 6746 8678 6758 8730
rect 6758 8678 6772 8730
rect 6796 8678 6810 8730
rect 6810 8678 6822 8730
rect 6822 8678 6852 8730
rect 6876 8678 6886 8730
rect 6886 8678 6932 8730
rect 6636 8676 6692 8678
rect 6716 8676 6772 8678
rect 6796 8676 6852 8678
rect 6876 8676 6932 8678
rect 6636 7642 6692 7644
rect 6716 7642 6772 7644
rect 6796 7642 6852 7644
rect 6876 7642 6932 7644
rect 6636 7590 6682 7642
rect 6682 7590 6692 7642
rect 6716 7590 6746 7642
rect 6746 7590 6758 7642
rect 6758 7590 6772 7642
rect 6796 7590 6810 7642
rect 6810 7590 6822 7642
rect 6822 7590 6852 7642
rect 6876 7590 6886 7642
rect 6886 7590 6932 7642
rect 6636 7588 6692 7590
rect 6716 7588 6772 7590
rect 6796 7588 6852 7590
rect 6876 7588 6932 7590
rect 6826 6724 6882 6760
rect 6826 6704 6828 6724
rect 6828 6704 6880 6724
rect 6880 6704 6882 6724
rect 6636 6554 6692 6556
rect 6716 6554 6772 6556
rect 6796 6554 6852 6556
rect 6876 6554 6932 6556
rect 6636 6502 6682 6554
rect 6682 6502 6692 6554
rect 6716 6502 6746 6554
rect 6746 6502 6758 6554
rect 6758 6502 6772 6554
rect 6796 6502 6810 6554
rect 6810 6502 6822 6554
rect 6822 6502 6852 6554
rect 6876 6502 6886 6554
rect 6886 6502 6932 6554
rect 6636 6500 6692 6502
rect 6716 6500 6772 6502
rect 6796 6500 6852 6502
rect 6876 6500 6932 6502
rect 6636 5466 6692 5468
rect 6716 5466 6772 5468
rect 6796 5466 6852 5468
rect 6876 5466 6932 5468
rect 6636 5414 6682 5466
rect 6682 5414 6692 5466
rect 6716 5414 6746 5466
rect 6746 5414 6758 5466
rect 6758 5414 6772 5466
rect 6796 5414 6810 5466
rect 6810 5414 6822 5466
rect 6822 5414 6852 5466
rect 6876 5414 6886 5466
rect 6886 5414 6932 5466
rect 6636 5412 6692 5414
rect 6716 5412 6772 5414
rect 6796 5412 6852 5414
rect 6876 5412 6932 5414
rect 6642 5072 6698 5128
rect 6636 4378 6692 4380
rect 6716 4378 6772 4380
rect 6796 4378 6852 4380
rect 6876 4378 6932 4380
rect 6636 4326 6682 4378
rect 6682 4326 6692 4378
rect 6716 4326 6746 4378
rect 6746 4326 6758 4378
rect 6758 4326 6772 4378
rect 6796 4326 6810 4378
rect 6810 4326 6822 4378
rect 6822 4326 6852 4378
rect 6876 4326 6886 4378
rect 6886 4326 6932 4378
rect 6636 4324 6692 4326
rect 6716 4324 6772 4326
rect 6796 4324 6852 4326
rect 6876 4324 6932 4326
rect 9477 21242 9533 21244
rect 9557 21242 9613 21244
rect 9637 21242 9693 21244
rect 9717 21242 9773 21244
rect 9477 21190 9523 21242
rect 9523 21190 9533 21242
rect 9557 21190 9587 21242
rect 9587 21190 9599 21242
rect 9599 21190 9613 21242
rect 9637 21190 9651 21242
rect 9651 21190 9663 21242
rect 9663 21190 9693 21242
rect 9717 21190 9727 21242
rect 9727 21190 9773 21242
rect 9477 21188 9533 21190
rect 9557 21188 9613 21190
rect 9637 21188 9693 21190
rect 9717 21188 9773 21190
rect 9477 20154 9533 20156
rect 9557 20154 9613 20156
rect 9637 20154 9693 20156
rect 9717 20154 9773 20156
rect 9477 20102 9523 20154
rect 9523 20102 9533 20154
rect 9557 20102 9587 20154
rect 9587 20102 9599 20154
rect 9599 20102 9613 20154
rect 9637 20102 9651 20154
rect 9651 20102 9663 20154
rect 9663 20102 9693 20154
rect 9717 20102 9727 20154
rect 9727 20102 9773 20154
rect 9477 20100 9533 20102
rect 9557 20100 9613 20102
rect 9637 20100 9693 20102
rect 9717 20100 9773 20102
rect 8482 10648 8538 10704
rect 7378 4936 7434 4992
rect 6550 3984 6606 4040
rect 7194 3576 7250 3632
rect 7102 3304 7158 3360
rect 6636 3290 6692 3292
rect 6716 3290 6772 3292
rect 6796 3290 6852 3292
rect 6876 3290 6932 3292
rect 6636 3238 6682 3290
rect 6682 3238 6692 3290
rect 6716 3238 6746 3290
rect 6746 3238 6758 3290
rect 6758 3238 6772 3290
rect 6796 3238 6810 3290
rect 6810 3238 6822 3290
rect 6822 3238 6852 3290
rect 6876 3238 6886 3290
rect 6886 3238 6932 3290
rect 6636 3236 6692 3238
rect 6716 3236 6772 3238
rect 6796 3236 6852 3238
rect 6876 3236 6932 3238
rect 9477 19066 9533 19068
rect 9557 19066 9613 19068
rect 9637 19066 9693 19068
rect 9717 19066 9773 19068
rect 9477 19014 9523 19066
rect 9523 19014 9533 19066
rect 9557 19014 9587 19066
rect 9587 19014 9599 19066
rect 9599 19014 9613 19066
rect 9637 19014 9651 19066
rect 9651 19014 9663 19066
rect 9663 19014 9693 19066
rect 9717 19014 9727 19066
rect 9727 19014 9773 19066
rect 9477 19012 9533 19014
rect 9557 19012 9613 19014
rect 9637 19012 9693 19014
rect 9717 19012 9773 19014
rect 9477 17978 9533 17980
rect 9557 17978 9613 17980
rect 9637 17978 9693 17980
rect 9717 17978 9773 17980
rect 9477 17926 9523 17978
rect 9523 17926 9533 17978
rect 9557 17926 9587 17978
rect 9587 17926 9599 17978
rect 9599 17926 9613 17978
rect 9637 17926 9651 17978
rect 9651 17926 9663 17978
rect 9663 17926 9693 17978
rect 9717 17926 9727 17978
rect 9727 17926 9773 17978
rect 9477 17924 9533 17926
rect 9557 17924 9613 17926
rect 9637 17924 9693 17926
rect 9717 17924 9773 17926
rect 9477 16890 9533 16892
rect 9557 16890 9613 16892
rect 9637 16890 9693 16892
rect 9717 16890 9773 16892
rect 9477 16838 9523 16890
rect 9523 16838 9533 16890
rect 9557 16838 9587 16890
rect 9587 16838 9599 16890
rect 9599 16838 9613 16890
rect 9637 16838 9651 16890
rect 9651 16838 9663 16890
rect 9663 16838 9693 16890
rect 9717 16838 9727 16890
rect 9727 16838 9773 16890
rect 9477 16836 9533 16838
rect 9557 16836 9613 16838
rect 9637 16836 9693 16838
rect 9717 16836 9773 16838
rect 9477 15802 9533 15804
rect 9557 15802 9613 15804
rect 9637 15802 9693 15804
rect 9717 15802 9773 15804
rect 9477 15750 9523 15802
rect 9523 15750 9533 15802
rect 9557 15750 9587 15802
rect 9587 15750 9599 15802
rect 9599 15750 9613 15802
rect 9637 15750 9651 15802
rect 9651 15750 9663 15802
rect 9663 15750 9693 15802
rect 9717 15750 9727 15802
rect 9727 15750 9773 15802
rect 9477 15748 9533 15750
rect 9557 15748 9613 15750
rect 9637 15748 9693 15750
rect 9717 15748 9773 15750
rect 9477 14714 9533 14716
rect 9557 14714 9613 14716
rect 9637 14714 9693 14716
rect 9717 14714 9773 14716
rect 9477 14662 9523 14714
rect 9523 14662 9533 14714
rect 9557 14662 9587 14714
rect 9587 14662 9599 14714
rect 9599 14662 9613 14714
rect 9637 14662 9651 14714
rect 9651 14662 9663 14714
rect 9663 14662 9693 14714
rect 9717 14662 9727 14714
rect 9727 14662 9773 14714
rect 9477 14660 9533 14662
rect 9557 14660 9613 14662
rect 9637 14660 9693 14662
rect 9717 14660 9773 14662
rect 9477 13626 9533 13628
rect 9557 13626 9613 13628
rect 9637 13626 9693 13628
rect 9717 13626 9773 13628
rect 9477 13574 9523 13626
rect 9523 13574 9533 13626
rect 9557 13574 9587 13626
rect 9587 13574 9599 13626
rect 9599 13574 9613 13626
rect 9637 13574 9651 13626
rect 9651 13574 9663 13626
rect 9663 13574 9693 13626
rect 9717 13574 9727 13626
rect 9727 13574 9773 13626
rect 9477 13572 9533 13574
rect 9557 13572 9613 13574
rect 9637 13572 9693 13574
rect 9717 13572 9773 13574
rect 9477 12538 9533 12540
rect 9557 12538 9613 12540
rect 9637 12538 9693 12540
rect 9717 12538 9773 12540
rect 9477 12486 9523 12538
rect 9523 12486 9533 12538
rect 9557 12486 9587 12538
rect 9587 12486 9599 12538
rect 9599 12486 9613 12538
rect 9637 12486 9651 12538
rect 9651 12486 9663 12538
rect 9663 12486 9693 12538
rect 9717 12486 9727 12538
rect 9727 12486 9773 12538
rect 9477 12484 9533 12486
rect 9557 12484 9613 12486
rect 9637 12484 9693 12486
rect 9717 12484 9773 12486
rect 10966 20868 11022 20904
rect 10966 20848 10968 20868
rect 10968 20848 11020 20868
rect 11020 20848 11022 20868
rect 9477 11450 9533 11452
rect 9557 11450 9613 11452
rect 9637 11450 9693 11452
rect 9717 11450 9773 11452
rect 9477 11398 9523 11450
rect 9523 11398 9533 11450
rect 9557 11398 9587 11450
rect 9587 11398 9599 11450
rect 9599 11398 9613 11450
rect 9637 11398 9651 11450
rect 9651 11398 9663 11450
rect 9663 11398 9693 11450
rect 9717 11398 9727 11450
rect 9727 11398 9773 11450
rect 9477 11396 9533 11398
rect 9557 11396 9613 11398
rect 9637 11396 9693 11398
rect 9717 11396 9773 11398
rect 9477 10362 9533 10364
rect 9557 10362 9613 10364
rect 9637 10362 9693 10364
rect 9717 10362 9773 10364
rect 9477 10310 9523 10362
rect 9523 10310 9533 10362
rect 9557 10310 9587 10362
rect 9587 10310 9599 10362
rect 9599 10310 9613 10362
rect 9637 10310 9651 10362
rect 9651 10310 9663 10362
rect 9663 10310 9693 10362
rect 9717 10310 9727 10362
rect 9727 10310 9773 10362
rect 9477 10308 9533 10310
rect 9557 10308 9613 10310
rect 9637 10308 9693 10310
rect 9717 10308 9773 10310
rect 9770 9560 9826 9616
rect 9477 9274 9533 9276
rect 9557 9274 9613 9276
rect 9637 9274 9693 9276
rect 9717 9274 9773 9276
rect 9477 9222 9523 9274
rect 9523 9222 9533 9274
rect 9557 9222 9587 9274
rect 9587 9222 9599 9274
rect 9599 9222 9613 9274
rect 9637 9222 9651 9274
rect 9651 9222 9663 9274
rect 9663 9222 9693 9274
rect 9717 9222 9727 9274
rect 9727 9222 9773 9274
rect 9477 9220 9533 9222
rect 9557 9220 9613 9222
rect 9637 9220 9693 9222
rect 9717 9220 9773 9222
rect 9477 8186 9533 8188
rect 9557 8186 9613 8188
rect 9637 8186 9693 8188
rect 9717 8186 9773 8188
rect 9477 8134 9523 8186
rect 9523 8134 9533 8186
rect 9557 8134 9587 8186
rect 9587 8134 9599 8186
rect 9599 8134 9613 8186
rect 9637 8134 9651 8186
rect 9651 8134 9663 8186
rect 9663 8134 9693 8186
rect 9717 8134 9727 8186
rect 9727 8134 9773 8186
rect 9477 8132 9533 8134
rect 9557 8132 9613 8134
rect 9637 8132 9693 8134
rect 9717 8132 9773 8134
rect 9477 7098 9533 7100
rect 9557 7098 9613 7100
rect 9637 7098 9693 7100
rect 9717 7098 9773 7100
rect 9477 7046 9523 7098
rect 9523 7046 9533 7098
rect 9557 7046 9587 7098
rect 9587 7046 9599 7098
rect 9599 7046 9613 7098
rect 9637 7046 9651 7098
rect 9651 7046 9663 7098
rect 9663 7046 9693 7098
rect 9717 7046 9727 7098
rect 9727 7046 9773 7098
rect 9477 7044 9533 7046
rect 9557 7044 9613 7046
rect 9637 7044 9693 7046
rect 9717 7044 9773 7046
rect 9477 6010 9533 6012
rect 9557 6010 9613 6012
rect 9637 6010 9693 6012
rect 9717 6010 9773 6012
rect 9477 5958 9523 6010
rect 9523 5958 9533 6010
rect 9557 5958 9587 6010
rect 9587 5958 9599 6010
rect 9599 5958 9613 6010
rect 9637 5958 9651 6010
rect 9651 5958 9663 6010
rect 9663 5958 9693 6010
rect 9717 5958 9727 6010
rect 9727 5958 9773 6010
rect 9477 5956 9533 5958
rect 9557 5956 9613 5958
rect 9637 5956 9693 5958
rect 9717 5956 9773 5958
rect 10230 9324 10232 9344
rect 10232 9324 10284 9344
rect 10284 9324 10286 9344
rect 10230 9288 10286 9324
rect 9477 4922 9533 4924
rect 9557 4922 9613 4924
rect 9637 4922 9693 4924
rect 9717 4922 9773 4924
rect 9477 4870 9523 4922
rect 9523 4870 9533 4922
rect 9557 4870 9587 4922
rect 9587 4870 9599 4922
rect 9599 4870 9613 4922
rect 9637 4870 9651 4922
rect 9651 4870 9663 4922
rect 9663 4870 9693 4922
rect 9717 4870 9727 4922
rect 9727 4870 9773 4922
rect 9477 4868 9533 4870
rect 9557 4868 9613 4870
rect 9637 4868 9693 4870
rect 9717 4868 9773 4870
rect 12317 21786 12373 21788
rect 12397 21786 12453 21788
rect 12477 21786 12533 21788
rect 12557 21786 12613 21788
rect 12317 21734 12363 21786
rect 12363 21734 12373 21786
rect 12397 21734 12427 21786
rect 12427 21734 12439 21786
rect 12439 21734 12453 21786
rect 12477 21734 12491 21786
rect 12491 21734 12503 21786
rect 12503 21734 12533 21786
rect 12557 21734 12567 21786
rect 12567 21734 12613 21786
rect 12317 21732 12373 21734
rect 12397 21732 12453 21734
rect 12477 21732 12533 21734
rect 12557 21732 12613 21734
rect 13174 21956 13230 21992
rect 13174 21936 13176 21956
rect 13176 21936 13228 21956
rect 13228 21936 13230 21956
rect 11242 13232 11298 13288
rect 10874 9324 10876 9344
rect 10876 9324 10928 9344
rect 10928 9324 10930 9344
rect 10874 9288 10930 9324
rect 10690 6024 10746 6080
rect 12530 21392 12586 21448
rect 12317 20698 12373 20700
rect 12397 20698 12453 20700
rect 12477 20698 12533 20700
rect 12557 20698 12613 20700
rect 12317 20646 12363 20698
rect 12363 20646 12373 20698
rect 12397 20646 12427 20698
rect 12427 20646 12439 20698
rect 12439 20646 12453 20698
rect 12477 20646 12491 20698
rect 12491 20646 12503 20698
rect 12503 20646 12533 20698
rect 12557 20646 12567 20698
rect 12567 20646 12613 20698
rect 12317 20644 12373 20646
rect 12397 20644 12453 20646
rect 12477 20644 12533 20646
rect 12557 20644 12613 20646
rect 12317 19610 12373 19612
rect 12397 19610 12453 19612
rect 12477 19610 12533 19612
rect 12557 19610 12613 19612
rect 12317 19558 12363 19610
rect 12363 19558 12373 19610
rect 12397 19558 12427 19610
rect 12427 19558 12439 19610
rect 12439 19558 12453 19610
rect 12477 19558 12491 19610
rect 12491 19558 12503 19610
rect 12503 19558 12533 19610
rect 12557 19558 12567 19610
rect 12567 19558 12613 19610
rect 12317 19556 12373 19558
rect 12397 19556 12453 19558
rect 12477 19556 12533 19558
rect 12557 19556 12613 19558
rect 12317 18522 12373 18524
rect 12397 18522 12453 18524
rect 12477 18522 12533 18524
rect 12557 18522 12613 18524
rect 12317 18470 12363 18522
rect 12363 18470 12373 18522
rect 12397 18470 12427 18522
rect 12427 18470 12439 18522
rect 12439 18470 12453 18522
rect 12477 18470 12491 18522
rect 12491 18470 12503 18522
rect 12503 18470 12533 18522
rect 12557 18470 12567 18522
rect 12567 18470 12613 18522
rect 12317 18468 12373 18470
rect 12397 18468 12453 18470
rect 12477 18468 12533 18470
rect 12557 18468 12613 18470
rect 12317 17434 12373 17436
rect 12397 17434 12453 17436
rect 12477 17434 12533 17436
rect 12557 17434 12613 17436
rect 12317 17382 12363 17434
rect 12363 17382 12373 17434
rect 12397 17382 12427 17434
rect 12427 17382 12439 17434
rect 12439 17382 12453 17434
rect 12477 17382 12491 17434
rect 12491 17382 12503 17434
rect 12503 17382 12533 17434
rect 12557 17382 12567 17434
rect 12567 17382 12613 17434
rect 12317 17380 12373 17382
rect 12397 17380 12453 17382
rect 12477 17380 12533 17382
rect 12557 17380 12613 17382
rect 13358 17620 13360 17640
rect 13360 17620 13412 17640
rect 13412 17620 13414 17640
rect 13358 17584 13414 17620
rect 12317 16346 12373 16348
rect 12397 16346 12453 16348
rect 12477 16346 12533 16348
rect 12557 16346 12613 16348
rect 12317 16294 12363 16346
rect 12363 16294 12373 16346
rect 12397 16294 12427 16346
rect 12427 16294 12439 16346
rect 12439 16294 12453 16346
rect 12477 16294 12491 16346
rect 12491 16294 12503 16346
rect 12503 16294 12533 16346
rect 12557 16294 12567 16346
rect 12567 16294 12613 16346
rect 12317 16292 12373 16294
rect 12397 16292 12453 16294
rect 12477 16292 12533 16294
rect 12557 16292 12613 16294
rect 11978 13232 12034 13288
rect 6636 2202 6692 2204
rect 6716 2202 6772 2204
rect 6796 2202 6852 2204
rect 6876 2202 6932 2204
rect 6636 2150 6682 2202
rect 6682 2150 6692 2202
rect 6716 2150 6746 2202
rect 6746 2150 6758 2202
rect 6758 2150 6772 2202
rect 6796 2150 6810 2202
rect 6810 2150 6822 2202
rect 6822 2150 6852 2202
rect 6876 2150 6886 2202
rect 6886 2150 6932 2202
rect 6636 2148 6692 2150
rect 6716 2148 6772 2150
rect 6796 2148 6852 2150
rect 6876 2148 6932 2150
rect 9477 3834 9533 3836
rect 9557 3834 9613 3836
rect 9637 3834 9693 3836
rect 9717 3834 9773 3836
rect 9477 3782 9523 3834
rect 9523 3782 9533 3834
rect 9557 3782 9587 3834
rect 9587 3782 9599 3834
rect 9599 3782 9613 3834
rect 9637 3782 9651 3834
rect 9651 3782 9663 3834
rect 9663 3782 9693 3834
rect 9717 3782 9727 3834
rect 9727 3782 9773 3834
rect 9477 3780 9533 3782
rect 9557 3780 9613 3782
rect 9637 3780 9693 3782
rect 9717 3780 9773 3782
rect 9477 2746 9533 2748
rect 9557 2746 9613 2748
rect 9637 2746 9693 2748
rect 9717 2746 9773 2748
rect 9477 2694 9523 2746
rect 9523 2694 9533 2746
rect 9557 2694 9587 2746
rect 9587 2694 9599 2746
rect 9599 2694 9613 2746
rect 9637 2694 9651 2746
rect 9651 2694 9663 2746
rect 9663 2694 9693 2746
rect 9717 2694 9727 2746
rect 9727 2694 9773 2746
rect 9477 2692 9533 2694
rect 9557 2692 9613 2694
rect 9637 2692 9693 2694
rect 9717 2692 9773 2694
rect 9954 3032 10010 3088
rect 11426 5208 11482 5264
rect 12317 15258 12373 15260
rect 12397 15258 12453 15260
rect 12477 15258 12533 15260
rect 12557 15258 12613 15260
rect 12317 15206 12363 15258
rect 12363 15206 12373 15258
rect 12397 15206 12427 15258
rect 12427 15206 12439 15258
rect 12439 15206 12453 15258
rect 12477 15206 12491 15258
rect 12491 15206 12503 15258
rect 12503 15206 12533 15258
rect 12557 15206 12567 15258
rect 12567 15206 12613 15258
rect 12317 15204 12373 15206
rect 12397 15204 12453 15206
rect 12477 15204 12533 15206
rect 12557 15204 12613 15206
rect 12317 14170 12373 14172
rect 12397 14170 12453 14172
rect 12477 14170 12533 14172
rect 12557 14170 12613 14172
rect 12317 14118 12363 14170
rect 12363 14118 12373 14170
rect 12397 14118 12427 14170
rect 12427 14118 12439 14170
rect 12439 14118 12453 14170
rect 12477 14118 12491 14170
rect 12491 14118 12503 14170
rect 12503 14118 12533 14170
rect 12557 14118 12567 14170
rect 12567 14118 12613 14170
rect 12317 14116 12373 14118
rect 12397 14116 12453 14118
rect 12477 14116 12533 14118
rect 12557 14116 12613 14118
rect 12317 13082 12373 13084
rect 12397 13082 12453 13084
rect 12477 13082 12533 13084
rect 12557 13082 12613 13084
rect 12317 13030 12363 13082
rect 12363 13030 12373 13082
rect 12397 13030 12427 13082
rect 12427 13030 12439 13082
rect 12439 13030 12453 13082
rect 12477 13030 12491 13082
rect 12491 13030 12503 13082
rect 12503 13030 12533 13082
rect 12557 13030 12567 13082
rect 12567 13030 12613 13082
rect 12317 13028 12373 13030
rect 12397 13028 12453 13030
rect 12477 13028 12533 13030
rect 12557 13028 12613 13030
rect 12317 11994 12373 11996
rect 12397 11994 12453 11996
rect 12477 11994 12533 11996
rect 12557 11994 12613 11996
rect 12317 11942 12363 11994
rect 12363 11942 12373 11994
rect 12397 11942 12427 11994
rect 12427 11942 12439 11994
rect 12439 11942 12453 11994
rect 12477 11942 12491 11994
rect 12491 11942 12503 11994
rect 12503 11942 12533 11994
rect 12557 11942 12567 11994
rect 12567 11942 12613 11994
rect 12317 11940 12373 11942
rect 12397 11940 12453 11942
rect 12477 11940 12533 11942
rect 12557 11940 12613 11942
rect 12317 10906 12373 10908
rect 12397 10906 12453 10908
rect 12477 10906 12533 10908
rect 12557 10906 12613 10908
rect 12317 10854 12363 10906
rect 12363 10854 12373 10906
rect 12397 10854 12427 10906
rect 12427 10854 12439 10906
rect 12439 10854 12453 10906
rect 12477 10854 12491 10906
rect 12491 10854 12503 10906
rect 12503 10854 12533 10906
rect 12557 10854 12567 10906
rect 12567 10854 12613 10906
rect 12317 10852 12373 10854
rect 12397 10852 12453 10854
rect 12477 10852 12533 10854
rect 12557 10852 12613 10854
rect 12317 9818 12373 9820
rect 12397 9818 12453 9820
rect 12477 9818 12533 9820
rect 12557 9818 12613 9820
rect 12317 9766 12363 9818
rect 12363 9766 12373 9818
rect 12397 9766 12427 9818
rect 12427 9766 12439 9818
rect 12439 9766 12453 9818
rect 12477 9766 12491 9818
rect 12491 9766 12503 9818
rect 12503 9766 12533 9818
rect 12557 9766 12567 9818
rect 12567 9766 12613 9818
rect 12317 9764 12373 9766
rect 12397 9764 12453 9766
rect 12477 9764 12533 9766
rect 12557 9764 12613 9766
rect 12162 9560 12218 9616
rect 12317 8730 12373 8732
rect 12397 8730 12453 8732
rect 12477 8730 12533 8732
rect 12557 8730 12613 8732
rect 12317 8678 12363 8730
rect 12363 8678 12373 8730
rect 12397 8678 12427 8730
rect 12427 8678 12439 8730
rect 12439 8678 12453 8730
rect 12477 8678 12491 8730
rect 12491 8678 12503 8730
rect 12503 8678 12533 8730
rect 12557 8678 12567 8730
rect 12567 8678 12613 8730
rect 12317 8676 12373 8678
rect 12397 8676 12453 8678
rect 12477 8676 12533 8678
rect 12557 8676 12613 8678
rect 12317 7642 12373 7644
rect 12397 7642 12453 7644
rect 12477 7642 12533 7644
rect 12557 7642 12613 7644
rect 12317 7590 12363 7642
rect 12363 7590 12373 7642
rect 12397 7590 12427 7642
rect 12427 7590 12439 7642
rect 12439 7590 12453 7642
rect 12477 7590 12491 7642
rect 12491 7590 12503 7642
rect 12503 7590 12533 7642
rect 12557 7590 12567 7642
rect 12567 7590 12613 7642
rect 12317 7588 12373 7590
rect 12397 7588 12453 7590
rect 12477 7588 12533 7590
rect 12557 7588 12613 7590
rect 11426 3460 11482 3496
rect 11426 3440 11428 3460
rect 11428 3440 11480 3460
rect 11480 3440 11482 3460
rect 11702 3304 11758 3360
rect 11794 3168 11850 3224
rect 13542 19236 13598 19272
rect 13542 19216 13544 19236
rect 13544 19216 13596 19236
rect 13596 19216 13598 19236
rect 13358 13368 13414 13424
rect 14186 21256 14242 21312
rect 15158 21242 15214 21244
rect 15238 21242 15294 21244
rect 15318 21242 15374 21244
rect 15398 21242 15454 21244
rect 15158 21190 15204 21242
rect 15204 21190 15214 21242
rect 15238 21190 15268 21242
rect 15268 21190 15280 21242
rect 15280 21190 15294 21242
rect 15318 21190 15332 21242
rect 15332 21190 15344 21242
rect 15344 21190 15374 21242
rect 15398 21190 15408 21242
rect 15408 21190 15454 21242
rect 15158 21188 15214 21190
rect 15238 21188 15294 21190
rect 15318 21188 15374 21190
rect 15398 21188 15454 21190
rect 20839 22330 20895 22332
rect 20919 22330 20975 22332
rect 20999 22330 21055 22332
rect 21079 22330 21135 22332
rect 20839 22278 20885 22330
rect 20885 22278 20895 22330
rect 20919 22278 20949 22330
rect 20949 22278 20961 22330
rect 20961 22278 20975 22330
rect 20999 22278 21013 22330
rect 21013 22278 21025 22330
rect 21025 22278 21055 22330
rect 21079 22278 21089 22330
rect 21089 22278 21135 22330
rect 20839 22276 20895 22278
rect 20919 22276 20975 22278
rect 20999 22276 21055 22278
rect 21079 22276 21135 22278
rect 20442 21972 20444 21992
rect 20444 21972 20496 21992
rect 20496 21972 20498 21992
rect 20442 21936 20498 21972
rect 17998 21786 18054 21788
rect 18078 21786 18134 21788
rect 18158 21786 18214 21788
rect 18238 21786 18294 21788
rect 17998 21734 18044 21786
rect 18044 21734 18054 21786
rect 18078 21734 18108 21786
rect 18108 21734 18120 21786
rect 18120 21734 18134 21786
rect 18158 21734 18172 21786
rect 18172 21734 18184 21786
rect 18184 21734 18214 21786
rect 18238 21734 18248 21786
rect 18248 21734 18294 21786
rect 17998 21732 18054 21734
rect 18078 21732 18134 21734
rect 18158 21732 18214 21734
rect 18238 21732 18294 21734
rect 14738 18808 14794 18864
rect 14462 17076 14464 17096
rect 14464 17076 14516 17096
rect 14516 17076 14518 17096
rect 14462 17040 14518 17076
rect 15158 20154 15214 20156
rect 15238 20154 15294 20156
rect 15318 20154 15374 20156
rect 15398 20154 15454 20156
rect 15158 20102 15204 20154
rect 15204 20102 15214 20154
rect 15238 20102 15268 20154
rect 15268 20102 15280 20154
rect 15280 20102 15294 20154
rect 15318 20102 15332 20154
rect 15332 20102 15344 20154
rect 15344 20102 15374 20154
rect 15398 20102 15408 20154
rect 15408 20102 15454 20154
rect 15158 20100 15214 20102
rect 15238 20100 15294 20102
rect 15318 20100 15374 20102
rect 15398 20100 15454 20102
rect 15158 19066 15214 19068
rect 15238 19066 15294 19068
rect 15318 19066 15374 19068
rect 15398 19066 15454 19068
rect 15158 19014 15204 19066
rect 15204 19014 15214 19066
rect 15238 19014 15268 19066
rect 15268 19014 15280 19066
rect 15280 19014 15294 19066
rect 15318 19014 15332 19066
rect 15332 19014 15344 19066
rect 15344 19014 15374 19066
rect 15398 19014 15408 19066
rect 15408 19014 15454 19066
rect 15158 19012 15214 19014
rect 15238 19012 15294 19014
rect 15318 19012 15374 19014
rect 15398 19012 15454 19014
rect 15014 18164 15016 18184
rect 15016 18164 15068 18184
rect 15068 18164 15070 18184
rect 15014 18128 15070 18164
rect 15158 17978 15214 17980
rect 15238 17978 15294 17980
rect 15318 17978 15374 17980
rect 15398 17978 15454 17980
rect 15158 17926 15204 17978
rect 15204 17926 15214 17978
rect 15238 17926 15268 17978
rect 15268 17926 15280 17978
rect 15280 17926 15294 17978
rect 15318 17926 15332 17978
rect 15332 17926 15344 17978
rect 15344 17926 15374 17978
rect 15398 17926 15408 17978
rect 15408 17926 15454 17978
rect 15158 17924 15214 17926
rect 15238 17924 15294 17926
rect 15318 17924 15374 17926
rect 15398 17924 15454 17926
rect 14830 16496 14886 16552
rect 15106 17584 15162 17640
rect 15158 16890 15214 16892
rect 15238 16890 15294 16892
rect 15318 16890 15374 16892
rect 15398 16890 15454 16892
rect 15158 16838 15204 16890
rect 15204 16838 15214 16890
rect 15238 16838 15268 16890
rect 15268 16838 15280 16890
rect 15280 16838 15294 16890
rect 15318 16838 15332 16890
rect 15332 16838 15344 16890
rect 15344 16838 15374 16890
rect 15398 16838 15408 16890
rect 15408 16838 15454 16890
rect 15158 16836 15214 16838
rect 15238 16836 15294 16838
rect 15318 16836 15374 16838
rect 15398 16836 15454 16838
rect 15014 15988 15016 16008
rect 15016 15988 15068 16008
rect 15068 15988 15070 16008
rect 15014 15952 15070 15988
rect 15842 19216 15898 19272
rect 15158 15802 15214 15804
rect 15238 15802 15294 15804
rect 15318 15802 15374 15804
rect 15398 15802 15454 15804
rect 15158 15750 15204 15802
rect 15204 15750 15214 15802
rect 15238 15750 15268 15802
rect 15268 15750 15280 15802
rect 15280 15750 15294 15802
rect 15318 15750 15332 15802
rect 15332 15750 15344 15802
rect 15344 15750 15374 15802
rect 15398 15750 15408 15802
rect 15408 15750 15454 15802
rect 15158 15748 15214 15750
rect 15238 15748 15294 15750
rect 15318 15748 15374 15750
rect 15398 15748 15454 15750
rect 14462 13776 14518 13832
rect 14462 12824 14518 12880
rect 15158 14714 15214 14716
rect 15238 14714 15294 14716
rect 15318 14714 15374 14716
rect 15398 14714 15454 14716
rect 15158 14662 15204 14714
rect 15204 14662 15214 14714
rect 15238 14662 15268 14714
rect 15268 14662 15280 14714
rect 15280 14662 15294 14714
rect 15318 14662 15332 14714
rect 15332 14662 15344 14714
rect 15344 14662 15374 14714
rect 15398 14662 15408 14714
rect 15408 14662 15454 14714
rect 15158 14660 15214 14662
rect 15238 14660 15294 14662
rect 15318 14660 15374 14662
rect 15398 14660 15454 14662
rect 15158 13626 15214 13628
rect 15238 13626 15294 13628
rect 15318 13626 15374 13628
rect 15398 13626 15454 13628
rect 15158 13574 15204 13626
rect 15204 13574 15214 13626
rect 15238 13574 15268 13626
rect 15268 13574 15280 13626
rect 15280 13574 15294 13626
rect 15318 13574 15332 13626
rect 15332 13574 15344 13626
rect 15344 13574 15374 13626
rect 15398 13574 15408 13626
rect 15408 13574 15454 13626
rect 15158 13572 15214 13574
rect 15238 13572 15294 13574
rect 15318 13572 15374 13574
rect 15398 13572 15454 13574
rect 15158 12538 15214 12540
rect 15238 12538 15294 12540
rect 15318 12538 15374 12540
rect 15398 12538 15454 12540
rect 15158 12486 15204 12538
rect 15204 12486 15214 12538
rect 15238 12486 15268 12538
rect 15268 12486 15280 12538
rect 15280 12486 15294 12538
rect 15318 12486 15332 12538
rect 15332 12486 15344 12538
rect 15344 12486 15374 12538
rect 15398 12486 15408 12538
rect 15408 12486 15454 12538
rect 15158 12484 15214 12486
rect 15238 12484 15294 12486
rect 15318 12484 15374 12486
rect 15398 12484 15454 12486
rect 15382 11736 15438 11792
rect 15158 11450 15214 11452
rect 15238 11450 15294 11452
rect 15318 11450 15374 11452
rect 15398 11450 15454 11452
rect 15158 11398 15204 11450
rect 15204 11398 15214 11450
rect 15238 11398 15268 11450
rect 15268 11398 15280 11450
rect 15280 11398 15294 11450
rect 15318 11398 15332 11450
rect 15332 11398 15344 11450
rect 15344 11398 15374 11450
rect 15398 11398 15408 11450
rect 15408 11398 15454 11450
rect 15158 11396 15214 11398
rect 15238 11396 15294 11398
rect 15318 11396 15374 11398
rect 15398 11396 15454 11398
rect 15198 10512 15254 10568
rect 15158 10362 15214 10364
rect 15238 10362 15294 10364
rect 15318 10362 15374 10364
rect 15398 10362 15454 10364
rect 15158 10310 15204 10362
rect 15204 10310 15214 10362
rect 15238 10310 15268 10362
rect 15268 10310 15280 10362
rect 15280 10310 15294 10362
rect 15318 10310 15332 10362
rect 15332 10310 15344 10362
rect 15344 10310 15374 10362
rect 15398 10310 15408 10362
rect 15408 10310 15454 10362
rect 15158 10308 15214 10310
rect 15238 10308 15294 10310
rect 15318 10308 15374 10310
rect 15398 10308 15454 10310
rect 17998 20698 18054 20700
rect 18078 20698 18134 20700
rect 18158 20698 18214 20700
rect 18238 20698 18294 20700
rect 17998 20646 18044 20698
rect 18044 20646 18054 20698
rect 18078 20646 18108 20698
rect 18108 20646 18120 20698
rect 18120 20646 18134 20698
rect 18158 20646 18172 20698
rect 18172 20646 18184 20698
rect 18184 20646 18214 20698
rect 18238 20646 18248 20698
rect 18248 20646 18294 20698
rect 17998 20644 18054 20646
rect 18078 20644 18134 20646
rect 18158 20644 18214 20646
rect 18238 20644 18294 20646
rect 17998 19610 18054 19612
rect 18078 19610 18134 19612
rect 18158 19610 18214 19612
rect 18238 19610 18294 19612
rect 17998 19558 18044 19610
rect 18044 19558 18054 19610
rect 18078 19558 18108 19610
rect 18108 19558 18120 19610
rect 18120 19558 18134 19610
rect 18158 19558 18172 19610
rect 18172 19558 18184 19610
rect 18184 19558 18214 19610
rect 18238 19558 18248 19610
rect 18248 19558 18294 19610
rect 17998 19556 18054 19558
rect 18078 19556 18134 19558
rect 18158 19556 18214 19558
rect 18238 19556 18294 19558
rect 16486 17584 16542 17640
rect 16670 15136 16726 15192
rect 16578 13096 16634 13152
rect 12317 6554 12373 6556
rect 12397 6554 12453 6556
rect 12477 6554 12533 6556
rect 12557 6554 12613 6556
rect 12317 6502 12363 6554
rect 12363 6502 12373 6554
rect 12397 6502 12427 6554
rect 12427 6502 12439 6554
rect 12439 6502 12453 6554
rect 12477 6502 12491 6554
rect 12491 6502 12503 6554
rect 12503 6502 12533 6554
rect 12557 6502 12567 6554
rect 12567 6502 12613 6554
rect 12317 6500 12373 6502
rect 12397 6500 12453 6502
rect 12477 6500 12533 6502
rect 12557 6500 12613 6502
rect 12317 5466 12373 5468
rect 12397 5466 12453 5468
rect 12477 5466 12533 5468
rect 12557 5466 12613 5468
rect 12317 5414 12363 5466
rect 12363 5414 12373 5466
rect 12397 5414 12427 5466
rect 12427 5414 12439 5466
rect 12439 5414 12453 5466
rect 12477 5414 12491 5466
rect 12491 5414 12503 5466
rect 12503 5414 12533 5466
rect 12557 5414 12567 5466
rect 12567 5414 12613 5466
rect 12317 5412 12373 5414
rect 12397 5412 12453 5414
rect 12477 5412 12533 5414
rect 12557 5412 12613 5414
rect 12254 5072 12310 5128
rect 12317 4378 12373 4380
rect 12397 4378 12453 4380
rect 12477 4378 12533 4380
rect 12557 4378 12613 4380
rect 12317 4326 12363 4378
rect 12363 4326 12373 4378
rect 12397 4326 12427 4378
rect 12427 4326 12439 4378
rect 12439 4326 12453 4378
rect 12477 4326 12491 4378
rect 12491 4326 12503 4378
rect 12503 4326 12533 4378
rect 12557 4326 12567 4378
rect 12567 4326 12613 4378
rect 12317 4324 12373 4326
rect 12397 4324 12453 4326
rect 12477 4324 12533 4326
rect 12557 4324 12613 4326
rect 12317 3290 12373 3292
rect 12397 3290 12453 3292
rect 12477 3290 12533 3292
rect 12557 3290 12613 3292
rect 12317 3238 12363 3290
rect 12363 3238 12373 3290
rect 12397 3238 12427 3290
rect 12427 3238 12439 3290
rect 12439 3238 12453 3290
rect 12477 3238 12491 3290
rect 12491 3238 12503 3290
rect 12503 3238 12533 3290
rect 12557 3238 12567 3290
rect 12567 3238 12613 3290
rect 12317 3236 12373 3238
rect 12397 3236 12453 3238
rect 12477 3236 12533 3238
rect 12557 3236 12613 3238
rect 13542 4120 13598 4176
rect 14002 6060 14004 6080
rect 14004 6060 14056 6080
rect 14056 6060 14058 6080
rect 14002 6024 14058 6060
rect 13726 3052 13782 3088
rect 13726 3032 13728 3052
rect 13728 3032 13780 3052
rect 13780 3032 13782 3052
rect 12317 2202 12373 2204
rect 12397 2202 12453 2204
rect 12477 2202 12533 2204
rect 12557 2202 12613 2204
rect 12317 2150 12363 2202
rect 12363 2150 12373 2202
rect 12397 2150 12427 2202
rect 12427 2150 12439 2202
rect 12439 2150 12453 2202
rect 12477 2150 12491 2202
rect 12491 2150 12503 2202
rect 12503 2150 12533 2202
rect 12557 2150 12567 2202
rect 12567 2150 12613 2202
rect 12317 2148 12373 2150
rect 12397 2148 12453 2150
rect 12477 2148 12533 2150
rect 12557 2148 12613 2150
rect 14554 2896 14610 2952
rect 15158 9274 15214 9276
rect 15238 9274 15294 9276
rect 15318 9274 15374 9276
rect 15398 9274 15454 9276
rect 15158 9222 15204 9274
rect 15204 9222 15214 9274
rect 15238 9222 15268 9274
rect 15268 9222 15280 9274
rect 15280 9222 15294 9274
rect 15318 9222 15332 9274
rect 15332 9222 15344 9274
rect 15344 9222 15374 9274
rect 15398 9222 15408 9274
rect 15408 9222 15454 9274
rect 15158 9220 15214 9222
rect 15238 9220 15294 9222
rect 15318 9220 15374 9222
rect 15398 9220 15454 9222
rect 15158 8186 15214 8188
rect 15238 8186 15294 8188
rect 15318 8186 15374 8188
rect 15398 8186 15454 8188
rect 15158 8134 15204 8186
rect 15204 8134 15214 8186
rect 15238 8134 15268 8186
rect 15268 8134 15280 8186
rect 15280 8134 15294 8186
rect 15318 8134 15332 8186
rect 15332 8134 15344 8186
rect 15344 8134 15374 8186
rect 15398 8134 15408 8186
rect 15408 8134 15454 8186
rect 15158 8132 15214 8134
rect 15238 8132 15294 8134
rect 15318 8132 15374 8134
rect 15398 8132 15454 8134
rect 15158 7098 15214 7100
rect 15238 7098 15294 7100
rect 15318 7098 15374 7100
rect 15398 7098 15454 7100
rect 15158 7046 15204 7098
rect 15204 7046 15214 7098
rect 15238 7046 15268 7098
rect 15268 7046 15280 7098
rect 15280 7046 15294 7098
rect 15318 7046 15332 7098
rect 15332 7046 15344 7098
rect 15344 7046 15374 7098
rect 15398 7046 15408 7098
rect 15408 7046 15454 7098
rect 15158 7044 15214 7046
rect 15238 7044 15294 7046
rect 15318 7044 15374 7046
rect 15398 7044 15454 7046
rect 15158 6010 15214 6012
rect 15238 6010 15294 6012
rect 15318 6010 15374 6012
rect 15398 6010 15454 6012
rect 15158 5958 15204 6010
rect 15204 5958 15214 6010
rect 15238 5958 15268 6010
rect 15268 5958 15280 6010
rect 15280 5958 15294 6010
rect 15318 5958 15332 6010
rect 15332 5958 15344 6010
rect 15344 5958 15374 6010
rect 15398 5958 15408 6010
rect 15408 5958 15454 6010
rect 15158 5956 15214 5958
rect 15238 5956 15294 5958
rect 15318 5956 15374 5958
rect 15398 5956 15454 5958
rect 15158 4922 15214 4924
rect 15238 4922 15294 4924
rect 15318 4922 15374 4924
rect 15398 4922 15454 4924
rect 15158 4870 15204 4922
rect 15204 4870 15214 4922
rect 15238 4870 15268 4922
rect 15268 4870 15280 4922
rect 15280 4870 15294 4922
rect 15318 4870 15332 4922
rect 15332 4870 15344 4922
rect 15344 4870 15374 4922
rect 15398 4870 15408 4922
rect 15408 4870 15454 4922
rect 15158 4868 15214 4870
rect 15238 4868 15294 4870
rect 15318 4868 15374 4870
rect 15398 4868 15454 4870
rect 15158 3834 15214 3836
rect 15238 3834 15294 3836
rect 15318 3834 15374 3836
rect 15398 3834 15454 3836
rect 15158 3782 15204 3834
rect 15204 3782 15214 3834
rect 15238 3782 15268 3834
rect 15268 3782 15280 3834
rect 15280 3782 15294 3834
rect 15318 3782 15332 3834
rect 15332 3782 15344 3834
rect 15344 3782 15374 3834
rect 15398 3782 15408 3834
rect 15408 3782 15454 3834
rect 15158 3780 15214 3782
rect 15238 3780 15294 3782
rect 15318 3780 15374 3782
rect 15398 3780 15454 3782
rect 14922 3576 14978 3632
rect 15158 2746 15214 2748
rect 15238 2746 15294 2748
rect 15318 2746 15374 2748
rect 15398 2746 15454 2748
rect 15158 2694 15204 2746
rect 15204 2694 15214 2746
rect 15238 2694 15268 2746
rect 15268 2694 15280 2746
rect 15280 2694 15294 2746
rect 15318 2694 15332 2746
rect 15332 2694 15344 2746
rect 15344 2694 15374 2746
rect 15398 2694 15408 2746
rect 15408 2694 15454 2746
rect 15158 2692 15214 2694
rect 15238 2692 15294 2694
rect 15318 2692 15374 2694
rect 15398 2692 15454 2694
rect 16854 13796 16910 13832
rect 16854 13776 16856 13796
rect 16856 13776 16908 13796
rect 16908 13776 16910 13796
rect 17998 18522 18054 18524
rect 18078 18522 18134 18524
rect 18158 18522 18214 18524
rect 18238 18522 18294 18524
rect 17998 18470 18044 18522
rect 18044 18470 18054 18522
rect 18078 18470 18108 18522
rect 18108 18470 18120 18522
rect 18120 18470 18134 18522
rect 18158 18470 18172 18522
rect 18172 18470 18184 18522
rect 18184 18470 18214 18522
rect 18238 18470 18248 18522
rect 18248 18470 18294 18522
rect 17998 18468 18054 18470
rect 18078 18468 18134 18470
rect 18158 18468 18214 18470
rect 18238 18468 18294 18470
rect 17682 18128 17738 18184
rect 17222 12844 17278 12880
rect 17222 12824 17224 12844
rect 17224 12824 17276 12844
rect 17276 12824 17278 12844
rect 17130 12280 17186 12336
rect 17038 11092 17040 11112
rect 17040 11092 17092 11112
rect 17092 11092 17094 11112
rect 17038 11056 17094 11092
rect 15842 5228 15898 5264
rect 15842 5208 15844 5228
rect 15844 5208 15896 5228
rect 15896 5208 15898 5228
rect 15934 4120 15990 4176
rect 17998 17434 18054 17436
rect 18078 17434 18134 17436
rect 18158 17434 18214 17436
rect 18238 17434 18294 17436
rect 17998 17382 18044 17434
rect 18044 17382 18054 17434
rect 18078 17382 18108 17434
rect 18108 17382 18120 17434
rect 18120 17382 18134 17434
rect 18158 17382 18172 17434
rect 18172 17382 18184 17434
rect 18184 17382 18214 17434
rect 18238 17382 18248 17434
rect 18248 17382 18294 17434
rect 17998 17380 18054 17382
rect 18078 17380 18134 17382
rect 18158 17380 18214 17382
rect 18238 17380 18294 17382
rect 17998 16346 18054 16348
rect 18078 16346 18134 16348
rect 18158 16346 18214 16348
rect 18238 16346 18294 16348
rect 17998 16294 18044 16346
rect 18044 16294 18054 16346
rect 18078 16294 18108 16346
rect 18108 16294 18120 16346
rect 18120 16294 18134 16346
rect 18158 16294 18172 16346
rect 18172 16294 18184 16346
rect 18184 16294 18214 16346
rect 18238 16294 18248 16346
rect 18248 16294 18294 16346
rect 17998 16292 18054 16294
rect 18078 16292 18134 16294
rect 18158 16292 18214 16294
rect 18238 16292 18294 16294
rect 17998 15258 18054 15260
rect 18078 15258 18134 15260
rect 18158 15258 18214 15260
rect 18238 15258 18294 15260
rect 17998 15206 18044 15258
rect 18044 15206 18054 15258
rect 18078 15206 18108 15258
rect 18108 15206 18120 15258
rect 18120 15206 18134 15258
rect 18158 15206 18172 15258
rect 18172 15206 18184 15258
rect 18184 15206 18214 15258
rect 18238 15206 18248 15258
rect 18248 15206 18294 15258
rect 17998 15204 18054 15206
rect 18078 15204 18134 15206
rect 18158 15204 18214 15206
rect 18238 15204 18294 15206
rect 17682 13096 17738 13152
rect 16302 4140 16358 4176
rect 16302 4120 16304 4140
rect 16304 4120 16356 4140
rect 16356 4120 16358 4140
rect 17998 14170 18054 14172
rect 18078 14170 18134 14172
rect 18158 14170 18214 14172
rect 18238 14170 18294 14172
rect 17998 14118 18044 14170
rect 18044 14118 18054 14170
rect 18078 14118 18108 14170
rect 18108 14118 18120 14170
rect 18120 14118 18134 14170
rect 18158 14118 18172 14170
rect 18172 14118 18184 14170
rect 18184 14118 18214 14170
rect 18238 14118 18248 14170
rect 18248 14118 18294 14170
rect 17998 14116 18054 14118
rect 18078 14116 18134 14118
rect 18158 14116 18214 14118
rect 18238 14116 18294 14118
rect 17998 13082 18054 13084
rect 18078 13082 18134 13084
rect 18158 13082 18214 13084
rect 18238 13082 18294 13084
rect 17998 13030 18044 13082
rect 18044 13030 18054 13082
rect 18078 13030 18108 13082
rect 18108 13030 18120 13082
rect 18120 13030 18134 13082
rect 18158 13030 18172 13082
rect 18172 13030 18184 13082
rect 18184 13030 18214 13082
rect 18238 13030 18248 13082
rect 18248 13030 18294 13082
rect 17998 13028 18054 13030
rect 18078 13028 18134 13030
rect 18158 13028 18214 13030
rect 18238 13028 18294 13030
rect 18602 17040 18658 17096
rect 19522 21392 19578 21448
rect 19614 20712 19670 20768
rect 17998 11994 18054 11996
rect 18078 11994 18134 11996
rect 18158 11994 18214 11996
rect 18238 11994 18294 11996
rect 17998 11942 18044 11994
rect 18044 11942 18054 11994
rect 18078 11942 18108 11994
rect 18108 11942 18120 11994
rect 18120 11942 18134 11994
rect 18158 11942 18172 11994
rect 18172 11942 18184 11994
rect 18184 11942 18214 11994
rect 18238 11942 18248 11994
rect 18248 11942 18294 11994
rect 17998 11940 18054 11942
rect 18078 11940 18134 11942
rect 18158 11940 18214 11942
rect 18238 11940 18294 11942
rect 17866 11736 17922 11792
rect 18786 13268 18788 13288
rect 18788 13268 18840 13288
rect 18840 13268 18842 13288
rect 18786 13232 18842 13268
rect 17998 10906 18054 10908
rect 18078 10906 18134 10908
rect 18158 10906 18214 10908
rect 18238 10906 18294 10908
rect 17998 10854 18044 10906
rect 18044 10854 18054 10906
rect 18078 10854 18108 10906
rect 18108 10854 18120 10906
rect 18120 10854 18134 10906
rect 18158 10854 18172 10906
rect 18172 10854 18184 10906
rect 18184 10854 18214 10906
rect 18238 10854 18248 10906
rect 18248 10854 18294 10906
rect 17998 10852 18054 10854
rect 18078 10852 18134 10854
rect 18158 10852 18214 10854
rect 18238 10852 18294 10854
rect 17774 9832 17830 9888
rect 17998 9818 18054 9820
rect 18078 9818 18134 9820
rect 18158 9818 18214 9820
rect 18238 9818 18294 9820
rect 17998 9766 18044 9818
rect 18044 9766 18054 9818
rect 18078 9766 18108 9818
rect 18108 9766 18120 9818
rect 18120 9766 18134 9818
rect 18158 9766 18172 9818
rect 18172 9766 18184 9818
rect 18184 9766 18214 9818
rect 18238 9766 18248 9818
rect 18248 9766 18294 9818
rect 17998 9764 18054 9766
rect 18078 9764 18134 9766
rect 18158 9764 18214 9766
rect 18238 9764 18294 9766
rect 17958 9632 18014 9688
rect 17998 8730 18054 8732
rect 18078 8730 18134 8732
rect 18158 8730 18214 8732
rect 18238 8730 18294 8732
rect 17998 8678 18044 8730
rect 18044 8678 18054 8730
rect 18078 8678 18108 8730
rect 18108 8678 18120 8730
rect 18120 8678 18134 8730
rect 18158 8678 18172 8730
rect 18172 8678 18184 8730
rect 18184 8678 18214 8730
rect 18238 8678 18248 8730
rect 18248 8678 18294 8730
rect 17998 8676 18054 8678
rect 18078 8676 18134 8678
rect 18158 8676 18214 8678
rect 18238 8676 18294 8678
rect 17998 7642 18054 7644
rect 18078 7642 18134 7644
rect 18158 7642 18214 7644
rect 18238 7642 18294 7644
rect 17998 7590 18044 7642
rect 18044 7590 18054 7642
rect 18078 7590 18108 7642
rect 18108 7590 18120 7642
rect 18120 7590 18134 7642
rect 18158 7590 18172 7642
rect 18172 7590 18184 7642
rect 18184 7590 18214 7642
rect 18238 7590 18248 7642
rect 18248 7590 18294 7642
rect 17998 7588 18054 7590
rect 18078 7588 18134 7590
rect 18158 7588 18214 7590
rect 18238 7588 18294 7590
rect 17998 6554 18054 6556
rect 18078 6554 18134 6556
rect 18158 6554 18214 6556
rect 18238 6554 18294 6556
rect 17998 6502 18044 6554
rect 18044 6502 18054 6554
rect 18078 6502 18108 6554
rect 18108 6502 18120 6554
rect 18120 6502 18134 6554
rect 18158 6502 18172 6554
rect 18172 6502 18184 6554
rect 18184 6502 18214 6554
rect 18238 6502 18248 6554
rect 18248 6502 18294 6554
rect 17998 6500 18054 6502
rect 18078 6500 18134 6502
rect 18158 6500 18214 6502
rect 18238 6500 18294 6502
rect 18694 6704 18750 6760
rect 17998 5466 18054 5468
rect 18078 5466 18134 5468
rect 18158 5466 18214 5468
rect 18238 5466 18294 5468
rect 17998 5414 18044 5466
rect 18044 5414 18054 5466
rect 18078 5414 18108 5466
rect 18108 5414 18120 5466
rect 18120 5414 18134 5466
rect 18158 5414 18172 5466
rect 18172 5414 18184 5466
rect 18184 5414 18214 5466
rect 18238 5414 18248 5466
rect 18248 5414 18294 5466
rect 17998 5412 18054 5414
rect 18078 5412 18134 5414
rect 18158 5412 18214 5414
rect 18238 5412 18294 5414
rect 17998 4378 18054 4380
rect 18078 4378 18134 4380
rect 18158 4378 18214 4380
rect 18238 4378 18294 4380
rect 17998 4326 18044 4378
rect 18044 4326 18054 4378
rect 18078 4326 18108 4378
rect 18108 4326 18120 4378
rect 18120 4326 18134 4378
rect 18158 4326 18172 4378
rect 18172 4326 18184 4378
rect 18184 4326 18214 4378
rect 18238 4326 18248 4378
rect 18248 4326 18294 4378
rect 17998 4324 18054 4326
rect 18078 4324 18134 4326
rect 18158 4324 18214 4326
rect 18238 4324 18294 4326
rect 18418 5072 18474 5128
rect 19062 15988 19064 16008
rect 19064 15988 19116 16008
rect 19116 15988 19118 16008
rect 19062 15952 19118 15988
rect 19430 16496 19486 16552
rect 20839 21242 20895 21244
rect 20919 21242 20975 21244
rect 20999 21242 21055 21244
rect 21079 21242 21135 21244
rect 20839 21190 20885 21242
rect 20885 21190 20895 21242
rect 20919 21190 20949 21242
rect 20949 21190 20961 21242
rect 20961 21190 20975 21242
rect 20999 21190 21013 21242
rect 21013 21190 21025 21242
rect 21025 21190 21055 21242
rect 21079 21190 21089 21242
rect 21089 21190 21135 21242
rect 20839 21188 20895 21190
rect 20919 21188 20975 21190
rect 20999 21188 21055 21190
rect 21079 21188 21135 21190
rect 21914 20868 21970 20904
rect 21914 20848 21916 20868
rect 21916 20848 21968 20868
rect 21968 20848 21970 20868
rect 19890 17992 19946 18048
rect 19154 12824 19210 12880
rect 19338 12300 19394 12336
rect 19338 12280 19340 12300
rect 19340 12280 19392 12300
rect 19392 12280 19394 12300
rect 23679 21786 23735 21788
rect 23759 21786 23815 21788
rect 23839 21786 23895 21788
rect 23919 21786 23975 21788
rect 23679 21734 23725 21786
rect 23725 21734 23735 21786
rect 23759 21734 23789 21786
rect 23789 21734 23801 21786
rect 23801 21734 23815 21786
rect 23839 21734 23853 21786
rect 23853 21734 23865 21786
rect 23865 21734 23895 21786
rect 23919 21734 23929 21786
rect 23929 21734 23975 21786
rect 23679 21732 23735 21734
rect 23759 21732 23815 21734
rect 23839 21732 23895 21734
rect 23919 21732 23975 21734
rect 23679 20698 23735 20700
rect 23759 20698 23815 20700
rect 23839 20698 23895 20700
rect 23919 20698 23975 20700
rect 23679 20646 23725 20698
rect 23725 20646 23735 20698
rect 23759 20646 23789 20698
rect 23789 20646 23801 20698
rect 23801 20646 23815 20698
rect 23839 20646 23853 20698
rect 23853 20646 23865 20698
rect 23865 20646 23895 20698
rect 23919 20646 23929 20698
rect 23929 20646 23975 20698
rect 23679 20644 23735 20646
rect 23759 20644 23815 20646
rect 23839 20644 23895 20646
rect 23919 20644 23975 20646
rect 19338 10512 19394 10568
rect 18970 8336 19026 8392
rect 20839 20154 20895 20156
rect 20919 20154 20975 20156
rect 20999 20154 21055 20156
rect 21079 20154 21135 20156
rect 20839 20102 20885 20154
rect 20885 20102 20895 20154
rect 20919 20102 20949 20154
rect 20949 20102 20961 20154
rect 20961 20102 20975 20154
rect 20999 20102 21013 20154
rect 21013 20102 21025 20154
rect 21025 20102 21055 20154
rect 21079 20102 21089 20154
rect 21089 20102 21135 20154
rect 20839 20100 20895 20102
rect 20919 20100 20975 20102
rect 20999 20100 21055 20102
rect 21079 20100 21135 20102
rect 20839 19066 20895 19068
rect 20919 19066 20975 19068
rect 20999 19066 21055 19068
rect 21079 19066 21135 19068
rect 20839 19014 20885 19066
rect 20885 19014 20895 19066
rect 20919 19014 20949 19066
rect 20949 19014 20961 19066
rect 20961 19014 20975 19066
rect 20999 19014 21013 19066
rect 21013 19014 21025 19066
rect 21025 19014 21055 19066
rect 21079 19014 21089 19066
rect 21089 19014 21135 19066
rect 20839 19012 20895 19014
rect 20919 19012 20975 19014
rect 20999 19012 21055 19014
rect 21079 19012 21135 19014
rect 20839 17978 20895 17980
rect 20919 17978 20975 17980
rect 20999 17978 21055 17980
rect 21079 17978 21135 17980
rect 20839 17926 20885 17978
rect 20885 17926 20895 17978
rect 20919 17926 20949 17978
rect 20949 17926 20961 17978
rect 20961 17926 20975 17978
rect 20999 17926 21013 17978
rect 21013 17926 21025 17978
rect 21025 17926 21055 17978
rect 21079 17926 21089 17978
rect 21089 17926 21135 17978
rect 20839 17924 20895 17926
rect 20919 17924 20975 17926
rect 20999 17924 21055 17926
rect 21079 17924 21135 17926
rect 23679 19610 23735 19612
rect 23759 19610 23815 19612
rect 23839 19610 23895 19612
rect 23919 19610 23975 19612
rect 23679 19558 23725 19610
rect 23725 19558 23735 19610
rect 23759 19558 23789 19610
rect 23789 19558 23801 19610
rect 23801 19558 23815 19610
rect 23839 19558 23853 19610
rect 23853 19558 23865 19610
rect 23865 19558 23895 19610
rect 23919 19558 23929 19610
rect 23929 19558 23975 19610
rect 23679 19556 23735 19558
rect 23759 19556 23815 19558
rect 23839 19556 23895 19558
rect 23919 19556 23975 19558
rect 23679 18522 23735 18524
rect 23759 18522 23815 18524
rect 23839 18522 23895 18524
rect 23919 18522 23975 18524
rect 23679 18470 23725 18522
rect 23725 18470 23735 18522
rect 23759 18470 23789 18522
rect 23789 18470 23801 18522
rect 23801 18470 23815 18522
rect 23839 18470 23853 18522
rect 23853 18470 23865 18522
rect 23865 18470 23895 18522
rect 23919 18470 23929 18522
rect 23929 18470 23975 18522
rect 23679 18468 23735 18470
rect 23759 18468 23815 18470
rect 23839 18468 23895 18470
rect 23919 18468 23975 18470
rect 20839 16890 20895 16892
rect 20919 16890 20975 16892
rect 20999 16890 21055 16892
rect 21079 16890 21135 16892
rect 20839 16838 20885 16890
rect 20885 16838 20895 16890
rect 20919 16838 20949 16890
rect 20949 16838 20961 16890
rect 20961 16838 20975 16890
rect 20999 16838 21013 16890
rect 21013 16838 21025 16890
rect 21025 16838 21055 16890
rect 21079 16838 21089 16890
rect 21089 16838 21135 16890
rect 20839 16836 20895 16838
rect 20919 16836 20975 16838
rect 20999 16836 21055 16838
rect 21079 16836 21135 16838
rect 20442 10512 20498 10568
rect 20839 15802 20895 15804
rect 20919 15802 20975 15804
rect 20999 15802 21055 15804
rect 21079 15802 21135 15804
rect 20839 15750 20885 15802
rect 20885 15750 20895 15802
rect 20919 15750 20949 15802
rect 20949 15750 20961 15802
rect 20961 15750 20975 15802
rect 20999 15750 21013 15802
rect 21013 15750 21025 15802
rect 21025 15750 21055 15802
rect 21079 15750 21089 15802
rect 21089 15750 21135 15802
rect 20839 15748 20895 15750
rect 20919 15748 20975 15750
rect 20999 15748 21055 15750
rect 21079 15748 21135 15750
rect 20839 14714 20895 14716
rect 20919 14714 20975 14716
rect 20999 14714 21055 14716
rect 21079 14714 21135 14716
rect 20839 14662 20885 14714
rect 20885 14662 20895 14714
rect 20919 14662 20949 14714
rect 20949 14662 20961 14714
rect 20961 14662 20975 14714
rect 20999 14662 21013 14714
rect 21013 14662 21025 14714
rect 21025 14662 21055 14714
rect 21079 14662 21089 14714
rect 21089 14662 21135 14714
rect 20839 14660 20895 14662
rect 20919 14660 20975 14662
rect 20999 14660 21055 14662
rect 21079 14660 21135 14662
rect 20839 13626 20895 13628
rect 20919 13626 20975 13628
rect 20999 13626 21055 13628
rect 21079 13626 21135 13628
rect 20839 13574 20885 13626
rect 20885 13574 20895 13626
rect 20919 13574 20949 13626
rect 20949 13574 20961 13626
rect 20961 13574 20975 13626
rect 20999 13574 21013 13626
rect 21013 13574 21025 13626
rect 21025 13574 21055 13626
rect 21079 13574 21089 13626
rect 21089 13574 21135 13626
rect 20839 13572 20895 13574
rect 20919 13572 20975 13574
rect 20999 13572 21055 13574
rect 21079 13572 21135 13574
rect 20839 12538 20895 12540
rect 20919 12538 20975 12540
rect 20999 12538 21055 12540
rect 21079 12538 21135 12540
rect 20839 12486 20885 12538
rect 20885 12486 20895 12538
rect 20919 12486 20949 12538
rect 20949 12486 20961 12538
rect 20961 12486 20975 12538
rect 20999 12486 21013 12538
rect 21013 12486 21025 12538
rect 21025 12486 21055 12538
rect 21079 12486 21089 12538
rect 21089 12486 21135 12538
rect 20839 12484 20895 12486
rect 20919 12484 20975 12486
rect 20999 12484 21055 12486
rect 21079 12484 21135 12486
rect 21086 12300 21142 12336
rect 21086 12280 21088 12300
rect 21088 12280 21140 12300
rect 21140 12280 21142 12300
rect 20839 11450 20895 11452
rect 20919 11450 20975 11452
rect 20999 11450 21055 11452
rect 21079 11450 21135 11452
rect 20839 11398 20885 11450
rect 20885 11398 20895 11450
rect 20919 11398 20949 11450
rect 20949 11398 20961 11450
rect 20961 11398 20975 11450
rect 20999 11398 21013 11450
rect 21013 11398 21025 11450
rect 21025 11398 21055 11450
rect 21079 11398 21089 11450
rect 21089 11398 21135 11450
rect 20839 11396 20895 11398
rect 20919 11396 20975 11398
rect 20999 11396 21055 11398
rect 21079 11396 21135 11398
rect 20839 10362 20895 10364
rect 20919 10362 20975 10364
rect 20999 10362 21055 10364
rect 21079 10362 21135 10364
rect 20839 10310 20885 10362
rect 20885 10310 20895 10362
rect 20919 10310 20949 10362
rect 20949 10310 20961 10362
rect 20961 10310 20975 10362
rect 20999 10310 21013 10362
rect 21013 10310 21025 10362
rect 21025 10310 21055 10362
rect 21079 10310 21089 10362
rect 21089 10310 21135 10362
rect 20839 10308 20895 10310
rect 20919 10308 20975 10310
rect 20999 10308 21055 10310
rect 21079 10308 21135 10310
rect 20839 9274 20895 9276
rect 20919 9274 20975 9276
rect 20999 9274 21055 9276
rect 21079 9274 21135 9276
rect 20839 9222 20885 9274
rect 20885 9222 20895 9274
rect 20919 9222 20949 9274
rect 20949 9222 20961 9274
rect 20961 9222 20975 9274
rect 20999 9222 21013 9274
rect 21013 9222 21025 9274
rect 21025 9222 21055 9274
rect 21079 9222 21089 9274
rect 21089 9222 21135 9274
rect 20839 9220 20895 9222
rect 20919 9220 20975 9222
rect 20999 9220 21055 9222
rect 21079 9220 21135 9222
rect 19246 5208 19302 5264
rect 18326 3440 18382 3496
rect 17998 3290 18054 3292
rect 18078 3290 18134 3292
rect 18158 3290 18214 3292
rect 18238 3290 18294 3292
rect 17998 3238 18044 3290
rect 18044 3238 18054 3290
rect 18078 3238 18108 3290
rect 18108 3238 18120 3290
rect 18120 3238 18134 3290
rect 18158 3238 18172 3290
rect 18172 3238 18184 3290
rect 18184 3238 18214 3290
rect 18238 3238 18248 3290
rect 18248 3238 18294 3290
rect 17998 3236 18054 3238
rect 18078 3236 18134 3238
rect 18158 3236 18214 3238
rect 18238 3236 18294 3238
rect 23679 17434 23735 17436
rect 23759 17434 23815 17436
rect 23839 17434 23895 17436
rect 23919 17434 23975 17436
rect 23679 17382 23725 17434
rect 23725 17382 23735 17434
rect 23759 17382 23789 17434
rect 23789 17382 23801 17434
rect 23801 17382 23815 17434
rect 23839 17382 23853 17434
rect 23853 17382 23865 17434
rect 23865 17382 23895 17434
rect 23919 17382 23929 17434
rect 23929 17382 23975 17434
rect 23679 17380 23735 17382
rect 23759 17380 23815 17382
rect 23839 17380 23895 17382
rect 23919 17380 23975 17382
rect 23679 16346 23735 16348
rect 23759 16346 23815 16348
rect 23839 16346 23895 16348
rect 23919 16346 23975 16348
rect 23679 16294 23725 16346
rect 23725 16294 23735 16346
rect 23759 16294 23789 16346
rect 23789 16294 23801 16346
rect 23801 16294 23815 16346
rect 23839 16294 23853 16346
rect 23853 16294 23865 16346
rect 23865 16294 23895 16346
rect 23919 16294 23929 16346
rect 23929 16294 23975 16346
rect 23679 16292 23735 16294
rect 23759 16292 23815 16294
rect 23839 16292 23895 16294
rect 23919 16292 23975 16294
rect 20839 8186 20895 8188
rect 20919 8186 20975 8188
rect 20999 8186 21055 8188
rect 21079 8186 21135 8188
rect 20839 8134 20885 8186
rect 20885 8134 20895 8186
rect 20919 8134 20949 8186
rect 20949 8134 20961 8186
rect 20961 8134 20975 8186
rect 20999 8134 21013 8186
rect 21013 8134 21025 8186
rect 21025 8134 21055 8186
rect 21079 8134 21089 8186
rect 21089 8134 21135 8186
rect 20839 8132 20895 8134
rect 20919 8132 20975 8134
rect 20999 8132 21055 8134
rect 21079 8132 21135 8134
rect 20839 7098 20895 7100
rect 20919 7098 20975 7100
rect 20999 7098 21055 7100
rect 21079 7098 21135 7100
rect 20839 7046 20885 7098
rect 20885 7046 20895 7098
rect 20919 7046 20949 7098
rect 20949 7046 20961 7098
rect 20961 7046 20975 7098
rect 20999 7046 21013 7098
rect 21013 7046 21025 7098
rect 21025 7046 21055 7098
rect 21079 7046 21089 7098
rect 21089 7046 21135 7098
rect 20839 7044 20895 7046
rect 20919 7044 20975 7046
rect 20999 7044 21055 7046
rect 21079 7044 21135 7046
rect 20839 6010 20895 6012
rect 20919 6010 20975 6012
rect 20999 6010 21055 6012
rect 21079 6010 21135 6012
rect 20839 5958 20885 6010
rect 20885 5958 20895 6010
rect 20919 5958 20949 6010
rect 20949 5958 20961 6010
rect 20961 5958 20975 6010
rect 20999 5958 21013 6010
rect 21013 5958 21025 6010
rect 21025 5958 21055 6010
rect 21079 5958 21089 6010
rect 21089 5958 21135 6010
rect 20839 5956 20895 5958
rect 20919 5956 20975 5958
rect 20999 5956 21055 5958
rect 21079 5956 21135 5958
rect 21178 5616 21234 5672
rect 20839 4922 20895 4924
rect 20919 4922 20975 4924
rect 20999 4922 21055 4924
rect 21079 4922 21135 4924
rect 20839 4870 20885 4922
rect 20885 4870 20895 4922
rect 20919 4870 20949 4922
rect 20949 4870 20961 4922
rect 20961 4870 20975 4922
rect 20999 4870 21013 4922
rect 21013 4870 21025 4922
rect 21025 4870 21055 4922
rect 21079 4870 21089 4922
rect 21089 4870 21135 4922
rect 20839 4868 20895 4870
rect 20919 4868 20975 4870
rect 20999 4868 21055 4870
rect 21079 4868 21135 4870
rect 22742 13368 22798 13424
rect 23679 15258 23735 15260
rect 23759 15258 23815 15260
rect 23839 15258 23895 15260
rect 23919 15258 23975 15260
rect 23679 15206 23725 15258
rect 23725 15206 23735 15258
rect 23759 15206 23789 15258
rect 23789 15206 23801 15258
rect 23801 15206 23815 15258
rect 23839 15206 23853 15258
rect 23853 15206 23865 15258
rect 23865 15206 23895 15258
rect 23919 15206 23929 15258
rect 23929 15206 23975 15258
rect 23679 15204 23735 15206
rect 23759 15204 23815 15206
rect 23839 15204 23895 15206
rect 23919 15204 23975 15206
rect 22006 8336 22062 8392
rect 22190 6860 22246 6896
rect 22190 6840 22192 6860
rect 22192 6840 22244 6860
rect 22244 6840 22246 6860
rect 23679 14170 23735 14172
rect 23759 14170 23815 14172
rect 23839 14170 23895 14172
rect 23919 14170 23975 14172
rect 23679 14118 23725 14170
rect 23725 14118 23735 14170
rect 23759 14118 23789 14170
rect 23789 14118 23801 14170
rect 23801 14118 23815 14170
rect 23839 14118 23853 14170
rect 23853 14118 23865 14170
rect 23865 14118 23895 14170
rect 23919 14118 23929 14170
rect 23929 14118 23975 14170
rect 23679 14116 23735 14118
rect 23759 14116 23815 14118
rect 23839 14116 23895 14118
rect 23919 14116 23975 14118
rect 23679 13082 23735 13084
rect 23759 13082 23815 13084
rect 23839 13082 23895 13084
rect 23919 13082 23975 13084
rect 23679 13030 23725 13082
rect 23725 13030 23735 13082
rect 23759 13030 23789 13082
rect 23789 13030 23801 13082
rect 23801 13030 23815 13082
rect 23839 13030 23853 13082
rect 23853 13030 23865 13082
rect 23865 13030 23895 13082
rect 23919 13030 23929 13082
rect 23929 13030 23975 13082
rect 23679 13028 23735 13030
rect 23759 13028 23815 13030
rect 23839 13028 23895 13030
rect 23919 13028 23975 13030
rect 23679 11994 23735 11996
rect 23759 11994 23815 11996
rect 23839 11994 23895 11996
rect 23919 11994 23975 11996
rect 23679 11942 23725 11994
rect 23725 11942 23735 11994
rect 23759 11942 23789 11994
rect 23789 11942 23801 11994
rect 23801 11942 23815 11994
rect 23839 11942 23853 11994
rect 23853 11942 23865 11994
rect 23865 11942 23895 11994
rect 23919 11942 23929 11994
rect 23929 11942 23975 11994
rect 23679 11940 23735 11942
rect 23759 11940 23815 11942
rect 23839 11940 23895 11942
rect 23919 11940 23975 11942
rect 23679 10906 23735 10908
rect 23759 10906 23815 10908
rect 23839 10906 23895 10908
rect 23919 10906 23975 10908
rect 23679 10854 23725 10906
rect 23725 10854 23735 10906
rect 23759 10854 23789 10906
rect 23789 10854 23801 10906
rect 23801 10854 23815 10906
rect 23839 10854 23853 10906
rect 23853 10854 23865 10906
rect 23865 10854 23895 10906
rect 23919 10854 23929 10906
rect 23929 10854 23975 10906
rect 23679 10852 23735 10854
rect 23759 10852 23815 10854
rect 23839 10852 23895 10854
rect 23919 10852 23975 10854
rect 23679 9818 23735 9820
rect 23759 9818 23815 9820
rect 23839 9818 23895 9820
rect 23919 9818 23975 9820
rect 23679 9766 23725 9818
rect 23725 9766 23735 9818
rect 23759 9766 23789 9818
rect 23789 9766 23801 9818
rect 23801 9766 23815 9818
rect 23839 9766 23853 9818
rect 23853 9766 23865 9818
rect 23865 9766 23895 9818
rect 23919 9766 23929 9818
rect 23929 9766 23975 9818
rect 23679 9764 23735 9766
rect 23759 9764 23815 9766
rect 23839 9764 23895 9766
rect 23919 9764 23975 9766
rect 23679 8730 23735 8732
rect 23759 8730 23815 8732
rect 23839 8730 23895 8732
rect 23919 8730 23975 8732
rect 23679 8678 23725 8730
rect 23725 8678 23735 8730
rect 23759 8678 23789 8730
rect 23789 8678 23801 8730
rect 23801 8678 23815 8730
rect 23839 8678 23853 8730
rect 23853 8678 23865 8730
rect 23865 8678 23895 8730
rect 23919 8678 23929 8730
rect 23929 8678 23975 8730
rect 23679 8676 23735 8678
rect 23759 8676 23815 8678
rect 23839 8676 23895 8678
rect 23919 8676 23975 8678
rect 23679 7642 23735 7644
rect 23759 7642 23815 7644
rect 23839 7642 23895 7644
rect 23919 7642 23975 7644
rect 23679 7590 23725 7642
rect 23725 7590 23735 7642
rect 23759 7590 23789 7642
rect 23789 7590 23801 7642
rect 23801 7590 23815 7642
rect 23839 7590 23853 7642
rect 23853 7590 23865 7642
rect 23865 7590 23895 7642
rect 23919 7590 23929 7642
rect 23929 7590 23975 7642
rect 23679 7588 23735 7590
rect 23759 7588 23815 7590
rect 23839 7588 23895 7590
rect 23919 7588 23975 7590
rect 23679 6554 23735 6556
rect 23759 6554 23815 6556
rect 23839 6554 23895 6556
rect 23919 6554 23975 6556
rect 23679 6502 23725 6554
rect 23725 6502 23735 6554
rect 23759 6502 23789 6554
rect 23789 6502 23801 6554
rect 23801 6502 23815 6554
rect 23839 6502 23853 6554
rect 23853 6502 23865 6554
rect 23865 6502 23895 6554
rect 23919 6502 23929 6554
rect 23929 6502 23975 6554
rect 23679 6500 23735 6502
rect 23759 6500 23815 6502
rect 23839 6500 23895 6502
rect 23919 6500 23975 6502
rect 23294 5616 23350 5672
rect 23679 5466 23735 5468
rect 23759 5466 23815 5468
rect 23839 5466 23895 5468
rect 23919 5466 23975 5468
rect 23679 5414 23725 5466
rect 23725 5414 23735 5466
rect 23759 5414 23789 5466
rect 23789 5414 23801 5466
rect 23801 5414 23815 5466
rect 23839 5414 23853 5466
rect 23853 5414 23865 5466
rect 23865 5414 23895 5466
rect 23919 5414 23929 5466
rect 23929 5414 23975 5466
rect 23679 5412 23735 5414
rect 23759 5412 23815 5414
rect 23839 5412 23895 5414
rect 23919 5412 23975 5414
rect 23679 4378 23735 4380
rect 23759 4378 23815 4380
rect 23839 4378 23895 4380
rect 23919 4378 23975 4380
rect 23679 4326 23725 4378
rect 23725 4326 23735 4378
rect 23759 4326 23789 4378
rect 23789 4326 23801 4378
rect 23801 4326 23815 4378
rect 23839 4326 23853 4378
rect 23853 4326 23865 4378
rect 23865 4326 23895 4378
rect 23919 4326 23929 4378
rect 23929 4326 23975 4378
rect 23679 4324 23735 4326
rect 23759 4324 23815 4326
rect 23839 4324 23895 4326
rect 23919 4324 23975 4326
rect 20839 3834 20895 3836
rect 20919 3834 20975 3836
rect 20999 3834 21055 3836
rect 21079 3834 21135 3836
rect 20839 3782 20885 3834
rect 20885 3782 20895 3834
rect 20919 3782 20949 3834
rect 20949 3782 20961 3834
rect 20961 3782 20975 3834
rect 20999 3782 21013 3834
rect 21013 3782 21025 3834
rect 21025 3782 21055 3834
rect 21079 3782 21089 3834
rect 21089 3782 21135 3834
rect 20839 3780 20895 3782
rect 20919 3780 20975 3782
rect 20999 3780 21055 3782
rect 21079 3780 21135 3782
rect 17998 2202 18054 2204
rect 18078 2202 18134 2204
rect 18158 2202 18214 2204
rect 18238 2202 18294 2204
rect 17998 2150 18044 2202
rect 18044 2150 18054 2202
rect 18078 2150 18108 2202
rect 18108 2150 18120 2202
rect 18120 2150 18134 2202
rect 18158 2150 18172 2202
rect 18172 2150 18184 2202
rect 18184 2150 18214 2202
rect 18238 2150 18248 2202
rect 18248 2150 18294 2202
rect 17998 2148 18054 2150
rect 18078 2148 18134 2150
rect 18158 2148 18214 2150
rect 18238 2148 18294 2150
rect 20839 2746 20895 2748
rect 20919 2746 20975 2748
rect 20999 2746 21055 2748
rect 21079 2746 21135 2748
rect 20839 2694 20885 2746
rect 20885 2694 20895 2746
rect 20919 2694 20949 2746
rect 20949 2694 20961 2746
rect 20961 2694 20975 2746
rect 20999 2694 21013 2746
rect 21013 2694 21025 2746
rect 21025 2694 21055 2746
rect 21079 2694 21089 2746
rect 21089 2694 21135 2746
rect 20839 2692 20895 2694
rect 20919 2692 20975 2694
rect 20999 2692 21055 2694
rect 21079 2692 21135 2694
rect 23679 3290 23735 3292
rect 23759 3290 23815 3292
rect 23839 3290 23895 3292
rect 23919 3290 23975 3292
rect 23679 3238 23725 3290
rect 23725 3238 23735 3290
rect 23759 3238 23789 3290
rect 23789 3238 23801 3290
rect 23801 3238 23815 3290
rect 23839 3238 23853 3290
rect 23853 3238 23865 3290
rect 23865 3238 23895 3290
rect 23919 3238 23929 3290
rect 23929 3238 23975 3290
rect 23679 3236 23735 3238
rect 23759 3236 23815 3238
rect 23839 3236 23895 3238
rect 23919 3236 23975 3238
rect 23679 2202 23735 2204
rect 23759 2202 23815 2204
rect 23839 2202 23895 2204
rect 23919 2202 23975 2204
rect 23679 2150 23725 2202
rect 23725 2150 23735 2202
rect 23759 2150 23789 2202
rect 23789 2150 23801 2202
rect 23801 2150 23815 2202
rect 23839 2150 23853 2202
rect 23853 2150 23865 2202
rect 23865 2150 23895 2202
rect 23919 2150 23929 2202
rect 23929 2150 23975 2202
rect 23679 2148 23735 2150
rect 23759 2148 23815 2150
rect 23839 2148 23895 2150
rect 23919 2148 23975 2150
<< metal3 >>
rect 3786 22336 4102 22337
rect 3786 22272 3792 22336
rect 3856 22272 3872 22336
rect 3936 22272 3952 22336
rect 4016 22272 4032 22336
rect 4096 22272 4102 22336
rect 3786 22271 4102 22272
rect 9467 22336 9783 22337
rect 9467 22272 9473 22336
rect 9537 22272 9553 22336
rect 9617 22272 9633 22336
rect 9697 22272 9713 22336
rect 9777 22272 9783 22336
rect 9467 22271 9783 22272
rect 15148 22336 15464 22337
rect 15148 22272 15154 22336
rect 15218 22272 15234 22336
rect 15298 22272 15314 22336
rect 15378 22272 15394 22336
rect 15458 22272 15464 22336
rect 15148 22271 15464 22272
rect 20829 22336 21145 22337
rect 20829 22272 20835 22336
rect 20899 22272 20915 22336
rect 20979 22272 20995 22336
rect 21059 22272 21075 22336
rect 21139 22272 21145 22336
rect 20829 22271 21145 22272
rect 13169 21994 13235 21997
rect 20437 21994 20503 21997
rect 13169 21992 20503 21994
rect 13169 21936 13174 21992
rect 13230 21936 20442 21992
rect 20498 21936 20503 21992
rect 13169 21934 20503 21936
rect 13169 21931 13235 21934
rect 20437 21931 20503 21934
rect 6626 21792 6942 21793
rect 6626 21728 6632 21792
rect 6696 21728 6712 21792
rect 6776 21728 6792 21792
rect 6856 21728 6872 21792
rect 6936 21728 6942 21792
rect 6626 21727 6942 21728
rect 12307 21792 12623 21793
rect 12307 21728 12313 21792
rect 12377 21728 12393 21792
rect 12457 21728 12473 21792
rect 12537 21728 12553 21792
rect 12617 21728 12623 21792
rect 12307 21727 12623 21728
rect 17988 21792 18304 21793
rect 17988 21728 17994 21792
rect 18058 21728 18074 21792
rect 18138 21728 18154 21792
rect 18218 21728 18234 21792
rect 18298 21728 18304 21792
rect 17988 21727 18304 21728
rect 23669 21792 23985 21793
rect 23669 21728 23675 21792
rect 23739 21728 23755 21792
rect 23819 21728 23835 21792
rect 23899 21728 23915 21792
rect 23979 21728 23985 21792
rect 23669 21727 23985 21728
rect 12525 21450 12591 21453
rect 19517 21450 19583 21453
rect 12525 21448 19583 21450
rect 12525 21392 12530 21448
rect 12586 21392 19522 21448
rect 19578 21392 19583 21448
rect 12525 21390 19583 21392
rect 12525 21387 12591 21390
rect 19517 21387 19583 21390
rect 14181 21316 14247 21317
rect 14181 21314 14228 21316
rect 14136 21312 14228 21314
rect 14136 21256 14186 21312
rect 14136 21254 14228 21256
rect 14181 21252 14228 21254
rect 14292 21252 14298 21316
rect 14181 21251 14247 21252
rect 3786 21248 4102 21249
rect 3786 21184 3792 21248
rect 3856 21184 3872 21248
rect 3936 21184 3952 21248
rect 4016 21184 4032 21248
rect 4096 21184 4102 21248
rect 3786 21183 4102 21184
rect 9467 21248 9783 21249
rect 9467 21184 9473 21248
rect 9537 21184 9553 21248
rect 9617 21184 9633 21248
rect 9697 21184 9713 21248
rect 9777 21184 9783 21248
rect 9467 21183 9783 21184
rect 15148 21248 15464 21249
rect 15148 21184 15154 21248
rect 15218 21184 15234 21248
rect 15298 21184 15314 21248
rect 15378 21184 15394 21248
rect 15458 21184 15464 21248
rect 15148 21183 15464 21184
rect 20829 21248 21145 21249
rect 20829 21184 20835 21248
rect 20899 21184 20915 21248
rect 20979 21184 20995 21248
rect 21059 21184 21075 21248
rect 21139 21184 21145 21248
rect 20829 21183 21145 21184
rect 10961 20906 11027 20909
rect 21909 20906 21975 20909
rect 10961 20904 21975 20906
rect 10961 20848 10966 20904
rect 11022 20848 21914 20904
rect 21970 20848 21975 20904
rect 10961 20846 21975 20848
rect 10961 20843 11027 20846
rect 21909 20843 21975 20846
rect 4613 20772 4679 20773
rect 4613 20768 4660 20772
rect 4724 20770 4730 20772
rect 19609 20770 19675 20773
rect 19742 20770 19748 20772
rect 4613 20712 4618 20768
rect 4613 20708 4660 20712
rect 4724 20710 4770 20770
rect 19609 20768 19748 20770
rect 19609 20712 19614 20768
rect 19670 20712 19748 20768
rect 19609 20710 19748 20712
rect 4724 20708 4730 20710
rect 4613 20707 4679 20708
rect 19609 20707 19675 20710
rect 19742 20708 19748 20710
rect 19812 20708 19818 20772
rect 6626 20704 6942 20705
rect 6626 20640 6632 20704
rect 6696 20640 6712 20704
rect 6776 20640 6792 20704
rect 6856 20640 6872 20704
rect 6936 20640 6942 20704
rect 6626 20639 6942 20640
rect 12307 20704 12623 20705
rect 12307 20640 12313 20704
rect 12377 20640 12393 20704
rect 12457 20640 12473 20704
rect 12537 20640 12553 20704
rect 12617 20640 12623 20704
rect 12307 20639 12623 20640
rect 17988 20704 18304 20705
rect 17988 20640 17994 20704
rect 18058 20640 18074 20704
rect 18138 20640 18154 20704
rect 18218 20640 18234 20704
rect 18298 20640 18304 20704
rect 17988 20639 18304 20640
rect 23669 20704 23985 20705
rect 23669 20640 23675 20704
rect 23739 20640 23755 20704
rect 23819 20640 23835 20704
rect 23899 20640 23915 20704
rect 23979 20640 23985 20704
rect 23669 20639 23985 20640
rect 3786 20160 4102 20161
rect 3786 20096 3792 20160
rect 3856 20096 3872 20160
rect 3936 20096 3952 20160
rect 4016 20096 4032 20160
rect 4096 20096 4102 20160
rect 3786 20095 4102 20096
rect 9467 20160 9783 20161
rect 9467 20096 9473 20160
rect 9537 20096 9553 20160
rect 9617 20096 9633 20160
rect 9697 20096 9713 20160
rect 9777 20096 9783 20160
rect 9467 20095 9783 20096
rect 15148 20160 15464 20161
rect 15148 20096 15154 20160
rect 15218 20096 15234 20160
rect 15298 20096 15314 20160
rect 15378 20096 15394 20160
rect 15458 20096 15464 20160
rect 15148 20095 15464 20096
rect 20829 20160 21145 20161
rect 20829 20096 20835 20160
rect 20899 20096 20915 20160
rect 20979 20096 20995 20160
rect 21059 20096 21075 20160
rect 21139 20096 21145 20160
rect 20829 20095 21145 20096
rect 6626 19616 6942 19617
rect 6626 19552 6632 19616
rect 6696 19552 6712 19616
rect 6776 19552 6792 19616
rect 6856 19552 6872 19616
rect 6936 19552 6942 19616
rect 6626 19551 6942 19552
rect 12307 19616 12623 19617
rect 12307 19552 12313 19616
rect 12377 19552 12393 19616
rect 12457 19552 12473 19616
rect 12537 19552 12553 19616
rect 12617 19552 12623 19616
rect 12307 19551 12623 19552
rect 17988 19616 18304 19617
rect 17988 19552 17994 19616
rect 18058 19552 18074 19616
rect 18138 19552 18154 19616
rect 18218 19552 18234 19616
rect 18298 19552 18304 19616
rect 17988 19551 18304 19552
rect 23669 19616 23985 19617
rect 23669 19552 23675 19616
rect 23739 19552 23755 19616
rect 23819 19552 23835 19616
rect 23899 19552 23915 19616
rect 23979 19552 23985 19616
rect 23669 19551 23985 19552
rect 5349 19412 5415 19413
rect 5349 19408 5396 19412
rect 5460 19410 5466 19412
rect 5349 19352 5354 19408
rect 5349 19348 5396 19352
rect 5460 19350 5506 19410
rect 5460 19348 5466 19350
rect 5349 19347 5415 19348
rect 13537 19274 13603 19277
rect 15837 19274 15903 19277
rect 13537 19272 15903 19274
rect 13537 19216 13542 19272
rect 13598 19216 15842 19272
rect 15898 19216 15903 19272
rect 13537 19214 15903 19216
rect 13537 19211 13603 19214
rect 15837 19211 15903 19214
rect 3786 19072 4102 19073
rect 3786 19008 3792 19072
rect 3856 19008 3872 19072
rect 3936 19008 3952 19072
rect 4016 19008 4032 19072
rect 4096 19008 4102 19072
rect 3786 19007 4102 19008
rect 9467 19072 9783 19073
rect 9467 19008 9473 19072
rect 9537 19008 9553 19072
rect 9617 19008 9633 19072
rect 9697 19008 9713 19072
rect 9777 19008 9783 19072
rect 9467 19007 9783 19008
rect 15148 19072 15464 19073
rect 15148 19008 15154 19072
rect 15218 19008 15234 19072
rect 15298 19008 15314 19072
rect 15378 19008 15394 19072
rect 15458 19008 15464 19072
rect 15148 19007 15464 19008
rect 20829 19072 21145 19073
rect 20829 19008 20835 19072
rect 20899 19008 20915 19072
rect 20979 19008 20995 19072
rect 21059 19008 21075 19072
rect 21139 19008 21145 19072
rect 20829 19007 21145 19008
rect 14733 18866 14799 18869
rect 14958 18866 14964 18868
rect 14733 18864 14964 18866
rect 14733 18808 14738 18864
rect 14794 18808 14964 18864
rect 14733 18806 14964 18808
rect 14733 18803 14799 18806
rect 14958 18804 14964 18806
rect 15028 18804 15034 18868
rect 6626 18528 6942 18529
rect 6626 18464 6632 18528
rect 6696 18464 6712 18528
rect 6776 18464 6792 18528
rect 6856 18464 6872 18528
rect 6936 18464 6942 18528
rect 6626 18463 6942 18464
rect 12307 18528 12623 18529
rect 12307 18464 12313 18528
rect 12377 18464 12393 18528
rect 12457 18464 12473 18528
rect 12537 18464 12553 18528
rect 12617 18464 12623 18528
rect 12307 18463 12623 18464
rect 17988 18528 18304 18529
rect 17988 18464 17994 18528
rect 18058 18464 18074 18528
rect 18138 18464 18154 18528
rect 18218 18464 18234 18528
rect 18298 18464 18304 18528
rect 17988 18463 18304 18464
rect 23669 18528 23985 18529
rect 23669 18464 23675 18528
rect 23739 18464 23755 18528
rect 23819 18464 23835 18528
rect 23899 18464 23915 18528
rect 23979 18464 23985 18528
rect 23669 18463 23985 18464
rect 15009 18186 15075 18189
rect 17677 18186 17743 18189
rect 15009 18184 17743 18186
rect 15009 18128 15014 18184
rect 15070 18128 17682 18184
rect 17738 18128 17743 18184
rect 15009 18126 17743 18128
rect 15009 18123 15075 18126
rect 17677 18123 17743 18126
rect 19885 18052 19951 18053
rect 19885 18048 19932 18052
rect 19996 18050 20002 18052
rect 19885 17992 19890 18048
rect 19885 17988 19932 17992
rect 19996 17990 20042 18050
rect 19996 17988 20002 17990
rect 19885 17987 19951 17988
rect 3786 17984 4102 17985
rect 3786 17920 3792 17984
rect 3856 17920 3872 17984
rect 3936 17920 3952 17984
rect 4016 17920 4032 17984
rect 4096 17920 4102 17984
rect 3786 17919 4102 17920
rect 9467 17984 9783 17985
rect 9467 17920 9473 17984
rect 9537 17920 9553 17984
rect 9617 17920 9633 17984
rect 9697 17920 9713 17984
rect 9777 17920 9783 17984
rect 9467 17919 9783 17920
rect 15148 17984 15464 17985
rect 15148 17920 15154 17984
rect 15218 17920 15234 17984
rect 15298 17920 15314 17984
rect 15378 17920 15394 17984
rect 15458 17920 15464 17984
rect 15148 17919 15464 17920
rect 20829 17984 21145 17985
rect 20829 17920 20835 17984
rect 20899 17920 20915 17984
rect 20979 17920 20995 17984
rect 21059 17920 21075 17984
rect 21139 17920 21145 17984
rect 20829 17919 21145 17920
rect 13353 17642 13419 17645
rect 15101 17642 15167 17645
rect 16481 17642 16547 17645
rect 13353 17640 16547 17642
rect 13353 17584 13358 17640
rect 13414 17584 15106 17640
rect 15162 17584 16486 17640
rect 16542 17584 16547 17640
rect 13353 17582 16547 17584
rect 13353 17579 13419 17582
rect 15101 17579 15167 17582
rect 16481 17579 16547 17582
rect 6626 17440 6942 17441
rect 6626 17376 6632 17440
rect 6696 17376 6712 17440
rect 6776 17376 6792 17440
rect 6856 17376 6872 17440
rect 6936 17376 6942 17440
rect 6626 17375 6942 17376
rect 12307 17440 12623 17441
rect 12307 17376 12313 17440
rect 12377 17376 12393 17440
rect 12457 17376 12473 17440
rect 12537 17376 12553 17440
rect 12617 17376 12623 17440
rect 12307 17375 12623 17376
rect 17988 17440 18304 17441
rect 17988 17376 17994 17440
rect 18058 17376 18074 17440
rect 18138 17376 18154 17440
rect 18218 17376 18234 17440
rect 18298 17376 18304 17440
rect 17988 17375 18304 17376
rect 23669 17440 23985 17441
rect 23669 17376 23675 17440
rect 23739 17376 23755 17440
rect 23819 17376 23835 17440
rect 23899 17376 23915 17440
rect 23979 17376 23985 17440
rect 23669 17375 23985 17376
rect 14457 17098 14523 17101
rect 18597 17098 18663 17101
rect 14457 17096 18663 17098
rect 14457 17040 14462 17096
rect 14518 17040 18602 17096
rect 18658 17040 18663 17096
rect 14457 17038 18663 17040
rect 14457 17035 14523 17038
rect 18597 17035 18663 17038
rect 3786 16896 4102 16897
rect 3786 16832 3792 16896
rect 3856 16832 3872 16896
rect 3936 16832 3952 16896
rect 4016 16832 4032 16896
rect 4096 16832 4102 16896
rect 3786 16831 4102 16832
rect 9467 16896 9783 16897
rect 9467 16832 9473 16896
rect 9537 16832 9553 16896
rect 9617 16832 9633 16896
rect 9697 16832 9713 16896
rect 9777 16832 9783 16896
rect 9467 16831 9783 16832
rect 15148 16896 15464 16897
rect 15148 16832 15154 16896
rect 15218 16832 15234 16896
rect 15298 16832 15314 16896
rect 15378 16832 15394 16896
rect 15458 16832 15464 16896
rect 15148 16831 15464 16832
rect 20829 16896 21145 16897
rect 20829 16832 20835 16896
rect 20899 16832 20915 16896
rect 20979 16832 20995 16896
rect 21059 16832 21075 16896
rect 21139 16832 21145 16896
rect 20829 16831 21145 16832
rect 6085 16690 6151 16693
rect 6310 16690 6316 16692
rect 6085 16688 6316 16690
rect 6085 16632 6090 16688
rect 6146 16632 6316 16688
rect 6085 16630 6316 16632
rect 6085 16627 6151 16630
rect 6310 16628 6316 16630
rect 6380 16628 6386 16692
rect 14825 16554 14891 16557
rect 19425 16554 19491 16557
rect 14825 16552 19491 16554
rect 14825 16496 14830 16552
rect 14886 16496 19430 16552
rect 19486 16496 19491 16552
rect 14825 16494 19491 16496
rect 14825 16491 14891 16494
rect 19425 16491 19491 16494
rect 6626 16352 6942 16353
rect 6626 16288 6632 16352
rect 6696 16288 6712 16352
rect 6776 16288 6792 16352
rect 6856 16288 6872 16352
rect 6936 16288 6942 16352
rect 6626 16287 6942 16288
rect 12307 16352 12623 16353
rect 12307 16288 12313 16352
rect 12377 16288 12393 16352
rect 12457 16288 12473 16352
rect 12537 16288 12553 16352
rect 12617 16288 12623 16352
rect 12307 16287 12623 16288
rect 17988 16352 18304 16353
rect 17988 16288 17994 16352
rect 18058 16288 18074 16352
rect 18138 16288 18154 16352
rect 18218 16288 18234 16352
rect 18298 16288 18304 16352
rect 17988 16287 18304 16288
rect 23669 16352 23985 16353
rect 23669 16288 23675 16352
rect 23739 16288 23755 16352
rect 23819 16288 23835 16352
rect 23899 16288 23915 16352
rect 23979 16288 23985 16352
rect 23669 16287 23985 16288
rect 15009 16010 15075 16013
rect 19057 16010 19123 16013
rect 15009 16008 19123 16010
rect 15009 15952 15014 16008
rect 15070 15952 19062 16008
rect 19118 15952 19123 16008
rect 15009 15950 19123 15952
rect 15009 15947 15075 15950
rect 19057 15947 19123 15950
rect 3786 15808 4102 15809
rect 3786 15744 3792 15808
rect 3856 15744 3872 15808
rect 3936 15744 3952 15808
rect 4016 15744 4032 15808
rect 4096 15744 4102 15808
rect 3786 15743 4102 15744
rect 9467 15808 9783 15809
rect 9467 15744 9473 15808
rect 9537 15744 9553 15808
rect 9617 15744 9633 15808
rect 9697 15744 9713 15808
rect 9777 15744 9783 15808
rect 9467 15743 9783 15744
rect 15148 15808 15464 15809
rect 15148 15744 15154 15808
rect 15218 15744 15234 15808
rect 15298 15744 15314 15808
rect 15378 15744 15394 15808
rect 15458 15744 15464 15808
rect 15148 15743 15464 15744
rect 20829 15808 21145 15809
rect 20829 15744 20835 15808
rect 20899 15744 20915 15808
rect 20979 15744 20995 15808
rect 21059 15744 21075 15808
rect 21139 15744 21145 15808
rect 20829 15743 21145 15744
rect 6626 15264 6942 15265
rect 6626 15200 6632 15264
rect 6696 15200 6712 15264
rect 6776 15200 6792 15264
rect 6856 15200 6872 15264
rect 6936 15200 6942 15264
rect 6626 15199 6942 15200
rect 12307 15264 12623 15265
rect 12307 15200 12313 15264
rect 12377 15200 12393 15264
rect 12457 15200 12473 15264
rect 12537 15200 12553 15264
rect 12617 15200 12623 15264
rect 12307 15199 12623 15200
rect 17988 15264 18304 15265
rect 17988 15200 17994 15264
rect 18058 15200 18074 15264
rect 18138 15200 18154 15264
rect 18218 15200 18234 15264
rect 18298 15200 18304 15264
rect 17988 15199 18304 15200
rect 23669 15264 23985 15265
rect 23669 15200 23675 15264
rect 23739 15200 23755 15264
rect 23819 15200 23835 15264
rect 23899 15200 23915 15264
rect 23979 15200 23985 15264
rect 23669 15199 23985 15200
rect 14222 15132 14228 15196
rect 14292 15194 14298 15196
rect 16665 15194 16731 15197
rect 14292 15192 16731 15194
rect 14292 15136 16670 15192
rect 16726 15136 16731 15192
rect 14292 15134 16731 15136
rect 14292 15132 14298 15134
rect 16665 15131 16731 15134
rect 3786 14720 4102 14721
rect 3786 14656 3792 14720
rect 3856 14656 3872 14720
rect 3936 14656 3952 14720
rect 4016 14656 4032 14720
rect 4096 14656 4102 14720
rect 3786 14655 4102 14656
rect 9467 14720 9783 14721
rect 9467 14656 9473 14720
rect 9537 14656 9553 14720
rect 9617 14656 9633 14720
rect 9697 14656 9713 14720
rect 9777 14656 9783 14720
rect 9467 14655 9783 14656
rect 15148 14720 15464 14721
rect 15148 14656 15154 14720
rect 15218 14656 15234 14720
rect 15298 14656 15314 14720
rect 15378 14656 15394 14720
rect 15458 14656 15464 14720
rect 15148 14655 15464 14656
rect 20829 14720 21145 14721
rect 20829 14656 20835 14720
rect 20899 14656 20915 14720
rect 20979 14656 20995 14720
rect 21059 14656 21075 14720
rect 21139 14656 21145 14720
rect 20829 14655 21145 14656
rect 6626 14176 6942 14177
rect 6626 14112 6632 14176
rect 6696 14112 6712 14176
rect 6776 14112 6792 14176
rect 6856 14112 6872 14176
rect 6936 14112 6942 14176
rect 6626 14111 6942 14112
rect 12307 14176 12623 14177
rect 12307 14112 12313 14176
rect 12377 14112 12393 14176
rect 12457 14112 12473 14176
rect 12537 14112 12553 14176
rect 12617 14112 12623 14176
rect 12307 14111 12623 14112
rect 17988 14176 18304 14177
rect 17988 14112 17994 14176
rect 18058 14112 18074 14176
rect 18138 14112 18154 14176
rect 18218 14112 18234 14176
rect 18298 14112 18304 14176
rect 17988 14111 18304 14112
rect 23669 14176 23985 14177
rect 23669 14112 23675 14176
rect 23739 14112 23755 14176
rect 23819 14112 23835 14176
rect 23899 14112 23915 14176
rect 23979 14112 23985 14176
rect 23669 14111 23985 14112
rect 14457 13834 14523 13837
rect 14590 13834 14596 13836
rect 14457 13832 14596 13834
rect 14457 13776 14462 13832
rect 14518 13776 14596 13832
rect 14457 13774 14596 13776
rect 14457 13771 14523 13774
rect 14590 13772 14596 13774
rect 14660 13772 14666 13836
rect 14958 13772 14964 13836
rect 15028 13834 15034 13836
rect 16849 13834 16915 13837
rect 15028 13832 16915 13834
rect 15028 13776 16854 13832
rect 16910 13776 16915 13832
rect 15028 13774 16915 13776
rect 15028 13772 15034 13774
rect 16849 13771 16915 13774
rect 3786 13632 4102 13633
rect 3786 13568 3792 13632
rect 3856 13568 3872 13632
rect 3936 13568 3952 13632
rect 4016 13568 4032 13632
rect 4096 13568 4102 13632
rect 3786 13567 4102 13568
rect 9467 13632 9783 13633
rect 9467 13568 9473 13632
rect 9537 13568 9553 13632
rect 9617 13568 9633 13632
rect 9697 13568 9713 13632
rect 9777 13568 9783 13632
rect 9467 13567 9783 13568
rect 15148 13632 15464 13633
rect 15148 13568 15154 13632
rect 15218 13568 15234 13632
rect 15298 13568 15314 13632
rect 15378 13568 15394 13632
rect 15458 13568 15464 13632
rect 15148 13567 15464 13568
rect 20829 13632 21145 13633
rect 20829 13568 20835 13632
rect 20899 13568 20915 13632
rect 20979 13568 20995 13632
rect 21059 13568 21075 13632
rect 21139 13568 21145 13632
rect 20829 13567 21145 13568
rect 13353 13426 13419 13429
rect 22737 13426 22803 13429
rect 13353 13424 22803 13426
rect 13353 13368 13358 13424
rect 13414 13368 22742 13424
rect 22798 13368 22803 13424
rect 13353 13366 22803 13368
rect 13353 13363 13419 13366
rect 22737 13363 22803 13366
rect 4889 13290 4955 13293
rect 5993 13290 6059 13293
rect 4889 13288 6059 13290
rect 4889 13232 4894 13288
rect 4950 13232 5998 13288
rect 6054 13232 6059 13288
rect 4889 13230 6059 13232
rect 4889 13227 4955 13230
rect 5993 13227 6059 13230
rect 11237 13290 11303 13293
rect 11973 13290 12039 13293
rect 18781 13290 18847 13293
rect 11237 13288 18847 13290
rect 11237 13232 11242 13288
rect 11298 13232 11978 13288
rect 12034 13232 18786 13288
rect 18842 13232 18847 13288
rect 11237 13230 18847 13232
rect 11237 13227 11303 13230
rect 11973 13227 12039 13230
rect 18781 13227 18847 13230
rect 16573 13154 16639 13157
rect 17677 13154 17743 13157
rect 16573 13152 17743 13154
rect 16573 13096 16578 13152
rect 16634 13096 17682 13152
rect 17738 13096 17743 13152
rect 16573 13094 17743 13096
rect 16573 13091 16639 13094
rect 17677 13091 17743 13094
rect 6626 13088 6942 13089
rect 6626 13024 6632 13088
rect 6696 13024 6712 13088
rect 6776 13024 6792 13088
rect 6856 13024 6872 13088
rect 6936 13024 6942 13088
rect 6626 13023 6942 13024
rect 12307 13088 12623 13089
rect 12307 13024 12313 13088
rect 12377 13024 12393 13088
rect 12457 13024 12473 13088
rect 12537 13024 12553 13088
rect 12617 13024 12623 13088
rect 12307 13023 12623 13024
rect 17988 13088 18304 13089
rect 17988 13024 17994 13088
rect 18058 13024 18074 13088
rect 18138 13024 18154 13088
rect 18218 13024 18234 13088
rect 18298 13024 18304 13088
rect 17988 13023 18304 13024
rect 23669 13088 23985 13089
rect 23669 13024 23675 13088
rect 23739 13024 23755 13088
rect 23819 13024 23835 13088
rect 23899 13024 23915 13088
rect 23979 13024 23985 13088
rect 23669 13023 23985 13024
rect 14457 12882 14523 12885
rect 17217 12882 17283 12885
rect 19149 12882 19215 12885
rect 14457 12880 19215 12882
rect 14457 12824 14462 12880
rect 14518 12824 17222 12880
rect 17278 12824 19154 12880
rect 19210 12824 19215 12880
rect 14457 12822 19215 12824
rect 14457 12819 14523 12822
rect 17217 12819 17283 12822
rect 19149 12819 19215 12822
rect 3786 12544 4102 12545
rect 3786 12480 3792 12544
rect 3856 12480 3872 12544
rect 3936 12480 3952 12544
rect 4016 12480 4032 12544
rect 4096 12480 4102 12544
rect 3786 12479 4102 12480
rect 9467 12544 9783 12545
rect 9467 12480 9473 12544
rect 9537 12480 9553 12544
rect 9617 12480 9633 12544
rect 9697 12480 9713 12544
rect 9777 12480 9783 12544
rect 9467 12479 9783 12480
rect 15148 12544 15464 12545
rect 15148 12480 15154 12544
rect 15218 12480 15234 12544
rect 15298 12480 15314 12544
rect 15378 12480 15394 12544
rect 15458 12480 15464 12544
rect 15148 12479 15464 12480
rect 20829 12544 21145 12545
rect 20829 12480 20835 12544
rect 20899 12480 20915 12544
rect 20979 12480 20995 12544
rect 21059 12480 21075 12544
rect 21139 12480 21145 12544
rect 20829 12479 21145 12480
rect 17125 12338 17191 12341
rect 19333 12338 19399 12341
rect 17125 12336 19399 12338
rect 17125 12280 17130 12336
rect 17186 12280 19338 12336
rect 19394 12280 19399 12336
rect 17125 12278 19399 12280
rect 17125 12275 17191 12278
rect 19333 12275 19399 12278
rect 19742 12276 19748 12340
rect 19812 12338 19818 12340
rect 21081 12338 21147 12341
rect 19812 12336 21147 12338
rect 19812 12280 21086 12336
rect 21142 12280 21147 12336
rect 19812 12278 21147 12280
rect 19812 12276 19818 12278
rect 21081 12275 21147 12278
rect 5441 12068 5507 12069
rect 5390 12004 5396 12068
rect 5460 12066 5507 12068
rect 5460 12064 5552 12066
rect 5502 12008 5552 12064
rect 5460 12006 5552 12008
rect 5460 12004 5507 12006
rect 5441 12003 5507 12004
rect 6626 12000 6942 12001
rect 6626 11936 6632 12000
rect 6696 11936 6712 12000
rect 6776 11936 6792 12000
rect 6856 11936 6872 12000
rect 6936 11936 6942 12000
rect 6626 11935 6942 11936
rect 12307 12000 12623 12001
rect 12307 11936 12313 12000
rect 12377 11936 12393 12000
rect 12457 11936 12473 12000
rect 12537 11936 12553 12000
rect 12617 11936 12623 12000
rect 12307 11935 12623 11936
rect 17988 12000 18304 12001
rect 17988 11936 17994 12000
rect 18058 11936 18074 12000
rect 18138 11936 18154 12000
rect 18218 11936 18234 12000
rect 18298 11936 18304 12000
rect 17988 11935 18304 11936
rect 23669 12000 23985 12001
rect 23669 11936 23675 12000
rect 23739 11936 23755 12000
rect 23819 11936 23835 12000
rect 23899 11936 23915 12000
rect 23979 11936 23985 12000
rect 23669 11935 23985 11936
rect 15377 11794 15443 11797
rect 17861 11794 17927 11797
rect 15377 11792 17927 11794
rect 15377 11736 15382 11792
rect 15438 11736 17866 11792
rect 17922 11736 17927 11792
rect 15377 11734 17927 11736
rect 15377 11731 15443 11734
rect 17861 11731 17927 11734
rect 3786 11456 4102 11457
rect 3786 11392 3792 11456
rect 3856 11392 3872 11456
rect 3936 11392 3952 11456
rect 4016 11392 4032 11456
rect 4096 11392 4102 11456
rect 3786 11391 4102 11392
rect 9467 11456 9783 11457
rect 9467 11392 9473 11456
rect 9537 11392 9553 11456
rect 9617 11392 9633 11456
rect 9697 11392 9713 11456
rect 9777 11392 9783 11456
rect 9467 11391 9783 11392
rect 15148 11456 15464 11457
rect 15148 11392 15154 11456
rect 15218 11392 15234 11456
rect 15298 11392 15314 11456
rect 15378 11392 15394 11456
rect 15458 11392 15464 11456
rect 15148 11391 15464 11392
rect 20829 11456 21145 11457
rect 20829 11392 20835 11456
rect 20899 11392 20915 11456
rect 20979 11392 20995 11456
rect 21059 11392 21075 11456
rect 21139 11392 21145 11456
rect 20829 11391 21145 11392
rect 17033 11114 17099 11117
rect 17718 11114 17724 11116
rect 17033 11112 17724 11114
rect 17033 11056 17038 11112
rect 17094 11056 17724 11112
rect 17033 11054 17724 11056
rect 17033 11051 17099 11054
rect 17718 11052 17724 11054
rect 17788 11052 17794 11116
rect 6626 10912 6942 10913
rect 6626 10848 6632 10912
rect 6696 10848 6712 10912
rect 6776 10848 6792 10912
rect 6856 10848 6872 10912
rect 6936 10848 6942 10912
rect 6626 10847 6942 10848
rect 12307 10912 12623 10913
rect 12307 10848 12313 10912
rect 12377 10848 12393 10912
rect 12457 10848 12473 10912
rect 12537 10848 12553 10912
rect 12617 10848 12623 10912
rect 12307 10847 12623 10848
rect 17988 10912 18304 10913
rect 17988 10848 17994 10912
rect 18058 10848 18074 10912
rect 18138 10848 18154 10912
rect 18218 10848 18234 10912
rect 18298 10848 18304 10912
rect 17988 10847 18304 10848
rect 23669 10912 23985 10913
rect 23669 10848 23675 10912
rect 23739 10848 23755 10912
rect 23819 10848 23835 10912
rect 23899 10848 23915 10912
rect 23979 10848 23985 10912
rect 23669 10847 23985 10848
rect 2957 10706 3023 10709
rect 8477 10706 8543 10709
rect 2957 10704 8543 10706
rect 2957 10648 2962 10704
rect 3018 10648 8482 10704
rect 8538 10648 8543 10704
rect 2957 10646 8543 10648
rect 2957 10643 3023 10646
rect 8477 10643 8543 10646
rect 15193 10570 15259 10573
rect 19333 10570 19399 10573
rect 20437 10570 20503 10573
rect 15193 10568 20503 10570
rect 15193 10512 15198 10568
rect 15254 10512 19338 10568
rect 19394 10512 20442 10568
rect 20498 10512 20503 10568
rect 15193 10510 20503 10512
rect 15193 10507 15259 10510
rect 19333 10507 19399 10510
rect 20437 10507 20503 10510
rect 3786 10368 4102 10369
rect 3786 10304 3792 10368
rect 3856 10304 3872 10368
rect 3936 10304 3952 10368
rect 4016 10304 4032 10368
rect 4096 10304 4102 10368
rect 3786 10303 4102 10304
rect 9467 10368 9783 10369
rect 9467 10304 9473 10368
rect 9537 10304 9553 10368
rect 9617 10304 9633 10368
rect 9697 10304 9713 10368
rect 9777 10304 9783 10368
rect 9467 10303 9783 10304
rect 15148 10368 15464 10369
rect 15148 10304 15154 10368
rect 15218 10304 15234 10368
rect 15298 10304 15314 10368
rect 15378 10304 15394 10368
rect 15458 10304 15464 10368
rect 15148 10303 15464 10304
rect 20829 10368 21145 10369
rect 20829 10304 20835 10368
rect 20899 10304 20915 10368
rect 20979 10304 20995 10368
rect 21059 10304 21075 10368
rect 21139 10304 21145 10368
rect 20829 10303 21145 10304
rect 17769 9890 17835 9893
rect 17726 9888 17835 9890
rect 17726 9832 17774 9888
rect 17830 9832 17835 9888
rect 17726 9827 17835 9832
rect 6626 9824 6942 9825
rect 6626 9760 6632 9824
rect 6696 9760 6712 9824
rect 6776 9760 6792 9824
rect 6856 9760 6872 9824
rect 6936 9760 6942 9824
rect 6626 9759 6942 9760
rect 12307 9824 12623 9825
rect 12307 9760 12313 9824
rect 12377 9760 12393 9824
rect 12457 9760 12473 9824
rect 12537 9760 12553 9824
rect 12617 9760 12623 9824
rect 12307 9759 12623 9760
rect 6310 9692 6316 9756
rect 6380 9692 6386 9756
rect 1669 9618 1735 9621
rect 4654 9618 4660 9620
rect 1669 9616 4660 9618
rect 1669 9560 1674 9616
rect 1730 9560 4660 9616
rect 1669 9558 4660 9560
rect 1669 9555 1735 9558
rect 4654 9556 4660 9558
rect 4724 9556 4730 9620
rect 4889 9618 4955 9621
rect 6318 9618 6378 9692
rect 17726 9690 17786 9827
rect 17988 9824 18304 9825
rect 17988 9760 17994 9824
rect 18058 9760 18074 9824
rect 18138 9760 18154 9824
rect 18218 9760 18234 9824
rect 18298 9760 18304 9824
rect 17988 9759 18304 9760
rect 23669 9824 23985 9825
rect 23669 9760 23675 9824
rect 23739 9760 23755 9824
rect 23819 9760 23835 9824
rect 23899 9760 23915 9824
rect 23979 9760 23985 9824
rect 23669 9759 23985 9760
rect 17953 9690 18019 9693
rect 17726 9688 18019 9690
rect 17726 9632 17958 9688
rect 18014 9632 18019 9688
rect 17726 9630 18019 9632
rect 17953 9627 18019 9630
rect 6545 9618 6611 9621
rect 4889 9616 6611 9618
rect 4889 9560 4894 9616
rect 4950 9560 6550 9616
rect 6606 9560 6611 9616
rect 4889 9558 6611 9560
rect 4889 9555 4955 9558
rect 6545 9555 6611 9558
rect 9765 9618 9831 9621
rect 12157 9618 12223 9621
rect 9765 9616 12223 9618
rect 9765 9560 9770 9616
rect 9826 9560 12162 9616
rect 12218 9560 12223 9616
rect 9765 9558 12223 9560
rect 9765 9555 9831 9558
rect 12157 9555 12223 9558
rect 1485 9482 1551 9485
rect 5717 9484 5783 9485
rect 5717 9482 5764 9484
rect 1485 9480 5764 9482
rect 1485 9424 1490 9480
rect 1546 9424 5722 9480
rect 1485 9422 5764 9424
rect 1485 9419 1551 9422
rect 5717 9420 5764 9422
rect 5828 9420 5834 9484
rect 5717 9419 5783 9420
rect 10225 9346 10291 9349
rect 10869 9346 10935 9349
rect 10225 9344 10935 9346
rect 10225 9288 10230 9344
rect 10286 9288 10874 9344
rect 10930 9288 10935 9344
rect 10225 9286 10935 9288
rect 10225 9283 10291 9286
rect 10869 9283 10935 9286
rect 3786 9280 4102 9281
rect 3786 9216 3792 9280
rect 3856 9216 3872 9280
rect 3936 9216 3952 9280
rect 4016 9216 4032 9280
rect 4096 9216 4102 9280
rect 3786 9215 4102 9216
rect 9467 9280 9783 9281
rect 9467 9216 9473 9280
rect 9537 9216 9553 9280
rect 9617 9216 9633 9280
rect 9697 9216 9713 9280
rect 9777 9216 9783 9280
rect 9467 9215 9783 9216
rect 15148 9280 15464 9281
rect 15148 9216 15154 9280
rect 15218 9216 15234 9280
rect 15298 9216 15314 9280
rect 15378 9216 15394 9280
rect 15458 9216 15464 9280
rect 15148 9215 15464 9216
rect 20829 9280 21145 9281
rect 20829 9216 20835 9280
rect 20899 9216 20915 9280
rect 20979 9216 20995 9280
rect 21059 9216 21075 9280
rect 21139 9216 21145 9280
rect 20829 9215 21145 9216
rect 6626 8736 6942 8737
rect 6626 8672 6632 8736
rect 6696 8672 6712 8736
rect 6776 8672 6792 8736
rect 6856 8672 6872 8736
rect 6936 8672 6942 8736
rect 6626 8671 6942 8672
rect 12307 8736 12623 8737
rect 12307 8672 12313 8736
rect 12377 8672 12393 8736
rect 12457 8672 12473 8736
rect 12537 8672 12553 8736
rect 12617 8672 12623 8736
rect 12307 8671 12623 8672
rect 17988 8736 18304 8737
rect 17988 8672 17994 8736
rect 18058 8672 18074 8736
rect 18138 8672 18154 8736
rect 18218 8672 18234 8736
rect 18298 8672 18304 8736
rect 17988 8671 18304 8672
rect 23669 8736 23985 8737
rect 23669 8672 23675 8736
rect 23739 8672 23755 8736
rect 23819 8672 23835 8736
rect 23899 8672 23915 8736
rect 23979 8672 23985 8736
rect 23669 8671 23985 8672
rect 18965 8394 19031 8397
rect 22001 8394 22067 8397
rect 18965 8392 22067 8394
rect 18965 8336 18970 8392
rect 19026 8336 22006 8392
rect 22062 8336 22067 8392
rect 18965 8334 22067 8336
rect 18965 8331 19031 8334
rect 22001 8331 22067 8334
rect 3786 8192 4102 8193
rect 3786 8128 3792 8192
rect 3856 8128 3872 8192
rect 3936 8128 3952 8192
rect 4016 8128 4032 8192
rect 4096 8128 4102 8192
rect 3786 8127 4102 8128
rect 9467 8192 9783 8193
rect 9467 8128 9473 8192
rect 9537 8128 9553 8192
rect 9617 8128 9633 8192
rect 9697 8128 9713 8192
rect 9777 8128 9783 8192
rect 9467 8127 9783 8128
rect 15148 8192 15464 8193
rect 15148 8128 15154 8192
rect 15218 8128 15234 8192
rect 15298 8128 15314 8192
rect 15378 8128 15394 8192
rect 15458 8128 15464 8192
rect 15148 8127 15464 8128
rect 20829 8192 21145 8193
rect 20829 8128 20835 8192
rect 20899 8128 20915 8192
rect 20979 8128 20995 8192
rect 21059 8128 21075 8192
rect 21139 8128 21145 8192
rect 20829 8127 21145 8128
rect 6626 7648 6942 7649
rect 6626 7584 6632 7648
rect 6696 7584 6712 7648
rect 6776 7584 6792 7648
rect 6856 7584 6872 7648
rect 6936 7584 6942 7648
rect 6626 7583 6942 7584
rect 12307 7648 12623 7649
rect 12307 7584 12313 7648
rect 12377 7584 12393 7648
rect 12457 7584 12473 7648
rect 12537 7584 12553 7648
rect 12617 7584 12623 7648
rect 12307 7583 12623 7584
rect 17988 7648 18304 7649
rect 17988 7584 17994 7648
rect 18058 7584 18074 7648
rect 18138 7584 18154 7648
rect 18218 7584 18234 7648
rect 18298 7584 18304 7648
rect 17988 7583 18304 7584
rect 23669 7648 23985 7649
rect 23669 7584 23675 7648
rect 23739 7584 23755 7648
rect 23819 7584 23835 7648
rect 23899 7584 23915 7648
rect 23979 7584 23985 7648
rect 23669 7583 23985 7584
rect 3786 7104 4102 7105
rect 3786 7040 3792 7104
rect 3856 7040 3872 7104
rect 3936 7040 3952 7104
rect 4016 7040 4032 7104
rect 4096 7040 4102 7104
rect 3786 7039 4102 7040
rect 9467 7104 9783 7105
rect 9467 7040 9473 7104
rect 9537 7040 9553 7104
rect 9617 7040 9633 7104
rect 9697 7040 9713 7104
rect 9777 7040 9783 7104
rect 9467 7039 9783 7040
rect 15148 7104 15464 7105
rect 15148 7040 15154 7104
rect 15218 7040 15234 7104
rect 15298 7040 15314 7104
rect 15378 7040 15394 7104
rect 15458 7040 15464 7104
rect 15148 7039 15464 7040
rect 20829 7104 21145 7105
rect 20829 7040 20835 7104
rect 20899 7040 20915 7104
rect 20979 7040 20995 7104
rect 21059 7040 21075 7104
rect 21139 7040 21145 7104
rect 20829 7039 21145 7040
rect 14590 6836 14596 6900
rect 14660 6898 14666 6900
rect 22185 6898 22251 6901
rect 14660 6896 22251 6898
rect 14660 6840 22190 6896
rect 22246 6840 22251 6896
rect 14660 6838 22251 6840
rect 14660 6836 14666 6838
rect 22185 6835 22251 6838
rect 6821 6762 6887 6765
rect 18689 6762 18755 6765
rect 6821 6760 18755 6762
rect 6821 6704 6826 6760
rect 6882 6704 18694 6760
rect 18750 6704 18755 6760
rect 6821 6702 18755 6704
rect 6821 6699 6887 6702
rect 18689 6699 18755 6702
rect 6626 6560 6942 6561
rect 6626 6496 6632 6560
rect 6696 6496 6712 6560
rect 6776 6496 6792 6560
rect 6856 6496 6872 6560
rect 6936 6496 6942 6560
rect 6626 6495 6942 6496
rect 12307 6560 12623 6561
rect 12307 6496 12313 6560
rect 12377 6496 12393 6560
rect 12457 6496 12473 6560
rect 12537 6496 12553 6560
rect 12617 6496 12623 6560
rect 12307 6495 12623 6496
rect 17988 6560 18304 6561
rect 17988 6496 17994 6560
rect 18058 6496 18074 6560
rect 18138 6496 18154 6560
rect 18218 6496 18234 6560
rect 18298 6496 18304 6560
rect 17988 6495 18304 6496
rect 23669 6560 23985 6561
rect 23669 6496 23675 6560
rect 23739 6496 23755 6560
rect 23819 6496 23835 6560
rect 23899 6496 23915 6560
rect 23979 6496 23985 6560
rect 23669 6495 23985 6496
rect 10685 6082 10751 6085
rect 13997 6082 14063 6085
rect 10685 6080 14063 6082
rect 10685 6024 10690 6080
rect 10746 6024 14002 6080
rect 14058 6024 14063 6080
rect 10685 6022 14063 6024
rect 10685 6019 10751 6022
rect 13997 6019 14063 6022
rect 3786 6016 4102 6017
rect 3786 5952 3792 6016
rect 3856 5952 3872 6016
rect 3936 5952 3952 6016
rect 4016 5952 4032 6016
rect 4096 5952 4102 6016
rect 3786 5951 4102 5952
rect 9467 6016 9783 6017
rect 9467 5952 9473 6016
rect 9537 5952 9553 6016
rect 9617 5952 9633 6016
rect 9697 5952 9713 6016
rect 9777 5952 9783 6016
rect 9467 5951 9783 5952
rect 15148 6016 15464 6017
rect 15148 5952 15154 6016
rect 15218 5952 15234 6016
rect 15298 5952 15314 6016
rect 15378 5952 15394 6016
rect 15458 5952 15464 6016
rect 15148 5951 15464 5952
rect 20829 6016 21145 6017
rect 20829 5952 20835 6016
rect 20899 5952 20915 6016
rect 20979 5952 20995 6016
rect 21059 5952 21075 6016
rect 21139 5952 21145 6016
rect 20829 5951 21145 5952
rect 3049 5674 3115 5677
rect 3601 5674 3667 5677
rect 3049 5672 3667 5674
rect 3049 5616 3054 5672
rect 3110 5616 3606 5672
rect 3662 5616 3667 5672
rect 3049 5614 3667 5616
rect 3049 5611 3115 5614
rect 3601 5611 3667 5614
rect 19926 5612 19932 5676
rect 19996 5674 20002 5676
rect 21173 5674 21239 5677
rect 23289 5674 23355 5677
rect 19996 5672 23355 5674
rect 19996 5616 21178 5672
rect 21234 5616 23294 5672
rect 23350 5616 23355 5672
rect 19996 5614 23355 5616
rect 19996 5612 20002 5614
rect 21173 5611 21239 5614
rect 23289 5611 23355 5614
rect 6626 5472 6942 5473
rect 6626 5408 6632 5472
rect 6696 5408 6712 5472
rect 6776 5408 6792 5472
rect 6856 5408 6872 5472
rect 6936 5408 6942 5472
rect 6626 5407 6942 5408
rect 12307 5472 12623 5473
rect 12307 5408 12313 5472
rect 12377 5408 12393 5472
rect 12457 5408 12473 5472
rect 12537 5408 12553 5472
rect 12617 5408 12623 5472
rect 12307 5407 12623 5408
rect 17988 5472 18304 5473
rect 17988 5408 17994 5472
rect 18058 5408 18074 5472
rect 18138 5408 18154 5472
rect 18218 5408 18234 5472
rect 18298 5408 18304 5472
rect 17988 5407 18304 5408
rect 23669 5472 23985 5473
rect 23669 5408 23675 5472
rect 23739 5408 23755 5472
rect 23819 5408 23835 5472
rect 23899 5408 23915 5472
rect 23979 5408 23985 5472
rect 23669 5407 23985 5408
rect 11421 5266 11487 5269
rect 15837 5266 15903 5269
rect 11421 5264 15903 5266
rect 11421 5208 11426 5264
rect 11482 5208 15842 5264
rect 15898 5208 15903 5264
rect 11421 5206 15903 5208
rect 11421 5203 11487 5206
rect 15837 5203 15903 5206
rect 17718 5204 17724 5268
rect 17788 5266 17794 5268
rect 19241 5266 19307 5269
rect 17788 5264 19307 5266
rect 17788 5208 19246 5264
rect 19302 5208 19307 5264
rect 17788 5206 19307 5208
rect 17788 5204 17794 5206
rect 19241 5203 19307 5206
rect 6637 5130 6703 5133
rect 12249 5130 12315 5133
rect 18413 5130 18479 5133
rect 6637 5128 18479 5130
rect 6637 5072 6642 5128
rect 6698 5072 12254 5128
rect 12310 5072 18418 5128
rect 18474 5072 18479 5128
rect 6637 5070 18479 5072
rect 6637 5067 6703 5070
rect 12249 5067 12315 5070
rect 18413 5067 18479 5070
rect 5809 4994 5875 4997
rect 7373 4994 7439 4997
rect 5809 4992 7439 4994
rect 5809 4936 5814 4992
rect 5870 4936 7378 4992
rect 7434 4936 7439 4992
rect 5809 4934 7439 4936
rect 5809 4931 5875 4934
rect 7373 4931 7439 4934
rect 3786 4928 4102 4929
rect 3786 4864 3792 4928
rect 3856 4864 3872 4928
rect 3936 4864 3952 4928
rect 4016 4864 4032 4928
rect 4096 4864 4102 4928
rect 3786 4863 4102 4864
rect 9467 4928 9783 4929
rect 9467 4864 9473 4928
rect 9537 4864 9553 4928
rect 9617 4864 9633 4928
rect 9697 4864 9713 4928
rect 9777 4864 9783 4928
rect 9467 4863 9783 4864
rect 15148 4928 15464 4929
rect 15148 4864 15154 4928
rect 15218 4864 15234 4928
rect 15298 4864 15314 4928
rect 15378 4864 15394 4928
rect 15458 4864 15464 4928
rect 15148 4863 15464 4864
rect 20829 4928 21145 4929
rect 20829 4864 20835 4928
rect 20899 4864 20915 4928
rect 20979 4864 20995 4928
rect 21059 4864 21075 4928
rect 21139 4864 21145 4928
rect 20829 4863 21145 4864
rect 6626 4384 6942 4385
rect 6626 4320 6632 4384
rect 6696 4320 6712 4384
rect 6776 4320 6792 4384
rect 6856 4320 6872 4384
rect 6936 4320 6942 4384
rect 6626 4319 6942 4320
rect 12307 4384 12623 4385
rect 12307 4320 12313 4384
rect 12377 4320 12393 4384
rect 12457 4320 12473 4384
rect 12537 4320 12553 4384
rect 12617 4320 12623 4384
rect 12307 4319 12623 4320
rect 17988 4384 18304 4385
rect 17988 4320 17994 4384
rect 18058 4320 18074 4384
rect 18138 4320 18154 4384
rect 18218 4320 18234 4384
rect 18298 4320 18304 4384
rect 17988 4319 18304 4320
rect 23669 4384 23985 4385
rect 23669 4320 23675 4384
rect 23739 4320 23755 4384
rect 23819 4320 23835 4384
rect 23899 4320 23915 4384
rect 23979 4320 23985 4384
rect 23669 4319 23985 4320
rect 13537 4178 13603 4181
rect 15929 4178 15995 4181
rect 16297 4178 16363 4181
rect 13537 4176 16363 4178
rect 13537 4120 13542 4176
rect 13598 4120 15934 4176
rect 15990 4120 16302 4176
rect 16358 4120 16363 4176
rect 13537 4118 16363 4120
rect 13537 4115 13603 4118
rect 15929 4115 15995 4118
rect 16297 4115 16363 4118
rect 5758 3980 5764 4044
rect 5828 4042 5834 4044
rect 6545 4042 6611 4045
rect 5828 4040 6611 4042
rect 5828 3984 6550 4040
rect 6606 3984 6611 4040
rect 5828 3982 6611 3984
rect 5828 3980 5834 3982
rect 6545 3979 6611 3982
rect 3786 3840 4102 3841
rect 3786 3776 3792 3840
rect 3856 3776 3872 3840
rect 3936 3776 3952 3840
rect 4016 3776 4032 3840
rect 4096 3776 4102 3840
rect 3786 3775 4102 3776
rect 9467 3840 9783 3841
rect 9467 3776 9473 3840
rect 9537 3776 9553 3840
rect 9617 3776 9633 3840
rect 9697 3776 9713 3840
rect 9777 3776 9783 3840
rect 9467 3775 9783 3776
rect 15148 3840 15464 3841
rect 15148 3776 15154 3840
rect 15218 3776 15234 3840
rect 15298 3776 15314 3840
rect 15378 3776 15394 3840
rect 15458 3776 15464 3840
rect 15148 3775 15464 3776
rect 20829 3840 21145 3841
rect 20829 3776 20835 3840
rect 20899 3776 20915 3840
rect 20979 3776 20995 3840
rect 21059 3776 21075 3840
rect 21139 3776 21145 3840
rect 20829 3775 21145 3776
rect 7189 3634 7255 3637
rect 14917 3634 14983 3637
rect 7189 3632 14983 3634
rect 7189 3576 7194 3632
rect 7250 3576 14922 3632
rect 14978 3576 14983 3632
rect 7189 3574 14983 3576
rect 7189 3571 7255 3574
rect 14917 3571 14983 3574
rect 5441 3498 5507 3501
rect 11421 3498 11487 3501
rect 18321 3498 18387 3501
rect 5441 3496 18387 3498
rect 5441 3440 5446 3496
rect 5502 3440 11426 3496
rect 11482 3440 18326 3496
rect 18382 3440 18387 3496
rect 5441 3438 18387 3440
rect 5441 3435 5507 3438
rect 11421 3435 11487 3438
rect 18321 3435 18387 3438
rect 7097 3362 7163 3365
rect 11697 3362 11763 3365
rect 7097 3360 11763 3362
rect 7097 3304 7102 3360
rect 7158 3304 11702 3360
rect 11758 3304 11763 3360
rect 7097 3302 11763 3304
rect 7097 3299 7163 3302
rect 11697 3299 11763 3302
rect 6626 3296 6942 3297
rect 6626 3232 6632 3296
rect 6696 3232 6712 3296
rect 6776 3232 6792 3296
rect 6856 3232 6872 3296
rect 6936 3232 6942 3296
rect 6626 3231 6942 3232
rect 12307 3296 12623 3297
rect 12307 3232 12313 3296
rect 12377 3232 12393 3296
rect 12457 3232 12473 3296
rect 12537 3232 12553 3296
rect 12617 3232 12623 3296
rect 12307 3231 12623 3232
rect 17988 3296 18304 3297
rect 17988 3232 17994 3296
rect 18058 3232 18074 3296
rect 18138 3232 18154 3296
rect 18218 3232 18234 3296
rect 18298 3232 18304 3296
rect 17988 3231 18304 3232
rect 23669 3296 23985 3297
rect 23669 3232 23675 3296
rect 23739 3232 23755 3296
rect 23819 3232 23835 3296
rect 23899 3232 23915 3296
rect 23979 3232 23985 3296
rect 23669 3231 23985 3232
rect 11789 3226 11855 3229
rect 7238 3224 11855 3226
rect 7238 3168 11794 3224
rect 11850 3168 11855 3224
rect 7238 3166 11855 3168
rect 4286 3028 4292 3092
rect 4356 3090 4362 3092
rect 5390 3090 5396 3092
rect 4356 3030 5396 3090
rect 4356 3028 4362 3030
rect 5390 3028 5396 3030
rect 5460 3090 5466 3092
rect 7238 3090 7298 3166
rect 11789 3163 11855 3166
rect 5460 3030 7298 3090
rect 9949 3090 10015 3093
rect 13721 3090 13787 3093
rect 9949 3088 13787 3090
rect 9949 3032 9954 3088
rect 10010 3032 13726 3088
rect 13782 3032 13787 3088
rect 9949 3030 13787 3032
rect 5460 3028 5466 3030
rect 9949 3027 10015 3030
rect 13721 3027 13787 3030
rect 2957 2954 3023 2957
rect 14549 2954 14615 2957
rect 2957 2952 14615 2954
rect 2957 2896 2962 2952
rect 3018 2896 14554 2952
rect 14610 2896 14615 2952
rect 2957 2894 14615 2896
rect 2957 2891 3023 2894
rect 14549 2891 14615 2894
rect 3786 2752 4102 2753
rect 3786 2688 3792 2752
rect 3856 2688 3872 2752
rect 3936 2688 3952 2752
rect 4016 2688 4032 2752
rect 4096 2688 4102 2752
rect 3786 2687 4102 2688
rect 9467 2752 9783 2753
rect 9467 2688 9473 2752
rect 9537 2688 9553 2752
rect 9617 2688 9633 2752
rect 9697 2688 9713 2752
rect 9777 2688 9783 2752
rect 9467 2687 9783 2688
rect 15148 2752 15464 2753
rect 15148 2688 15154 2752
rect 15218 2688 15234 2752
rect 15298 2688 15314 2752
rect 15378 2688 15394 2752
rect 15458 2688 15464 2752
rect 15148 2687 15464 2688
rect 20829 2752 21145 2753
rect 20829 2688 20835 2752
rect 20899 2688 20915 2752
rect 20979 2688 20995 2752
rect 21059 2688 21075 2752
rect 21139 2688 21145 2752
rect 20829 2687 21145 2688
rect 3417 2546 3483 2549
rect 4286 2546 4292 2548
rect 3417 2544 4292 2546
rect 3417 2488 3422 2544
rect 3478 2488 4292 2544
rect 3417 2486 4292 2488
rect 3417 2483 3483 2486
rect 4286 2484 4292 2486
rect 4356 2484 4362 2548
rect 6626 2208 6942 2209
rect 6626 2144 6632 2208
rect 6696 2144 6712 2208
rect 6776 2144 6792 2208
rect 6856 2144 6872 2208
rect 6936 2144 6942 2208
rect 6626 2143 6942 2144
rect 12307 2208 12623 2209
rect 12307 2144 12313 2208
rect 12377 2144 12393 2208
rect 12457 2144 12473 2208
rect 12537 2144 12553 2208
rect 12617 2144 12623 2208
rect 12307 2143 12623 2144
rect 17988 2208 18304 2209
rect 17988 2144 17994 2208
rect 18058 2144 18074 2208
rect 18138 2144 18154 2208
rect 18218 2144 18234 2208
rect 18298 2144 18304 2208
rect 17988 2143 18304 2144
rect 23669 2208 23985 2209
rect 23669 2144 23675 2208
rect 23739 2144 23755 2208
rect 23819 2144 23835 2208
rect 23899 2144 23915 2208
rect 23979 2144 23985 2208
rect 23669 2143 23985 2144
<< via3 >>
rect 3792 22332 3856 22336
rect 3792 22276 3796 22332
rect 3796 22276 3852 22332
rect 3852 22276 3856 22332
rect 3792 22272 3856 22276
rect 3872 22332 3936 22336
rect 3872 22276 3876 22332
rect 3876 22276 3932 22332
rect 3932 22276 3936 22332
rect 3872 22272 3936 22276
rect 3952 22332 4016 22336
rect 3952 22276 3956 22332
rect 3956 22276 4012 22332
rect 4012 22276 4016 22332
rect 3952 22272 4016 22276
rect 4032 22332 4096 22336
rect 4032 22276 4036 22332
rect 4036 22276 4092 22332
rect 4092 22276 4096 22332
rect 4032 22272 4096 22276
rect 9473 22332 9537 22336
rect 9473 22276 9477 22332
rect 9477 22276 9533 22332
rect 9533 22276 9537 22332
rect 9473 22272 9537 22276
rect 9553 22332 9617 22336
rect 9553 22276 9557 22332
rect 9557 22276 9613 22332
rect 9613 22276 9617 22332
rect 9553 22272 9617 22276
rect 9633 22332 9697 22336
rect 9633 22276 9637 22332
rect 9637 22276 9693 22332
rect 9693 22276 9697 22332
rect 9633 22272 9697 22276
rect 9713 22332 9777 22336
rect 9713 22276 9717 22332
rect 9717 22276 9773 22332
rect 9773 22276 9777 22332
rect 9713 22272 9777 22276
rect 15154 22332 15218 22336
rect 15154 22276 15158 22332
rect 15158 22276 15214 22332
rect 15214 22276 15218 22332
rect 15154 22272 15218 22276
rect 15234 22332 15298 22336
rect 15234 22276 15238 22332
rect 15238 22276 15294 22332
rect 15294 22276 15298 22332
rect 15234 22272 15298 22276
rect 15314 22332 15378 22336
rect 15314 22276 15318 22332
rect 15318 22276 15374 22332
rect 15374 22276 15378 22332
rect 15314 22272 15378 22276
rect 15394 22332 15458 22336
rect 15394 22276 15398 22332
rect 15398 22276 15454 22332
rect 15454 22276 15458 22332
rect 15394 22272 15458 22276
rect 20835 22332 20899 22336
rect 20835 22276 20839 22332
rect 20839 22276 20895 22332
rect 20895 22276 20899 22332
rect 20835 22272 20899 22276
rect 20915 22332 20979 22336
rect 20915 22276 20919 22332
rect 20919 22276 20975 22332
rect 20975 22276 20979 22332
rect 20915 22272 20979 22276
rect 20995 22332 21059 22336
rect 20995 22276 20999 22332
rect 20999 22276 21055 22332
rect 21055 22276 21059 22332
rect 20995 22272 21059 22276
rect 21075 22332 21139 22336
rect 21075 22276 21079 22332
rect 21079 22276 21135 22332
rect 21135 22276 21139 22332
rect 21075 22272 21139 22276
rect 6632 21788 6696 21792
rect 6632 21732 6636 21788
rect 6636 21732 6692 21788
rect 6692 21732 6696 21788
rect 6632 21728 6696 21732
rect 6712 21788 6776 21792
rect 6712 21732 6716 21788
rect 6716 21732 6772 21788
rect 6772 21732 6776 21788
rect 6712 21728 6776 21732
rect 6792 21788 6856 21792
rect 6792 21732 6796 21788
rect 6796 21732 6852 21788
rect 6852 21732 6856 21788
rect 6792 21728 6856 21732
rect 6872 21788 6936 21792
rect 6872 21732 6876 21788
rect 6876 21732 6932 21788
rect 6932 21732 6936 21788
rect 6872 21728 6936 21732
rect 12313 21788 12377 21792
rect 12313 21732 12317 21788
rect 12317 21732 12373 21788
rect 12373 21732 12377 21788
rect 12313 21728 12377 21732
rect 12393 21788 12457 21792
rect 12393 21732 12397 21788
rect 12397 21732 12453 21788
rect 12453 21732 12457 21788
rect 12393 21728 12457 21732
rect 12473 21788 12537 21792
rect 12473 21732 12477 21788
rect 12477 21732 12533 21788
rect 12533 21732 12537 21788
rect 12473 21728 12537 21732
rect 12553 21788 12617 21792
rect 12553 21732 12557 21788
rect 12557 21732 12613 21788
rect 12613 21732 12617 21788
rect 12553 21728 12617 21732
rect 17994 21788 18058 21792
rect 17994 21732 17998 21788
rect 17998 21732 18054 21788
rect 18054 21732 18058 21788
rect 17994 21728 18058 21732
rect 18074 21788 18138 21792
rect 18074 21732 18078 21788
rect 18078 21732 18134 21788
rect 18134 21732 18138 21788
rect 18074 21728 18138 21732
rect 18154 21788 18218 21792
rect 18154 21732 18158 21788
rect 18158 21732 18214 21788
rect 18214 21732 18218 21788
rect 18154 21728 18218 21732
rect 18234 21788 18298 21792
rect 18234 21732 18238 21788
rect 18238 21732 18294 21788
rect 18294 21732 18298 21788
rect 18234 21728 18298 21732
rect 23675 21788 23739 21792
rect 23675 21732 23679 21788
rect 23679 21732 23735 21788
rect 23735 21732 23739 21788
rect 23675 21728 23739 21732
rect 23755 21788 23819 21792
rect 23755 21732 23759 21788
rect 23759 21732 23815 21788
rect 23815 21732 23819 21788
rect 23755 21728 23819 21732
rect 23835 21788 23899 21792
rect 23835 21732 23839 21788
rect 23839 21732 23895 21788
rect 23895 21732 23899 21788
rect 23835 21728 23899 21732
rect 23915 21788 23979 21792
rect 23915 21732 23919 21788
rect 23919 21732 23975 21788
rect 23975 21732 23979 21788
rect 23915 21728 23979 21732
rect 14228 21312 14292 21316
rect 14228 21256 14242 21312
rect 14242 21256 14292 21312
rect 14228 21252 14292 21256
rect 3792 21244 3856 21248
rect 3792 21188 3796 21244
rect 3796 21188 3852 21244
rect 3852 21188 3856 21244
rect 3792 21184 3856 21188
rect 3872 21244 3936 21248
rect 3872 21188 3876 21244
rect 3876 21188 3932 21244
rect 3932 21188 3936 21244
rect 3872 21184 3936 21188
rect 3952 21244 4016 21248
rect 3952 21188 3956 21244
rect 3956 21188 4012 21244
rect 4012 21188 4016 21244
rect 3952 21184 4016 21188
rect 4032 21244 4096 21248
rect 4032 21188 4036 21244
rect 4036 21188 4092 21244
rect 4092 21188 4096 21244
rect 4032 21184 4096 21188
rect 9473 21244 9537 21248
rect 9473 21188 9477 21244
rect 9477 21188 9533 21244
rect 9533 21188 9537 21244
rect 9473 21184 9537 21188
rect 9553 21244 9617 21248
rect 9553 21188 9557 21244
rect 9557 21188 9613 21244
rect 9613 21188 9617 21244
rect 9553 21184 9617 21188
rect 9633 21244 9697 21248
rect 9633 21188 9637 21244
rect 9637 21188 9693 21244
rect 9693 21188 9697 21244
rect 9633 21184 9697 21188
rect 9713 21244 9777 21248
rect 9713 21188 9717 21244
rect 9717 21188 9773 21244
rect 9773 21188 9777 21244
rect 9713 21184 9777 21188
rect 15154 21244 15218 21248
rect 15154 21188 15158 21244
rect 15158 21188 15214 21244
rect 15214 21188 15218 21244
rect 15154 21184 15218 21188
rect 15234 21244 15298 21248
rect 15234 21188 15238 21244
rect 15238 21188 15294 21244
rect 15294 21188 15298 21244
rect 15234 21184 15298 21188
rect 15314 21244 15378 21248
rect 15314 21188 15318 21244
rect 15318 21188 15374 21244
rect 15374 21188 15378 21244
rect 15314 21184 15378 21188
rect 15394 21244 15458 21248
rect 15394 21188 15398 21244
rect 15398 21188 15454 21244
rect 15454 21188 15458 21244
rect 15394 21184 15458 21188
rect 20835 21244 20899 21248
rect 20835 21188 20839 21244
rect 20839 21188 20895 21244
rect 20895 21188 20899 21244
rect 20835 21184 20899 21188
rect 20915 21244 20979 21248
rect 20915 21188 20919 21244
rect 20919 21188 20975 21244
rect 20975 21188 20979 21244
rect 20915 21184 20979 21188
rect 20995 21244 21059 21248
rect 20995 21188 20999 21244
rect 20999 21188 21055 21244
rect 21055 21188 21059 21244
rect 20995 21184 21059 21188
rect 21075 21244 21139 21248
rect 21075 21188 21079 21244
rect 21079 21188 21135 21244
rect 21135 21188 21139 21244
rect 21075 21184 21139 21188
rect 4660 20768 4724 20772
rect 4660 20712 4674 20768
rect 4674 20712 4724 20768
rect 4660 20708 4724 20712
rect 19748 20708 19812 20772
rect 6632 20700 6696 20704
rect 6632 20644 6636 20700
rect 6636 20644 6692 20700
rect 6692 20644 6696 20700
rect 6632 20640 6696 20644
rect 6712 20700 6776 20704
rect 6712 20644 6716 20700
rect 6716 20644 6772 20700
rect 6772 20644 6776 20700
rect 6712 20640 6776 20644
rect 6792 20700 6856 20704
rect 6792 20644 6796 20700
rect 6796 20644 6852 20700
rect 6852 20644 6856 20700
rect 6792 20640 6856 20644
rect 6872 20700 6936 20704
rect 6872 20644 6876 20700
rect 6876 20644 6932 20700
rect 6932 20644 6936 20700
rect 6872 20640 6936 20644
rect 12313 20700 12377 20704
rect 12313 20644 12317 20700
rect 12317 20644 12373 20700
rect 12373 20644 12377 20700
rect 12313 20640 12377 20644
rect 12393 20700 12457 20704
rect 12393 20644 12397 20700
rect 12397 20644 12453 20700
rect 12453 20644 12457 20700
rect 12393 20640 12457 20644
rect 12473 20700 12537 20704
rect 12473 20644 12477 20700
rect 12477 20644 12533 20700
rect 12533 20644 12537 20700
rect 12473 20640 12537 20644
rect 12553 20700 12617 20704
rect 12553 20644 12557 20700
rect 12557 20644 12613 20700
rect 12613 20644 12617 20700
rect 12553 20640 12617 20644
rect 17994 20700 18058 20704
rect 17994 20644 17998 20700
rect 17998 20644 18054 20700
rect 18054 20644 18058 20700
rect 17994 20640 18058 20644
rect 18074 20700 18138 20704
rect 18074 20644 18078 20700
rect 18078 20644 18134 20700
rect 18134 20644 18138 20700
rect 18074 20640 18138 20644
rect 18154 20700 18218 20704
rect 18154 20644 18158 20700
rect 18158 20644 18214 20700
rect 18214 20644 18218 20700
rect 18154 20640 18218 20644
rect 18234 20700 18298 20704
rect 18234 20644 18238 20700
rect 18238 20644 18294 20700
rect 18294 20644 18298 20700
rect 18234 20640 18298 20644
rect 23675 20700 23739 20704
rect 23675 20644 23679 20700
rect 23679 20644 23735 20700
rect 23735 20644 23739 20700
rect 23675 20640 23739 20644
rect 23755 20700 23819 20704
rect 23755 20644 23759 20700
rect 23759 20644 23815 20700
rect 23815 20644 23819 20700
rect 23755 20640 23819 20644
rect 23835 20700 23899 20704
rect 23835 20644 23839 20700
rect 23839 20644 23895 20700
rect 23895 20644 23899 20700
rect 23835 20640 23899 20644
rect 23915 20700 23979 20704
rect 23915 20644 23919 20700
rect 23919 20644 23975 20700
rect 23975 20644 23979 20700
rect 23915 20640 23979 20644
rect 3792 20156 3856 20160
rect 3792 20100 3796 20156
rect 3796 20100 3852 20156
rect 3852 20100 3856 20156
rect 3792 20096 3856 20100
rect 3872 20156 3936 20160
rect 3872 20100 3876 20156
rect 3876 20100 3932 20156
rect 3932 20100 3936 20156
rect 3872 20096 3936 20100
rect 3952 20156 4016 20160
rect 3952 20100 3956 20156
rect 3956 20100 4012 20156
rect 4012 20100 4016 20156
rect 3952 20096 4016 20100
rect 4032 20156 4096 20160
rect 4032 20100 4036 20156
rect 4036 20100 4092 20156
rect 4092 20100 4096 20156
rect 4032 20096 4096 20100
rect 9473 20156 9537 20160
rect 9473 20100 9477 20156
rect 9477 20100 9533 20156
rect 9533 20100 9537 20156
rect 9473 20096 9537 20100
rect 9553 20156 9617 20160
rect 9553 20100 9557 20156
rect 9557 20100 9613 20156
rect 9613 20100 9617 20156
rect 9553 20096 9617 20100
rect 9633 20156 9697 20160
rect 9633 20100 9637 20156
rect 9637 20100 9693 20156
rect 9693 20100 9697 20156
rect 9633 20096 9697 20100
rect 9713 20156 9777 20160
rect 9713 20100 9717 20156
rect 9717 20100 9773 20156
rect 9773 20100 9777 20156
rect 9713 20096 9777 20100
rect 15154 20156 15218 20160
rect 15154 20100 15158 20156
rect 15158 20100 15214 20156
rect 15214 20100 15218 20156
rect 15154 20096 15218 20100
rect 15234 20156 15298 20160
rect 15234 20100 15238 20156
rect 15238 20100 15294 20156
rect 15294 20100 15298 20156
rect 15234 20096 15298 20100
rect 15314 20156 15378 20160
rect 15314 20100 15318 20156
rect 15318 20100 15374 20156
rect 15374 20100 15378 20156
rect 15314 20096 15378 20100
rect 15394 20156 15458 20160
rect 15394 20100 15398 20156
rect 15398 20100 15454 20156
rect 15454 20100 15458 20156
rect 15394 20096 15458 20100
rect 20835 20156 20899 20160
rect 20835 20100 20839 20156
rect 20839 20100 20895 20156
rect 20895 20100 20899 20156
rect 20835 20096 20899 20100
rect 20915 20156 20979 20160
rect 20915 20100 20919 20156
rect 20919 20100 20975 20156
rect 20975 20100 20979 20156
rect 20915 20096 20979 20100
rect 20995 20156 21059 20160
rect 20995 20100 20999 20156
rect 20999 20100 21055 20156
rect 21055 20100 21059 20156
rect 20995 20096 21059 20100
rect 21075 20156 21139 20160
rect 21075 20100 21079 20156
rect 21079 20100 21135 20156
rect 21135 20100 21139 20156
rect 21075 20096 21139 20100
rect 6632 19612 6696 19616
rect 6632 19556 6636 19612
rect 6636 19556 6692 19612
rect 6692 19556 6696 19612
rect 6632 19552 6696 19556
rect 6712 19612 6776 19616
rect 6712 19556 6716 19612
rect 6716 19556 6772 19612
rect 6772 19556 6776 19612
rect 6712 19552 6776 19556
rect 6792 19612 6856 19616
rect 6792 19556 6796 19612
rect 6796 19556 6852 19612
rect 6852 19556 6856 19612
rect 6792 19552 6856 19556
rect 6872 19612 6936 19616
rect 6872 19556 6876 19612
rect 6876 19556 6932 19612
rect 6932 19556 6936 19612
rect 6872 19552 6936 19556
rect 12313 19612 12377 19616
rect 12313 19556 12317 19612
rect 12317 19556 12373 19612
rect 12373 19556 12377 19612
rect 12313 19552 12377 19556
rect 12393 19612 12457 19616
rect 12393 19556 12397 19612
rect 12397 19556 12453 19612
rect 12453 19556 12457 19612
rect 12393 19552 12457 19556
rect 12473 19612 12537 19616
rect 12473 19556 12477 19612
rect 12477 19556 12533 19612
rect 12533 19556 12537 19612
rect 12473 19552 12537 19556
rect 12553 19612 12617 19616
rect 12553 19556 12557 19612
rect 12557 19556 12613 19612
rect 12613 19556 12617 19612
rect 12553 19552 12617 19556
rect 17994 19612 18058 19616
rect 17994 19556 17998 19612
rect 17998 19556 18054 19612
rect 18054 19556 18058 19612
rect 17994 19552 18058 19556
rect 18074 19612 18138 19616
rect 18074 19556 18078 19612
rect 18078 19556 18134 19612
rect 18134 19556 18138 19612
rect 18074 19552 18138 19556
rect 18154 19612 18218 19616
rect 18154 19556 18158 19612
rect 18158 19556 18214 19612
rect 18214 19556 18218 19612
rect 18154 19552 18218 19556
rect 18234 19612 18298 19616
rect 18234 19556 18238 19612
rect 18238 19556 18294 19612
rect 18294 19556 18298 19612
rect 18234 19552 18298 19556
rect 23675 19612 23739 19616
rect 23675 19556 23679 19612
rect 23679 19556 23735 19612
rect 23735 19556 23739 19612
rect 23675 19552 23739 19556
rect 23755 19612 23819 19616
rect 23755 19556 23759 19612
rect 23759 19556 23815 19612
rect 23815 19556 23819 19612
rect 23755 19552 23819 19556
rect 23835 19612 23899 19616
rect 23835 19556 23839 19612
rect 23839 19556 23895 19612
rect 23895 19556 23899 19612
rect 23835 19552 23899 19556
rect 23915 19612 23979 19616
rect 23915 19556 23919 19612
rect 23919 19556 23975 19612
rect 23975 19556 23979 19612
rect 23915 19552 23979 19556
rect 5396 19408 5460 19412
rect 5396 19352 5410 19408
rect 5410 19352 5460 19408
rect 5396 19348 5460 19352
rect 3792 19068 3856 19072
rect 3792 19012 3796 19068
rect 3796 19012 3852 19068
rect 3852 19012 3856 19068
rect 3792 19008 3856 19012
rect 3872 19068 3936 19072
rect 3872 19012 3876 19068
rect 3876 19012 3932 19068
rect 3932 19012 3936 19068
rect 3872 19008 3936 19012
rect 3952 19068 4016 19072
rect 3952 19012 3956 19068
rect 3956 19012 4012 19068
rect 4012 19012 4016 19068
rect 3952 19008 4016 19012
rect 4032 19068 4096 19072
rect 4032 19012 4036 19068
rect 4036 19012 4092 19068
rect 4092 19012 4096 19068
rect 4032 19008 4096 19012
rect 9473 19068 9537 19072
rect 9473 19012 9477 19068
rect 9477 19012 9533 19068
rect 9533 19012 9537 19068
rect 9473 19008 9537 19012
rect 9553 19068 9617 19072
rect 9553 19012 9557 19068
rect 9557 19012 9613 19068
rect 9613 19012 9617 19068
rect 9553 19008 9617 19012
rect 9633 19068 9697 19072
rect 9633 19012 9637 19068
rect 9637 19012 9693 19068
rect 9693 19012 9697 19068
rect 9633 19008 9697 19012
rect 9713 19068 9777 19072
rect 9713 19012 9717 19068
rect 9717 19012 9773 19068
rect 9773 19012 9777 19068
rect 9713 19008 9777 19012
rect 15154 19068 15218 19072
rect 15154 19012 15158 19068
rect 15158 19012 15214 19068
rect 15214 19012 15218 19068
rect 15154 19008 15218 19012
rect 15234 19068 15298 19072
rect 15234 19012 15238 19068
rect 15238 19012 15294 19068
rect 15294 19012 15298 19068
rect 15234 19008 15298 19012
rect 15314 19068 15378 19072
rect 15314 19012 15318 19068
rect 15318 19012 15374 19068
rect 15374 19012 15378 19068
rect 15314 19008 15378 19012
rect 15394 19068 15458 19072
rect 15394 19012 15398 19068
rect 15398 19012 15454 19068
rect 15454 19012 15458 19068
rect 15394 19008 15458 19012
rect 20835 19068 20899 19072
rect 20835 19012 20839 19068
rect 20839 19012 20895 19068
rect 20895 19012 20899 19068
rect 20835 19008 20899 19012
rect 20915 19068 20979 19072
rect 20915 19012 20919 19068
rect 20919 19012 20975 19068
rect 20975 19012 20979 19068
rect 20915 19008 20979 19012
rect 20995 19068 21059 19072
rect 20995 19012 20999 19068
rect 20999 19012 21055 19068
rect 21055 19012 21059 19068
rect 20995 19008 21059 19012
rect 21075 19068 21139 19072
rect 21075 19012 21079 19068
rect 21079 19012 21135 19068
rect 21135 19012 21139 19068
rect 21075 19008 21139 19012
rect 14964 18804 15028 18868
rect 6632 18524 6696 18528
rect 6632 18468 6636 18524
rect 6636 18468 6692 18524
rect 6692 18468 6696 18524
rect 6632 18464 6696 18468
rect 6712 18524 6776 18528
rect 6712 18468 6716 18524
rect 6716 18468 6772 18524
rect 6772 18468 6776 18524
rect 6712 18464 6776 18468
rect 6792 18524 6856 18528
rect 6792 18468 6796 18524
rect 6796 18468 6852 18524
rect 6852 18468 6856 18524
rect 6792 18464 6856 18468
rect 6872 18524 6936 18528
rect 6872 18468 6876 18524
rect 6876 18468 6932 18524
rect 6932 18468 6936 18524
rect 6872 18464 6936 18468
rect 12313 18524 12377 18528
rect 12313 18468 12317 18524
rect 12317 18468 12373 18524
rect 12373 18468 12377 18524
rect 12313 18464 12377 18468
rect 12393 18524 12457 18528
rect 12393 18468 12397 18524
rect 12397 18468 12453 18524
rect 12453 18468 12457 18524
rect 12393 18464 12457 18468
rect 12473 18524 12537 18528
rect 12473 18468 12477 18524
rect 12477 18468 12533 18524
rect 12533 18468 12537 18524
rect 12473 18464 12537 18468
rect 12553 18524 12617 18528
rect 12553 18468 12557 18524
rect 12557 18468 12613 18524
rect 12613 18468 12617 18524
rect 12553 18464 12617 18468
rect 17994 18524 18058 18528
rect 17994 18468 17998 18524
rect 17998 18468 18054 18524
rect 18054 18468 18058 18524
rect 17994 18464 18058 18468
rect 18074 18524 18138 18528
rect 18074 18468 18078 18524
rect 18078 18468 18134 18524
rect 18134 18468 18138 18524
rect 18074 18464 18138 18468
rect 18154 18524 18218 18528
rect 18154 18468 18158 18524
rect 18158 18468 18214 18524
rect 18214 18468 18218 18524
rect 18154 18464 18218 18468
rect 18234 18524 18298 18528
rect 18234 18468 18238 18524
rect 18238 18468 18294 18524
rect 18294 18468 18298 18524
rect 18234 18464 18298 18468
rect 23675 18524 23739 18528
rect 23675 18468 23679 18524
rect 23679 18468 23735 18524
rect 23735 18468 23739 18524
rect 23675 18464 23739 18468
rect 23755 18524 23819 18528
rect 23755 18468 23759 18524
rect 23759 18468 23815 18524
rect 23815 18468 23819 18524
rect 23755 18464 23819 18468
rect 23835 18524 23899 18528
rect 23835 18468 23839 18524
rect 23839 18468 23895 18524
rect 23895 18468 23899 18524
rect 23835 18464 23899 18468
rect 23915 18524 23979 18528
rect 23915 18468 23919 18524
rect 23919 18468 23975 18524
rect 23975 18468 23979 18524
rect 23915 18464 23979 18468
rect 19932 18048 19996 18052
rect 19932 17992 19946 18048
rect 19946 17992 19996 18048
rect 19932 17988 19996 17992
rect 3792 17980 3856 17984
rect 3792 17924 3796 17980
rect 3796 17924 3852 17980
rect 3852 17924 3856 17980
rect 3792 17920 3856 17924
rect 3872 17980 3936 17984
rect 3872 17924 3876 17980
rect 3876 17924 3932 17980
rect 3932 17924 3936 17980
rect 3872 17920 3936 17924
rect 3952 17980 4016 17984
rect 3952 17924 3956 17980
rect 3956 17924 4012 17980
rect 4012 17924 4016 17980
rect 3952 17920 4016 17924
rect 4032 17980 4096 17984
rect 4032 17924 4036 17980
rect 4036 17924 4092 17980
rect 4092 17924 4096 17980
rect 4032 17920 4096 17924
rect 9473 17980 9537 17984
rect 9473 17924 9477 17980
rect 9477 17924 9533 17980
rect 9533 17924 9537 17980
rect 9473 17920 9537 17924
rect 9553 17980 9617 17984
rect 9553 17924 9557 17980
rect 9557 17924 9613 17980
rect 9613 17924 9617 17980
rect 9553 17920 9617 17924
rect 9633 17980 9697 17984
rect 9633 17924 9637 17980
rect 9637 17924 9693 17980
rect 9693 17924 9697 17980
rect 9633 17920 9697 17924
rect 9713 17980 9777 17984
rect 9713 17924 9717 17980
rect 9717 17924 9773 17980
rect 9773 17924 9777 17980
rect 9713 17920 9777 17924
rect 15154 17980 15218 17984
rect 15154 17924 15158 17980
rect 15158 17924 15214 17980
rect 15214 17924 15218 17980
rect 15154 17920 15218 17924
rect 15234 17980 15298 17984
rect 15234 17924 15238 17980
rect 15238 17924 15294 17980
rect 15294 17924 15298 17980
rect 15234 17920 15298 17924
rect 15314 17980 15378 17984
rect 15314 17924 15318 17980
rect 15318 17924 15374 17980
rect 15374 17924 15378 17980
rect 15314 17920 15378 17924
rect 15394 17980 15458 17984
rect 15394 17924 15398 17980
rect 15398 17924 15454 17980
rect 15454 17924 15458 17980
rect 15394 17920 15458 17924
rect 20835 17980 20899 17984
rect 20835 17924 20839 17980
rect 20839 17924 20895 17980
rect 20895 17924 20899 17980
rect 20835 17920 20899 17924
rect 20915 17980 20979 17984
rect 20915 17924 20919 17980
rect 20919 17924 20975 17980
rect 20975 17924 20979 17980
rect 20915 17920 20979 17924
rect 20995 17980 21059 17984
rect 20995 17924 20999 17980
rect 20999 17924 21055 17980
rect 21055 17924 21059 17980
rect 20995 17920 21059 17924
rect 21075 17980 21139 17984
rect 21075 17924 21079 17980
rect 21079 17924 21135 17980
rect 21135 17924 21139 17980
rect 21075 17920 21139 17924
rect 6632 17436 6696 17440
rect 6632 17380 6636 17436
rect 6636 17380 6692 17436
rect 6692 17380 6696 17436
rect 6632 17376 6696 17380
rect 6712 17436 6776 17440
rect 6712 17380 6716 17436
rect 6716 17380 6772 17436
rect 6772 17380 6776 17436
rect 6712 17376 6776 17380
rect 6792 17436 6856 17440
rect 6792 17380 6796 17436
rect 6796 17380 6852 17436
rect 6852 17380 6856 17436
rect 6792 17376 6856 17380
rect 6872 17436 6936 17440
rect 6872 17380 6876 17436
rect 6876 17380 6932 17436
rect 6932 17380 6936 17436
rect 6872 17376 6936 17380
rect 12313 17436 12377 17440
rect 12313 17380 12317 17436
rect 12317 17380 12373 17436
rect 12373 17380 12377 17436
rect 12313 17376 12377 17380
rect 12393 17436 12457 17440
rect 12393 17380 12397 17436
rect 12397 17380 12453 17436
rect 12453 17380 12457 17436
rect 12393 17376 12457 17380
rect 12473 17436 12537 17440
rect 12473 17380 12477 17436
rect 12477 17380 12533 17436
rect 12533 17380 12537 17436
rect 12473 17376 12537 17380
rect 12553 17436 12617 17440
rect 12553 17380 12557 17436
rect 12557 17380 12613 17436
rect 12613 17380 12617 17436
rect 12553 17376 12617 17380
rect 17994 17436 18058 17440
rect 17994 17380 17998 17436
rect 17998 17380 18054 17436
rect 18054 17380 18058 17436
rect 17994 17376 18058 17380
rect 18074 17436 18138 17440
rect 18074 17380 18078 17436
rect 18078 17380 18134 17436
rect 18134 17380 18138 17436
rect 18074 17376 18138 17380
rect 18154 17436 18218 17440
rect 18154 17380 18158 17436
rect 18158 17380 18214 17436
rect 18214 17380 18218 17436
rect 18154 17376 18218 17380
rect 18234 17436 18298 17440
rect 18234 17380 18238 17436
rect 18238 17380 18294 17436
rect 18294 17380 18298 17436
rect 18234 17376 18298 17380
rect 23675 17436 23739 17440
rect 23675 17380 23679 17436
rect 23679 17380 23735 17436
rect 23735 17380 23739 17436
rect 23675 17376 23739 17380
rect 23755 17436 23819 17440
rect 23755 17380 23759 17436
rect 23759 17380 23815 17436
rect 23815 17380 23819 17436
rect 23755 17376 23819 17380
rect 23835 17436 23899 17440
rect 23835 17380 23839 17436
rect 23839 17380 23895 17436
rect 23895 17380 23899 17436
rect 23835 17376 23899 17380
rect 23915 17436 23979 17440
rect 23915 17380 23919 17436
rect 23919 17380 23975 17436
rect 23975 17380 23979 17436
rect 23915 17376 23979 17380
rect 3792 16892 3856 16896
rect 3792 16836 3796 16892
rect 3796 16836 3852 16892
rect 3852 16836 3856 16892
rect 3792 16832 3856 16836
rect 3872 16892 3936 16896
rect 3872 16836 3876 16892
rect 3876 16836 3932 16892
rect 3932 16836 3936 16892
rect 3872 16832 3936 16836
rect 3952 16892 4016 16896
rect 3952 16836 3956 16892
rect 3956 16836 4012 16892
rect 4012 16836 4016 16892
rect 3952 16832 4016 16836
rect 4032 16892 4096 16896
rect 4032 16836 4036 16892
rect 4036 16836 4092 16892
rect 4092 16836 4096 16892
rect 4032 16832 4096 16836
rect 9473 16892 9537 16896
rect 9473 16836 9477 16892
rect 9477 16836 9533 16892
rect 9533 16836 9537 16892
rect 9473 16832 9537 16836
rect 9553 16892 9617 16896
rect 9553 16836 9557 16892
rect 9557 16836 9613 16892
rect 9613 16836 9617 16892
rect 9553 16832 9617 16836
rect 9633 16892 9697 16896
rect 9633 16836 9637 16892
rect 9637 16836 9693 16892
rect 9693 16836 9697 16892
rect 9633 16832 9697 16836
rect 9713 16892 9777 16896
rect 9713 16836 9717 16892
rect 9717 16836 9773 16892
rect 9773 16836 9777 16892
rect 9713 16832 9777 16836
rect 15154 16892 15218 16896
rect 15154 16836 15158 16892
rect 15158 16836 15214 16892
rect 15214 16836 15218 16892
rect 15154 16832 15218 16836
rect 15234 16892 15298 16896
rect 15234 16836 15238 16892
rect 15238 16836 15294 16892
rect 15294 16836 15298 16892
rect 15234 16832 15298 16836
rect 15314 16892 15378 16896
rect 15314 16836 15318 16892
rect 15318 16836 15374 16892
rect 15374 16836 15378 16892
rect 15314 16832 15378 16836
rect 15394 16892 15458 16896
rect 15394 16836 15398 16892
rect 15398 16836 15454 16892
rect 15454 16836 15458 16892
rect 15394 16832 15458 16836
rect 20835 16892 20899 16896
rect 20835 16836 20839 16892
rect 20839 16836 20895 16892
rect 20895 16836 20899 16892
rect 20835 16832 20899 16836
rect 20915 16892 20979 16896
rect 20915 16836 20919 16892
rect 20919 16836 20975 16892
rect 20975 16836 20979 16892
rect 20915 16832 20979 16836
rect 20995 16892 21059 16896
rect 20995 16836 20999 16892
rect 20999 16836 21055 16892
rect 21055 16836 21059 16892
rect 20995 16832 21059 16836
rect 21075 16892 21139 16896
rect 21075 16836 21079 16892
rect 21079 16836 21135 16892
rect 21135 16836 21139 16892
rect 21075 16832 21139 16836
rect 6316 16628 6380 16692
rect 6632 16348 6696 16352
rect 6632 16292 6636 16348
rect 6636 16292 6692 16348
rect 6692 16292 6696 16348
rect 6632 16288 6696 16292
rect 6712 16348 6776 16352
rect 6712 16292 6716 16348
rect 6716 16292 6772 16348
rect 6772 16292 6776 16348
rect 6712 16288 6776 16292
rect 6792 16348 6856 16352
rect 6792 16292 6796 16348
rect 6796 16292 6852 16348
rect 6852 16292 6856 16348
rect 6792 16288 6856 16292
rect 6872 16348 6936 16352
rect 6872 16292 6876 16348
rect 6876 16292 6932 16348
rect 6932 16292 6936 16348
rect 6872 16288 6936 16292
rect 12313 16348 12377 16352
rect 12313 16292 12317 16348
rect 12317 16292 12373 16348
rect 12373 16292 12377 16348
rect 12313 16288 12377 16292
rect 12393 16348 12457 16352
rect 12393 16292 12397 16348
rect 12397 16292 12453 16348
rect 12453 16292 12457 16348
rect 12393 16288 12457 16292
rect 12473 16348 12537 16352
rect 12473 16292 12477 16348
rect 12477 16292 12533 16348
rect 12533 16292 12537 16348
rect 12473 16288 12537 16292
rect 12553 16348 12617 16352
rect 12553 16292 12557 16348
rect 12557 16292 12613 16348
rect 12613 16292 12617 16348
rect 12553 16288 12617 16292
rect 17994 16348 18058 16352
rect 17994 16292 17998 16348
rect 17998 16292 18054 16348
rect 18054 16292 18058 16348
rect 17994 16288 18058 16292
rect 18074 16348 18138 16352
rect 18074 16292 18078 16348
rect 18078 16292 18134 16348
rect 18134 16292 18138 16348
rect 18074 16288 18138 16292
rect 18154 16348 18218 16352
rect 18154 16292 18158 16348
rect 18158 16292 18214 16348
rect 18214 16292 18218 16348
rect 18154 16288 18218 16292
rect 18234 16348 18298 16352
rect 18234 16292 18238 16348
rect 18238 16292 18294 16348
rect 18294 16292 18298 16348
rect 18234 16288 18298 16292
rect 23675 16348 23739 16352
rect 23675 16292 23679 16348
rect 23679 16292 23735 16348
rect 23735 16292 23739 16348
rect 23675 16288 23739 16292
rect 23755 16348 23819 16352
rect 23755 16292 23759 16348
rect 23759 16292 23815 16348
rect 23815 16292 23819 16348
rect 23755 16288 23819 16292
rect 23835 16348 23899 16352
rect 23835 16292 23839 16348
rect 23839 16292 23895 16348
rect 23895 16292 23899 16348
rect 23835 16288 23899 16292
rect 23915 16348 23979 16352
rect 23915 16292 23919 16348
rect 23919 16292 23975 16348
rect 23975 16292 23979 16348
rect 23915 16288 23979 16292
rect 3792 15804 3856 15808
rect 3792 15748 3796 15804
rect 3796 15748 3852 15804
rect 3852 15748 3856 15804
rect 3792 15744 3856 15748
rect 3872 15804 3936 15808
rect 3872 15748 3876 15804
rect 3876 15748 3932 15804
rect 3932 15748 3936 15804
rect 3872 15744 3936 15748
rect 3952 15804 4016 15808
rect 3952 15748 3956 15804
rect 3956 15748 4012 15804
rect 4012 15748 4016 15804
rect 3952 15744 4016 15748
rect 4032 15804 4096 15808
rect 4032 15748 4036 15804
rect 4036 15748 4092 15804
rect 4092 15748 4096 15804
rect 4032 15744 4096 15748
rect 9473 15804 9537 15808
rect 9473 15748 9477 15804
rect 9477 15748 9533 15804
rect 9533 15748 9537 15804
rect 9473 15744 9537 15748
rect 9553 15804 9617 15808
rect 9553 15748 9557 15804
rect 9557 15748 9613 15804
rect 9613 15748 9617 15804
rect 9553 15744 9617 15748
rect 9633 15804 9697 15808
rect 9633 15748 9637 15804
rect 9637 15748 9693 15804
rect 9693 15748 9697 15804
rect 9633 15744 9697 15748
rect 9713 15804 9777 15808
rect 9713 15748 9717 15804
rect 9717 15748 9773 15804
rect 9773 15748 9777 15804
rect 9713 15744 9777 15748
rect 15154 15804 15218 15808
rect 15154 15748 15158 15804
rect 15158 15748 15214 15804
rect 15214 15748 15218 15804
rect 15154 15744 15218 15748
rect 15234 15804 15298 15808
rect 15234 15748 15238 15804
rect 15238 15748 15294 15804
rect 15294 15748 15298 15804
rect 15234 15744 15298 15748
rect 15314 15804 15378 15808
rect 15314 15748 15318 15804
rect 15318 15748 15374 15804
rect 15374 15748 15378 15804
rect 15314 15744 15378 15748
rect 15394 15804 15458 15808
rect 15394 15748 15398 15804
rect 15398 15748 15454 15804
rect 15454 15748 15458 15804
rect 15394 15744 15458 15748
rect 20835 15804 20899 15808
rect 20835 15748 20839 15804
rect 20839 15748 20895 15804
rect 20895 15748 20899 15804
rect 20835 15744 20899 15748
rect 20915 15804 20979 15808
rect 20915 15748 20919 15804
rect 20919 15748 20975 15804
rect 20975 15748 20979 15804
rect 20915 15744 20979 15748
rect 20995 15804 21059 15808
rect 20995 15748 20999 15804
rect 20999 15748 21055 15804
rect 21055 15748 21059 15804
rect 20995 15744 21059 15748
rect 21075 15804 21139 15808
rect 21075 15748 21079 15804
rect 21079 15748 21135 15804
rect 21135 15748 21139 15804
rect 21075 15744 21139 15748
rect 6632 15260 6696 15264
rect 6632 15204 6636 15260
rect 6636 15204 6692 15260
rect 6692 15204 6696 15260
rect 6632 15200 6696 15204
rect 6712 15260 6776 15264
rect 6712 15204 6716 15260
rect 6716 15204 6772 15260
rect 6772 15204 6776 15260
rect 6712 15200 6776 15204
rect 6792 15260 6856 15264
rect 6792 15204 6796 15260
rect 6796 15204 6852 15260
rect 6852 15204 6856 15260
rect 6792 15200 6856 15204
rect 6872 15260 6936 15264
rect 6872 15204 6876 15260
rect 6876 15204 6932 15260
rect 6932 15204 6936 15260
rect 6872 15200 6936 15204
rect 12313 15260 12377 15264
rect 12313 15204 12317 15260
rect 12317 15204 12373 15260
rect 12373 15204 12377 15260
rect 12313 15200 12377 15204
rect 12393 15260 12457 15264
rect 12393 15204 12397 15260
rect 12397 15204 12453 15260
rect 12453 15204 12457 15260
rect 12393 15200 12457 15204
rect 12473 15260 12537 15264
rect 12473 15204 12477 15260
rect 12477 15204 12533 15260
rect 12533 15204 12537 15260
rect 12473 15200 12537 15204
rect 12553 15260 12617 15264
rect 12553 15204 12557 15260
rect 12557 15204 12613 15260
rect 12613 15204 12617 15260
rect 12553 15200 12617 15204
rect 17994 15260 18058 15264
rect 17994 15204 17998 15260
rect 17998 15204 18054 15260
rect 18054 15204 18058 15260
rect 17994 15200 18058 15204
rect 18074 15260 18138 15264
rect 18074 15204 18078 15260
rect 18078 15204 18134 15260
rect 18134 15204 18138 15260
rect 18074 15200 18138 15204
rect 18154 15260 18218 15264
rect 18154 15204 18158 15260
rect 18158 15204 18214 15260
rect 18214 15204 18218 15260
rect 18154 15200 18218 15204
rect 18234 15260 18298 15264
rect 18234 15204 18238 15260
rect 18238 15204 18294 15260
rect 18294 15204 18298 15260
rect 18234 15200 18298 15204
rect 23675 15260 23739 15264
rect 23675 15204 23679 15260
rect 23679 15204 23735 15260
rect 23735 15204 23739 15260
rect 23675 15200 23739 15204
rect 23755 15260 23819 15264
rect 23755 15204 23759 15260
rect 23759 15204 23815 15260
rect 23815 15204 23819 15260
rect 23755 15200 23819 15204
rect 23835 15260 23899 15264
rect 23835 15204 23839 15260
rect 23839 15204 23895 15260
rect 23895 15204 23899 15260
rect 23835 15200 23899 15204
rect 23915 15260 23979 15264
rect 23915 15204 23919 15260
rect 23919 15204 23975 15260
rect 23975 15204 23979 15260
rect 23915 15200 23979 15204
rect 14228 15132 14292 15196
rect 3792 14716 3856 14720
rect 3792 14660 3796 14716
rect 3796 14660 3852 14716
rect 3852 14660 3856 14716
rect 3792 14656 3856 14660
rect 3872 14716 3936 14720
rect 3872 14660 3876 14716
rect 3876 14660 3932 14716
rect 3932 14660 3936 14716
rect 3872 14656 3936 14660
rect 3952 14716 4016 14720
rect 3952 14660 3956 14716
rect 3956 14660 4012 14716
rect 4012 14660 4016 14716
rect 3952 14656 4016 14660
rect 4032 14716 4096 14720
rect 4032 14660 4036 14716
rect 4036 14660 4092 14716
rect 4092 14660 4096 14716
rect 4032 14656 4096 14660
rect 9473 14716 9537 14720
rect 9473 14660 9477 14716
rect 9477 14660 9533 14716
rect 9533 14660 9537 14716
rect 9473 14656 9537 14660
rect 9553 14716 9617 14720
rect 9553 14660 9557 14716
rect 9557 14660 9613 14716
rect 9613 14660 9617 14716
rect 9553 14656 9617 14660
rect 9633 14716 9697 14720
rect 9633 14660 9637 14716
rect 9637 14660 9693 14716
rect 9693 14660 9697 14716
rect 9633 14656 9697 14660
rect 9713 14716 9777 14720
rect 9713 14660 9717 14716
rect 9717 14660 9773 14716
rect 9773 14660 9777 14716
rect 9713 14656 9777 14660
rect 15154 14716 15218 14720
rect 15154 14660 15158 14716
rect 15158 14660 15214 14716
rect 15214 14660 15218 14716
rect 15154 14656 15218 14660
rect 15234 14716 15298 14720
rect 15234 14660 15238 14716
rect 15238 14660 15294 14716
rect 15294 14660 15298 14716
rect 15234 14656 15298 14660
rect 15314 14716 15378 14720
rect 15314 14660 15318 14716
rect 15318 14660 15374 14716
rect 15374 14660 15378 14716
rect 15314 14656 15378 14660
rect 15394 14716 15458 14720
rect 15394 14660 15398 14716
rect 15398 14660 15454 14716
rect 15454 14660 15458 14716
rect 15394 14656 15458 14660
rect 20835 14716 20899 14720
rect 20835 14660 20839 14716
rect 20839 14660 20895 14716
rect 20895 14660 20899 14716
rect 20835 14656 20899 14660
rect 20915 14716 20979 14720
rect 20915 14660 20919 14716
rect 20919 14660 20975 14716
rect 20975 14660 20979 14716
rect 20915 14656 20979 14660
rect 20995 14716 21059 14720
rect 20995 14660 20999 14716
rect 20999 14660 21055 14716
rect 21055 14660 21059 14716
rect 20995 14656 21059 14660
rect 21075 14716 21139 14720
rect 21075 14660 21079 14716
rect 21079 14660 21135 14716
rect 21135 14660 21139 14716
rect 21075 14656 21139 14660
rect 6632 14172 6696 14176
rect 6632 14116 6636 14172
rect 6636 14116 6692 14172
rect 6692 14116 6696 14172
rect 6632 14112 6696 14116
rect 6712 14172 6776 14176
rect 6712 14116 6716 14172
rect 6716 14116 6772 14172
rect 6772 14116 6776 14172
rect 6712 14112 6776 14116
rect 6792 14172 6856 14176
rect 6792 14116 6796 14172
rect 6796 14116 6852 14172
rect 6852 14116 6856 14172
rect 6792 14112 6856 14116
rect 6872 14172 6936 14176
rect 6872 14116 6876 14172
rect 6876 14116 6932 14172
rect 6932 14116 6936 14172
rect 6872 14112 6936 14116
rect 12313 14172 12377 14176
rect 12313 14116 12317 14172
rect 12317 14116 12373 14172
rect 12373 14116 12377 14172
rect 12313 14112 12377 14116
rect 12393 14172 12457 14176
rect 12393 14116 12397 14172
rect 12397 14116 12453 14172
rect 12453 14116 12457 14172
rect 12393 14112 12457 14116
rect 12473 14172 12537 14176
rect 12473 14116 12477 14172
rect 12477 14116 12533 14172
rect 12533 14116 12537 14172
rect 12473 14112 12537 14116
rect 12553 14172 12617 14176
rect 12553 14116 12557 14172
rect 12557 14116 12613 14172
rect 12613 14116 12617 14172
rect 12553 14112 12617 14116
rect 17994 14172 18058 14176
rect 17994 14116 17998 14172
rect 17998 14116 18054 14172
rect 18054 14116 18058 14172
rect 17994 14112 18058 14116
rect 18074 14172 18138 14176
rect 18074 14116 18078 14172
rect 18078 14116 18134 14172
rect 18134 14116 18138 14172
rect 18074 14112 18138 14116
rect 18154 14172 18218 14176
rect 18154 14116 18158 14172
rect 18158 14116 18214 14172
rect 18214 14116 18218 14172
rect 18154 14112 18218 14116
rect 18234 14172 18298 14176
rect 18234 14116 18238 14172
rect 18238 14116 18294 14172
rect 18294 14116 18298 14172
rect 18234 14112 18298 14116
rect 23675 14172 23739 14176
rect 23675 14116 23679 14172
rect 23679 14116 23735 14172
rect 23735 14116 23739 14172
rect 23675 14112 23739 14116
rect 23755 14172 23819 14176
rect 23755 14116 23759 14172
rect 23759 14116 23815 14172
rect 23815 14116 23819 14172
rect 23755 14112 23819 14116
rect 23835 14172 23899 14176
rect 23835 14116 23839 14172
rect 23839 14116 23895 14172
rect 23895 14116 23899 14172
rect 23835 14112 23899 14116
rect 23915 14172 23979 14176
rect 23915 14116 23919 14172
rect 23919 14116 23975 14172
rect 23975 14116 23979 14172
rect 23915 14112 23979 14116
rect 14596 13772 14660 13836
rect 14964 13772 15028 13836
rect 3792 13628 3856 13632
rect 3792 13572 3796 13628
rect 3796 13572 3852 13628
rect 3852 13572 3856 13628
rect 3792 13568 3856 13572
rect 3872 13628 3936 13632
rect 3872 13572 3876 13628
rect 3876 13572 3932 13628
rect 3932 13572 3936 13628
rect 3872 13568 3936 13572
rect 3952 13628 4016 13632
rect 3952 13572 3956 13628
rect 3956 13572 4012 13628
rect 4012 13572 4016 13628
rect 3952 13568 4016 13572
rect 4032 13628 4096 13632
rect 4032 13572 4036 13628
rect 4036 13572 4092 13628
rect 4092 13572 4096 13628
rect 4032 13568 4096 13572
rect 9473 13628 9537 13632
rect 9473 13572 9477 13628
rect 9477 13572 9533 13628
rect 9533 13572 9537 13628
rect 9473 13568 9537 13572
rect 9553 13628 9617 13632
rect 9553 13572 9557 13628
rect 9557 13572 9613 13628
rect 9613 13572 9617 13628
rect 9553 13568 9617 13572
rect 9633 13628 9697 13632
rect 9633 13572 9637 13628
rect 9637 13572 9693 13628
rect 9693 13572 9697 13628
rect 9633 13568 9697 13572
rect 9713 13628 9777 13632
rect 9713 13572 9717 13628
rect 9717 13572 9773 13628
rect 9773 13572 9777 13628
rect 9713 13568 9777 13572
rect 15154 13628 15218 13632
rect 15154 13572 15158 13628
rect 15158 13572 15214 13628
rect 15214 13572 15218 13628
rect 15154 13568 15218 13572
rect 15234 13628 15298 13632
rect 15234 13572 15238 13628
rect 15238 13572 15294 13628
rect 15294 13572 15298 13628
rect 15234 13568 15298 13572
rect 15314 13628 15378 13632
rect 15314 13572 15318 13628
rect 15318 13572 15374 13628
rect 15374 13572 15378 13628
rect 15314 13568 15378 13572
rect 15394 13628 15458 13632
rect 15394 13572 15398 13628
rect 15398 13572 15454 13628
rect 15454 13572 15458 13628
rect 15394 13568 15458 13572
rect 20835 13628 20899 13632
rect 20835 13572 20839 13628
rect 20839 13572 20895 13628
rect 20895 13572 20899 13628
rect 20835 13568 20899 13572
rect 20915 13628 20979 13632
rect 20915 13572 20919 13628
rect 20919 13572 20975 13628
rect 20975 13572 20979 13628
rect 20915 13568 20979 13572
rect 20995 13628 21059 13632
rect 20995 13572 20999 13628
rect 20999 13572 21055 13628
rect 21055 13572 21059 13628
rect 20995 13568 21059 13572
rect 21075 13628 21139 13632
rect 21075 13572 21079 13628
rect 21079 13572 21135 13628
rect 21135 13572 21139 13628
rect 21075 13568 21139 13572
rect 6632 13084 6696 13088
rect 6632 13028 6636 13084
rect 6636 13028 6692 13084
rect 6692 13028 6696 13084
rect 6632 13024 6696 13028
rect 6712 13084 6776 13088
rect 6712 13028 6716 13084
rect 6716 13028 6772 13084
rect 6772 13028 6776 13084
rect 6712 13024 6776 13028
rect 6792 13084 6856 13088
rect 6792 13028 6796 13084
rect 6796 13028 6852 13084
rect 6852 13028 6856 13084
rect 6792 13024 6856 13028
rect 6872 13084 6936 13088
rect 6872 13028 6876 13084
rect 6876 13028 6932 13084
rect 6932 13028 6936 13084
rect 6872 13024 6936 13028
rect 12313 13084 12377 13088
rect 12313 13028 12317 13084
rect 12317 13028 12373 13084
rect 12373 13028 12377 13084
rect 12313 13024 12377 13028
rect 12393 13084 12457 13088
rect 12393 13028 12397 13084
rect 12397 13028 12453 13084
rect 12453 13028 12457 13084
rect 12393 13024 12457 13028
rect 12473 13084 12537 13088
rect 12473 13028 12477 13084
rect 12477 13028 12533 13084
rect 12533 13028 12537 13084
rect 12473 13024 12537 13028
rect 12553 13084 12617 13088
rect 12553 13028 12557 13084
rect 12557 13028 12613 13084
rect 12613 13028 12617 13084
rect 12553 13024 12617 13028
rect 17994 13084 18058 13088
rect 17994 13028 17998 13084
rect 17998 13028 18054 13084
rect 18054 13028 18058 13084
rect 17994 13024 18058 13028
rect 18074 13084 18138 13088
rect 18074 13028 18078 13084
rect 18078 13028 18134 13084
rect 18134 13028 18138 13084
rect 18074 13024 18138 13028
rect 18154 13084 18218 13088
rect 18154 13028 18158 13084
rect 18158 13028 18214 13084
rect 18214 13028 18218 13084
rect 18154 13024 18218 13028
rect 18234 13084 18298 13088
rect 18234 13028 18238 13084
rect 18238 13028 18294 13084
rect 18294 13028 18298 13084
rect 18234 13024 18298 13028
rect 23675 13084 23739 13088
rect 23675 13028 23679 13084
rect 23679 13028 23735 13084
rect 23735 13028 23739 13084
rect 23675 13024 23739 13028
rect 23755 13084 23819 13088
rect 23755 13028 23759 13084
rect 23759 13028 23815 13084
rect 23815 13028 23819 13084
rect 23755 13024 23819 13028
rect 23835 13084 23899 13088
rect 23835 13028 23839 13084
rect 23839 13028 23895 13084
rect 23895 13028 23899 13084
rect 23835 13024 23899 13028
rect 23915 13084 23979 13088
rect 23915 13028 23919 13084
rect 23919 13028 23975 13084
rect 23975 13028 23979 13084
rect 23915 13024 23979 13028
rect 3792 12540 3856 12544
rect 3792 12484 3796 12540
rect 3796 12484 3852 12540
rect 3852 12484 3856 12540
rect 3792 12480 3856 12484
rect 3872 12540 3936 12544
rect 3872 12484 3876 12540
rect 3876 12484 3932 12540
rect 3932 12484 3936 12540
rect 3872 12480 3936 12484
rect 3952 12540 4016 12544
rect 3952 12484 3956 12540
rect 3956 12484 4012 12540
rect 4012 12484 4016 12540
rect 3952 12480 4016 12484
rect 4032 12540 4096 12544
rect 4032 12484 4036 12540
rect 4036 12484 4092 12540
rect 4092 12484 4096 12540
rect 4032 12480 4096 12484
rect 9473 12540 9537 12544
rect 9473 12484 9477 12540
rect 9477 12484 9533 12540
rect 9533 12484 9537 12540
rect 9473 12480 9537 12484
rect 9553 12540 9617 12544
rect 9553 12484 9557 12540
rect 9557 12484 9613 12540
rect 9613 12484 9617 12540
rect 9553 12480 9617 12484
rect 9633 12540 9697 12544
rect 9633 12484 9637 12540
rect 9637 12484 9693 12540
rect 9693 12484 9697 12540
rect 9633 12480 9697 12484
rect 9713 12540 9777 12544
rect 9713 12484 9717 12540
rect 9717 12484 9773 12540
rect 9773 12484 9777 12540
rect 9713 12480 9777 12484
rect 15154 12540 15218 12544
rect 15154 12484 15158 12540
rect 15158 12484 15214 12540
rect 15214 12484 15218 12540
rect 15154 12480 15218 12484
rect 15234 12540 15298 12544
rect 15234 12484 15238 12540
rect 15238 12484 15294 12540
rect 15294 12484 15298 12540
rect 15234 12480 15298 12484
rect 15314 12540 15378 12544
rect 15314 12484 15318 12540
rect 15318 12484 15374 12540
rect 15374 12484 15378 12540
rect 15314 12480 15378 12484
rect 15394 12540 15458 12544
rect 15394 12484 15398 12540
rect 15398 12484 15454 12540
rect 15454 12484 15458 12540
rect 15394 12480 15458 12484
rect 20835 12540 20899 12544
rect 20835 12484 20839 12540
rect 20839 12484 20895 12540
rect 20895 12484 20899 12540
rect 20835 12480 20899 12484
rect 20915 12540 20979 12544
rect 20915 12484 20919 12540
rect 20919 12484 20975 12540
rect 20975 12484 20979 12540
rect 20915 12480 20979 12484
rect 20995 12540 21059 12544
rect 20995 12484 20999 12540
rect 20999 12484 21055 12540
rect 21055 12484 21059 12540
rect 20995 12480 21059 12484
rect 21075 12540 21139 12544
rect 21075 12484 21079 12540
rect 21079 12484 21135 12540
rect 21135 12484 21139 12540
rect 21075 12480 21139 12484
rect 19748 12276 19812 12340
rect 5396 12064 5460 12068
rect 5396 12008 5446 12064
rect 5446 12008 5460 12064
rect 5396 12004 5460 12008
rect 6632 11996 6696 12000
rect 6632 11940 6636 11996
rect 6636 11940 6692 11996
rect 6692 11940 6696 11996
rect 6632 11936 6696 11940
rect 6712 11996 6776 12000
rect 6712 11940 6716 11996
rect 6716 11940 6772 11996
rect 6772 11940 6776 11996
rect 6712 11936 6776 11940
rect 6792 11996 6856 12000
rect 6792 11940 6796 11996
rect 6796 11940 6852 11996
rect 6852 11940 6856 11996
rect 6792 11936 6856 11940
rect 6872 11996 6936 12000
rect 6872 11940 6876 11996
rect 6876 11940 6932 11996
rect 6932 11940 6936 11996
rect 6872 11936 6936 11940
rect 12313 11996 12377 12000
rect 12313 11940 12317 11996
rect 12317 11940 12373 11996
rect 12373 11940 12377 11996
rect 12313 11936 12377 11940
rect 12393 11996 12457 12000
rect 12393 11940 12397 11996
rect 12397 11940 12453 11996
rect 12453 11940 12457 11996
rect 12393 11936 12457 11940
rect 12473 11996 12537 12000
rect 12473 11940 12477 11996
rect 12477 11940 12533 11996
rect 12533 11940 12537 11996
rect 12473 11936 12537 11940
rect 12553 11996 12617 12000
rect 12553 11940 12557 11996
rect 12557 11940 12613 11996
rect 12613 11940 12617 11996
rect 12553 11936 12617 11940
rect 17994 11996 18058 12000
rect 17994 11940 17998 11996
rect 17998 11940 18054 11996
rect 18054 11940 18058 11996
rect 17994 11936 18058 11940
rect 18074 11996 18138 12000
rect 18074 11940 18078 11996
rect 18078 11940 18134 11996
rect 18134 11940 18138 11996
rect 18074 11936 18138 11940
rect 18154 11996 18218 12000
rect 18154 11940 18158 11996
rect 18158 11940 18214 11996
rect 18214 11940 18218 11996
rect 18154 11936 18218 11940
rect 18234 11996 18298 12000
rect 18234 11940 18238 11996
rect 18238 11940 18294 11996
rect 18294 11940 18298 11996
rect 18234 11936 18298 11940
rect 23675 11996 23739 12000
rect 23675 11940 23679 11996
rect 23679 11940 23735 11996
rect 23735 11940 23739 11996
rect 23675 11936 23739 11940
rect 23755 11996 23819 12000
rect 23755 11940 23759 11996
rect 23759 11940 23815 11996
rect 23815 11940 23819 11996
rect 23755 11936 23819 11940
rect 23835 11996 23899 12000
rect 23835 11940 23839 11996
rect 23839 11940 23895 11996
rect 23895 11940 23899 11996
rect 23835 11936 23899 11940
rect 23915 11996 23979 12000
rect 23915 11940 23919 11996
rect 23919 11940 23975 11996
rect 23975 11940 23979 11996
rect 23915 11936 23979 11940
rect 3792 11452 3856 11456
rect 3792 11396 3796 11452
rect 3796 11396 3852 11452
rect 3852 11396 3856 11452
rect 3792 11392 3856 11396
rect 3872 11452 3936 11456
rect 3872 11396 3876 11452
rect 3876 11396 3932 11452
rect 3932 11396 3936 11452
rect 3872 11392 3936 11396
rect 3952 11452 4016 11456
rect 3952 11396 3956 11452
rect 3956 11396 4012 11452
rect 4012 11396 4016 11452
rect 3952 11392 4016 11396
rect 4032 11452 4096 11456
rect 4032 11396 4036 11452
rect 4036 11396 4092 11452
rect 4092 11396 4096 11452
rect 4032 11392 4096 11396
rect 9473 11452 9537 11456
rect 9473 11396 9477 11452
rect 9477 11396 9533 11452
rect 9533 11396 9537 11452
rect 9473 11392 9537 11396
rect 9553 11452 9617 11456
rect 9553 11396 9557 11452
rect 9557 11396 9613 11452
rect 9613 11396 9617 11452
rect 9553 11392 9617 11396
rect 9633 11452 9697 11456
rect 9633 11396 9637 11452
rect 9637 11396 9693 11452
rect 9693 11396 9697 11452
rect 9633 11392 9697 11396
rect 9713 11452 9777 11456
rect 9713 11396 9717 11452
rect 9717 11396 9773 11452
rect 9773 11396 9777 11452
rect 9713 11392 9777 11396
rect 15154 11452 15218 11456
rect 15154 11396 15158 11452
rect 15158 11396 15214 11452
rect 15214 11396 15218 11452
rect 15154 11392 15218 11396
rect 15234 11452 15298 11456
rect 15234 11396 15238 11452
rect 15238 11396 15294 11452
rect 15294 11396 15298 11452
rect 15234 11392 15298 11396
rect 15314 11452 15378 11456
rect 15314 11396 15318 11452
rect 15318 11396 15374 11452
rect 15374 11396 15378 11452
rect 15314 11392 15378 11396
rect 15394 11452 15458 11456
rect 15394 11396 15398 11452
rect 15398 11396 15454 11452
rect 15454 11396 15458 11452
rect 15394 11392 15458 11396
rect 20835 11452 20899 11456
rect 20835 11396 20839 11452
rect 20839 11396 20895 11452
rect 20895 11396 20899 11452
rect 20835 11392 20899 11396
rect 20915 11452 20979 11456
rect 20915 11396 20919 11452
rect 20919 11396 20975 11452
rect 20975 11396 20979 11452
rect 20915 11392 20979 11396
rect 20995 11452 21059 11456
rect 20995 11396 20999 11452
rect 20999 11396 21055 11452
rect 21055 11396 21059 11452
rect 20995 11392 21059 11396
rect 21075 11452 21139 11456
rect 21075 11396 21079 11452
rect 21079 11396 21135 11452
rect 21135 11396 21139 11452
rect 21075 11392 21139 11396
rect 17724 11052 17788 11116
rect 6632 10908 6696 10912
rect 6632 10852 6636 10908
rect 6636 10852 6692 10908
rect 6692 10852 6696 10908
rect 6632 10848 6696 10852
rect 6712 10908 6776 10912
rect 6712 10852 6716 10908
rect 6716 10852 6772 10908
rect 6772 10852 6776 10908
rect 6712 10848 6776 10852
rect 6792 10908 6856 10912
rect 6792 10852 6796 10908
rect 6796 10852 6852 10908
rect 6852 10852 6856 10908
rect 6792 10848 6856 10852
rect 6872 10908 6936 10912
rect 6872 10852 6876 10908
rect 6876 10852 6932 10908
rect 6932 10852 6936 10908
rect 6872 10848 6936 10852
rect 12313 10908 12377 10912
rect 12313 10852 12317 10908
rect 12317 10852 12373 10908
rect 12373 10852 12377 10908
rect 12313 10848 12377 10852
rect 12393 10908 12457 10912
rect 12393 10852 12397 10908
rect 12397 10852 12453 10908
rect 12453 10852 12457 10908
rect 12393 10848 12457 10852
rect 12473 10908 12537 10912
rect 12473 10852 12477 10908
rect 12477 10852 12533 10908
rect 12533 10852 12537 10908
rect 12473 10848 12537 10852
rect 12553 10908 12617 10912
rect 12553 10852 12557 10908
rect 12557 10852 12613 10908
rect 12613 10852 12617 10908
rect 12553 10848 12617 10852
rect 17994 10908 18058 10912
rect 17994 10852 17998 10908
rect 17998 10852 18054 10908
rect 18054 10852 18058 10908
rect 17994 10848 18058 10852
rect 18074 10908 18138 10912
rect 18074 10852 18078 10908
rect 18078 10852 18134 10908
rect 18134 10852 18138 10908
rect 18074 10848 18138 10852
rect 18154 10908 18218 10912
rect 18154 10852 18158 10908
rect 18158 10852 18214 10908
rect 18214 10852 18218 10908
rect 18154 10848 18218 10852
rect 18234 10908 18298 10912
rect 18234 10852 18238 10908
rect 18238 10852 18294 10908
rect 18294 10852 18298 10908
rect 18234 10848 18298 10852
rect 23675 10908 23739 10912
rect 23675 10852 23679 10908
rect 23679 10852 23735 10908
rect 23735 10852 23739 10908
rect 23675 10848 23739 10852
rect 23755 10908 23819 10912
rect 23755 10852 23759 10908
rect 23759 10852 23815 10908
rect 23815 10852 23819 10908
rect 23755 10848 23819 10852
rect 23835 10908 23899 10912
rect 23835 10852 23839 10908
rect 23839 10852 23895 10908
rect 23895 10852 23899 10908
rect 23835 10848 23899 10852
rect 23915 10908 23979 10912
rect 23915 10852 23919 10908
rect 23919 10852 23975 10908
rect 23975 10852 23979 10908
rect 23915 10848 23979 10852
rect 3792 10364 3856 10368
rect 3792 10308 3796 10364
rect 3796 10308 3852 10364
rect 3852 10308 3856 10364
rect 3792 10304 3856 10308
rect 3872 10364 3936 10368
rect 3872 10308 3876 10364
rect 3876 10308 3932 10364
rect 3932 10308 3936 10364
rect 3872 10304 3936 10308
rect 3952 10364 4016 10368
rect 3952 10308 3956 10364
rect 3956 10308 4012 10364
rect 4012 10308 4016 10364
rect 3952 10304 4016 10308
rect 4032 10364 4096 10368
rect 4032 10308 4036 10364
rect 4036 10308 4092 10364
rect 4092 10308 4096 10364
rect 4032 10304 4096 10308
rect 9473 10364 9537 10368
rect 9473 10308 9477 10364
rect 9477 10308 9533 10364
rect 9533 10308 9537 10364
rect 9473 10304 9537 10308
rect 9553 10364 9617 10368
rect 9553 10308 9557 10364
rect 9557 10308 9613 10364
rect 9613 10308 9617 10364
rect 9553 10304 9617 10308
rect 9633 10364 9697 10368
rect 9633 10308 9637 10364
rect 9637 10308 9693 10364
rect 9693 10308 9697 10364
rect 9633 10304 9697 10308
rect 9713 10364 9777 10368
rect 9713 10308 9717 10364
rect 9717 10308 9773 10364
rect 9773 10308 9777 10364
rect 9713 10304 9777 10308
rect 15154 10364 15218 10368
rect 15154 10308 15158 10364
rect 15158 10308 15214 10364
rect 15214 10308 15218 10364
rect 15154 10304 15218 10308
rect 15234 10364 15298 10368
rect 15234 10308 15238 10364
rect 15238 10308 15294 10364
rect 15294 10308 15298 10364
rect 15234 10304 15298 10308
rect 15314 10364 15378 10368
rect 15314 10308 15318 10364
rect 15318 10308 15374 10364
rect 15374 10308 15378 10364
rect 15314 10304 15378 10308
rect 15394 10364 15458 10368
rect 15394 10308 15398 10364
rect 15398 10308 15454 10364
rect 15454 10308 15458 10364
rect 15394 10304 15458 10308
rect 20835 10364 20899 10368
rect 20835 10308 20839 10364
rect 20839 10308 20895 10364
rect 20895 10308 20899 10364
rect 20835 10304 20899 10308
rect 20915 10364 20979 10368
rect 20915 10308 20919 10364
rect 20919 10308 20975 10364
rect 20975 10308 20979 10364
rect 20915 10304 20979 10308
rect 20995 10364 21059 10368
rect 20995 10308 20999 10364
rect 20999 10308 21055 10364
rect 21055 10308 21059 10364
rect 20995 10304 21059 10308
rect 21075 10364 21139 10368
rect 21075 10308 21079 10364
rect 21079 10308 21135 10364
rect 21135 10308 21139 10364
rect 21075 10304 21139 10308
rect 6632 9820 6696 9824
rect 6632 9764 6636 9820
rect 6636 9764 6692 9820
rect 6692 9764 6696 9820
rect 6632 9760 6696 9764
rect 6712 9820 6776 9824
rect 6712 9764 6716 9820
rect 6716 9764 6772 9820
rect 6772 9764 6776 9820
rect 6712 9760 6776 9764
rect 6792 9820 6856 9824
rect 6792 9764 6796 9820
rect 6796 9764 6852 9820
rect 6852 9764 6856 9820
rect 6792 9760 6856 9764
rect 6872 9820 6936 9824
rect 6872 9764 6876 9820
rect 6876 9764 6932 9820
rect 6932 9764 6936 9820
rect 6872 9760 6936 9764
rect 12313 9820 12377 9824
rect 12313 9764 12317 9820
rect 12317 9764 12373 9820
rect 12373 9764 12377 9820
rect 12313 9760 12377 9764
rect 12393 9820 12457 9824
rect 12393 9764 12397 9820
rect 12397 9764 12453 9820
rect 12453 9764 12457 9820
rect 12393 9760 12457 9764
rect 12473 9820 12537 9824
rect 12473 9764 12477 9820
rect 12477 9764 12533 9820
rect 12533 9764 12537 9820
rect 12473 9760 12537 9764
rect 12553 9820 12617 9824
rect 12553 9764 12557 9820
rect 12557 9764 12613 9820
rect 12613 9764 12617 9820
rect 12553 9760 12617 9764
rect 6316 9692 6380 9756
rect 4660 9556 4724 9620
rect 17994 9820 18058 9824
rect 17994 9764 17998 9820
rect 17998 9764 18054 9820
rect 18054 9764 18058 9820
rect 17994 9760 18058 9764
rect 18074 9820 18138 9824
rect 18074 9764 18078 9820
rect 18078 9764 18134 9820
rect 18134 9764 18138 9820
rect 18074 9760 18138 9764
rect 18154 9820 18218 9824
rect 18154 9764 18158 9820
rect 18158 9764 18214 9820
rect 18214 9764 18218 9820
rect 18154 9760 18218 9764
rect 18234 9820 18298 9824
rect 18234 9764 18238 9820
rect 18238 9764 18294 9820
rect 18294 9764 18298 9820
rect 18234 9760 18298 9764
rect 23675 9820 23739 9824
rect 23675 9764 23679 9820
rect 23679 9764 23735 9820
rect 23735 9764 23739 9820
rect 23675 9760 23739 9764
rect 23755 9820 23819 9824
rect 23755 9764 23759 9820
rect 23759 9764 23815 9820
rect 23815 9764 23819 9820
rect 23755 9760 23819 9764
rect 23835 9820 23899 9824
rect 23835 9764 23839 9820
rect 23839 9764 23895 9820
rect 23895 9764 23899 9820
rect 23835 9760 23899 9764
rect 23915 9820 23979 9824
rect 23915 9764 23919 9820
rect 23919 9764 23975 9820
rect 23975 9764 23979 9820
rect 23915 9760 23979 9764
rect 5764 9480 5828 9484
rect 5764 9424 5778 9480
rect 5778 9424 5828 9480
rect 5764 9420 5828 9424
rect 3792 9276 3856 9280
rect 3792 9220 3796 9276
rect 3796 9220 3852 9276
rect 3852 9220 3856 9276
rect 3792 9216 3856 9220
rect 3872 9276 3936 9280
rect 3872 9220 3876 9276
rect 3876 9220 3932 9276
rect 3932 9220 3936 9276
rect 3872 9216 3936 9220
rect 3952 9276 4016 9280
rect 3952 9220 3956 9276
rect 3956 9220 4012 9276
rect 4012 9220 4016 9276
rect 3952 9216 4016 9220
rect 4032 9276 4096 9280
rect 4032 9220 4036 9276
rect 4036 9220 4092 9276
rect 4092 9220 4096 9276
rect 4032 9216 4096 9220
rect 9473 9276 9537 9280
rect 9473 9220 9477 9276
rect 9477 9220 9533 9276
rect 9533 9220 9537 9276
rect 9473 9216 9537 9220
rect 9553 9276 9617 9280
rect 9553 9220 9557 9276
rect 9557 9220 9613 9276
rect 9613 9220 9617 9276
rect 9553 9216 9617 9220
rect 9633 9276 9697 9280
rect 9633 9220 9637 9276
rect 9637 9220 9693 9276
rect 9693 9220 9697 9276
rect 9633 9216 9697 9220
rect 9713 9276 9777 9280
rect 9713 9220 9717 9276
rect 9717 9220 9773 9276
rect 9773 9220 9777 9276
rect 9713 9216 9777 9220
rect 15154 9276 15218 9280
rect 15154 9220 15158 9276
rect 15158 9220 15214 9276
rect 15214 9220 15218 9276
rect 15154 9216 15218 9220
rect 15234 9276 15298 9280
rect 15234 9220 15238 9276
rect 15238 9220 15294 9276
rect 15294 9220 15298 9276
rect 15234 9216 15298 9220
rect 15314 9276 15378 9280
rect 15314 9220 15318 9276
rect 15318 9220 15374 9276
rect 15374 9220 15378 9276
rect 15314 9216 15378 9220
rect 15394 9276 15458 9280
rect 15394 9220 15398 9276
rect 15398 9220 15454 9276
rect 15454 9220 15458 9276
rect 15394 9216 15458 9220
rect 20835 9276 20899 9280
rect 20835 9220 20839 9276
rect 20839 9220 20895 9276
rect 20895 9220 20899 9276
rect 20835 9216 20899 9220
rect 20915 9276 20979 9280
rect 20915 9220 20919 9276
rect 20919 9220 20975 9276
rect 20975 9220 20979 9276
rect 20915 9216 20979 9220
rect 20995 9276 21059 9280
rect 20995 9220 20999 9276
rect 20999 9220 21055 9276
rect 21055 9220 21059 9276
rect 20995 9216 21059 9220
rect 21075 9276 21139 9280
rect 21075 9220 21079 9276
rect 21079 9220 21135 9276
rect 21135 9220 21139 9276
rect 21075 9216 21139 9220
rect 6632 8732 6696 8736
rect 6632 8676 6636 8732
rect 6636 8676 6692 8732
rect 6692 8676 6696 8732
rect 6632 8672 6696 8676
rect 6712 8732 6776 8736
rect 6712 8676 6716 8732
rect 6716 8676 6772 8732
rect 6772 8676 6776 8732
rect 6712 8672 6776 8676
rect 6792 8732 6856 8736
rect 6792 8676 6796 8732
rect 6796 8676 6852 8732
rect 6852 8676 6856 8732
rect 6792 8672 6856 8676
rect 6872 8732 6936 8736
rect 6872 8676 6876 8732
rect 6876 8676 6932 8732
rect 6932 8676 6936 8732
rect 6872 8672 6936 8676
rect 12313 8732 12377 8736
rect 12313 8676 12317 8732
rect 12317 8676 12373 8732
rect 12373 8676 12377 8732
rect 12313 8672 12377 8676
rect 12393 8732 12457 8736
rect 12393 8676 12397 8732
rect 12397 8676 12453 8732
rect 12453 8676 12457 8732
rect 12393 8672 12457 8676
rect 12473 8732 12537 8736
rect 12473 8676 12477 8732
rect 12477 8676 12533 8732
rect 12533 8676 12537 8732
rect 12473 8672 12537 8676
rect 12553 8732 12617 8736
rect 12553 8676 12557 8732
rect 12557 8676 12613 8732
rect 12613 8676 12617 8732
rect 12553 8672 12617 8676
rect 17994 8732 18058 8736
rect 17994 8676 17998 8732
rect 17998 8676 18054 8732
rect 18054 8676 18058 8732
rect 17994 8672 18058 8676
rect 18074 8732 18138 8736
rect 18074 8676 18078 8732
rect 18078 8676 18134 8732
rect 18134 8676 18138 8732
rect 18074 8672 18138 8676
rect 18154 8732 18218 8736
rect 18154 8676 18158 8732
rect 18158 8676 18214 8732
rect 18214 8676 18218 8732
rect 18154 8672 18218 8676
rect 18234 8732 18298 8736
rect 18234 8676 18238 8732
rect 18238 8676 18294 8732
rect 18294 8676 18298 8732
rect 18234 8672 18298 8676
rect 23675 8732 23739 8736
rect 23675 8676 23679 8732
rect 23679 8676 23735 8732
rect 23735 8676 23739 8732
rect 23675 8672 23739 8676
rect 23755 8732 23819 8736
rect 23755 8676 23759 8732
rect 23759 8676 23815 8732
rect 23815 8676 23819 8732
rect 23755 8672 23819 8676
rect 23835 8732 23899 8736
rect 23835 8676 23839 8732
rect 23839 8676 23895 8732
rect 23895 8676 23899 8732
rect 23835 8672 23899 8676
rect 23915 8732 23979 8736
rect 23915 8676 23919 8732
rect 23919 8676 23975 8732
rect 23975 8676 23979 8732
rect 23915 8672 23979 8676
rect 3792 8188 3856 8192
rect 3792 8132 3796 8188
rect 3796 8132 3852 8188
rect 3852 8132 3856 8188
rect 3792 8128 3856 8132
rect 3872 8188 3936 8192
rect 3872 8132 3876 8188
rect 3876 8132 3932 8188
rect 3932 8132 3936 8188
rect 3872 8128 3936 8132
rect 3952 8188 4016 8192
rect 3952 8132 3956 8188
rect 3956 8132 4012 8188
rect 4012 8132 4016 8188
rect 3952 8128 4016 8132
rect 4032 8188 4096 8192
rect 4032 8132 4036 8188
rect 4036 8132 4092 8188
rect 4092 8132 4096 8188
rect 4032 8128 4096 8132
rect 9473 8188 9537 8192
rect 9473 8132 9477 8188
rect 9477 8132 9533 8188
rect 9533 8132 9537 8188
rect 9473 8128 9537 8132
rect 9553 8188 9617 8192
rect 9553 8132 9557 8188
rect 9557 8132 9613 8188
rect 9613 8132 9617 8188
rect 9553 8128 9617 8132
rect 9633 8188 9697 8192
rect 9633 8132 9637 8188
rect 9637 8132 9693 8188
rect 9693 8132 9697 8188
rect 9633 8128 9697 8132
rect 9713 8188 9777 8192
rect 9713 8132 9717 8188
rect 9717 8132 9773 8188
rect 9773 8132 9777 8188
rect 9713 8128 9777 8132
rect 15154 8188 15218 8192
rect 15154 8132 15158 8188
rect 15158 8132 15214 8188
rect 15214 8132 15218 8188
rect 15154 8128 15218 8132
rect 15234 8188 15298 8192
rect 15234 8132 15238 8188
rect 15238 8132 15294 8188
rect 15294 8132 15298 8188
rect 15234 8128 15298 8132
rect 15314 8188 15378 8192
rect 15314 8132 15318 8188
rect 15318 8132 15374 8188
rect 15374 8132 15378 8188
rect 15314 8128 15378 8132
rect 15394 8188 15458 8192
rect 15394 8132 15398 8188
rect 15398 8132 15454 8188
rect 15454 8132 15458 8188
rect 15394 8128 15458 8132
rect 20835 8188 20899 8192
rect 20835 8132 20839 8188
rect 20839 8132 20895 8188
rect 20895 8132 20899 8188
rect 20835 8128 20899 8132
rect 20915 8188 20979 8192
rect 20915 8132 20919 8188
rect 20919 8132 20975 8188
rect 20975 8132 20979 8188
rect 20915 8128 20979 8132
rect 20995 8188 21059 8192
rect 20995 8132 20999 8188
rect 20999 8132 21055 8188
rect 21055 8132 21059 8188
rect 20995 8128 21059 8132
rect 21075 8188 21139 8192
rect 21075 8132 21079 8188
rect 21079 8132 21135 8188
rect 21135 8132 21139 8188
rect 21075 8128 21139 8132
rect 6632 7644 6696 7648
rect 6632 7588 6636 7644
rect 6636 7588 6692 7644
rect 6692 7588 6696 7644
rect 6632 7584 6696 7588
rect 6712 7644 6776 7648
rect 6712 7588 6716 7644
rect 6716 7588 6772 7644
rect 6772 7588 6776 7644
rect 6712 7584 6776 7588
rect 6792 7644 6856 7648
rect 6792 7588 6796 7644
rect 6796 7588 6852 7644
rect 6852 7588 6856 7644
rect 6792 7584 6856 7588
rect 6872 7644 6936 7648
rect 6872 7588 6876 7644
rect 6876 7588 6932 7644
rect 6932 7588 6936 7644
rect 6872 7584 6936 7588
rect 12313 7644 12377 7648
rect 12313 7588 12317 7644
rect 12317 7588 12373 7644
rect 12373 7588 12377 7644
rect 12313 7584 12377 7588
rect 12393 7644 12457 7648
rect 12393 7588 12397 7644
rect 12397 7588 12453 7644
rect 12453 7588 12457 7644
rect 12393 7584 12457 7588
rect 12473 7644 12537 7648
rect 12473 7588 12477 7644
rect 12477 7588 12533 7644
rect 12533 7588 12537 7644
rect 12473 7584 12537 7588
rect 12553 7644 12617 7648
rect 12553 7588 12557 7644
rect 12557 7588 12613 7644
rect 12613 7588 12617 7644
rect 12553 7584 12617 7588
rect 17994 7644 18058 7648
rect 17994 7588 17998 7644
rect 17998 7588 18054 7644
rect 18054 7588 18058 7644
rect 17994 7584 18058 7588
rect 18074 7644 18138 7648
rect 18074 7588 18078 7644
rect 18078 7588 18134 7644
rect 18134 7588 18138 7644
rect 18074 7584 18138 7588
rect 18154 7644 18218 7648
rect 18154 7588 18158 7644
rect 18158 7588 18214 7644
rect 18214 7588 18218 7644
rect 18154 7584 18218 7588
rect 18234 7644 18298 7648
rect 18234 7588 18238 7644
rect 18238 7588 18294 7644
rect 18294 7588 18298 7644
rect 18234 7584 18298 7588
rect 23675 7644 23739 7648
rect 23675 7588 23679 7644
rect 23679 7588 23735 7644
rect 23735 7588 23739 7644
rect 23675 7584 23739 7588
rect 23755 7644 23819 7648
rect 23755 7588 23759 7644
rect 23759 7588 23815 7644
rect 23815 7588 23819 7644
rect 23755 7584 23819 7588
rect 23835 7644 23899 7648
rect 23835 7588 23839 7644
rect 23839 7588 23895 7644
rect 23895 7588 23899 7644
rect 23835 7584 23899 7588
rect 23915 7644 23979 7648
rect 23915 7588 23919 7644
rect 23919 7588 23975 7644
rect 23975 7588 23979 7644
rect 23915 7584 23979 7588
rect 3792 7100 3856 7104
rect 3792 7044 3796 7100
rect 3796 7044 3852 7100
rect 3852 7044 3856 7100
rect 3792 7040 3856 7044
rect 3872 7100 3936 7104
rect 3872 7044 3876 7100
rect 3876 7044 3932 7100
rect 3932 7044 3936 7100
rect 3872 7040 3936 7044
rect 3952 7100 4016 7104
rect 3952 7044 3956 7100
rect 3956 7044 4012 7100
rect 4012 7044 4016 7100
rect 3952 7040 4016 7044
rect 4032 7100 4096 7104
rect 4032 7044 4036 7100
rect 4036 7044 4092 7100
rect 4092 7044 4096 7100
rect 4032 7040 4096 7044
rect 9473 7100 9537 7104
rect 9473 7044 9477 7100
rect 9477 7044 9533 7100
rect 9533 7044 9537 7100
rect 9473 7040 9537 7044
rect 9553 7100 9617 7104
rect 9553 7044 9557 7100
rect 9557 7044 9613 7100
rect 9613 7044 9617 7100
rect 9553 7040 9617 7044
rect 9633 7100 9697 7104
rect 9633 7044 9637 7100
rect 9637 7044 9693 7100
rect 9693 7044 9697 7100
rect 9633 7040 9697 7044
rect 9713 7100 9777 7104
rect 9713 7044 9717 7100
rect 9717 7044 9773 7100
rect 9773 7044 9777 7100
rect 9713 7040 9777 7044
rect 15154 7100 15218 7104
rect 15154 7044 15158 7100
rect 15158 7044 15214 7100
rect 15214 7044 15218 7100
rect 15154 7040 15218 7044
rect 15234 7100 15298 7104
rect 15234 7044 15238 7100
rect 15238 7044 15294 7100
rect 15294 7044 15298 7100
rect 15234 7040 15298 7044
rect 15314 7100 15378 7104
rect 15314 7044 15318 7100
rect 15318 7044 15374 7100
rect 15374 7044 15378 7100
rect 15314 7040 15378 7044
rect 15394 7100 15458 7104
rect 15394 7044 15398 7100
rect 15398 7044 15454 7100
rect 15454 7044 15458 7100
rect 15394 7040 15458 7044
rect 20835 7100 20899 7104
rect 20835 7044 20839 7100
rect 20839 7044 20895 7100
rect 20895 7044 20899 7100
rect 20835 7040 20899 7044
rect 20915 7100 20979 7104
rect 20915 7044 20919 7100
rect 20919 7044 20975 7100
rect 20975 7044 20979 7100
rect 20915 7040 20979 7044
rect 20995 7100 21059 7104
rect 20995 7044 20999 7100
rect 20999 7044 21055 7100
rect 21055 7044 21059 7100
rect 20995 7040 21059 7044
rect 21075 7100 21139 7104
rect 21075 7044 21079 7100
rect 21079 7044 21135 7100
rect 21135 7044 21139 7100
rect 21075 7040 21139 7044
rect 14596 6836 14660 6900
rect 6632 6556 6696 6560
rect 6632 6500 6636 6556
rect 6636 6500 6692 6556
rect 6692 6500 6696 6556
rect 6632 6496 6696 6500
rect 6712 6556 6776 6560
rect 6712 6500 6716 6556
rect 6716 6500 6772 6556
rect 6772 6500 6776 6556
rect 6712 6496 6776 6500
rect 6792 6556 6856 6560
rect 6792 6500 6796 6556
rect 6796 6500 6852 6556
rect 6852 6500 6856 6556
rect 6792 6496 6856 6500
rect 6872 6556 6936 6560
rect 6872 6500 6876 6556
rect 6876 6500 6932 6556
rect 6932 6500 6936 6556
rect 6872 6496 6936 6500
rect 12313 6556 12377 6560
rect 12313 6500 12317 6556
rect 12317 6500 12373 6556
rect 12373 6500 12377 6556
rect 12313 6496 12377 6500
rect 12393 6556 12457 6560
rect 12393 6500 12397 6556
rect 12397 6500 12453 6556
rect 12453 6500 12457 6556
rect 12393 6496 12457 6500
rect 12473 6556 12537 6560
rect 12473 6500 12477 6556
rect 12477 6500 12533 6556
rect 12533 6500 12537 6556
rect 12473 6496 12537 6500
rect 12553 6556 12617 6560
rect 12553 6500 12557 6556
rect 12557 6500 12613 6556
rect 12613 6500 12617 6556
rect 12553 6496 12617 6500
rect 17994 6556 18058 6560
rect 17994 6500 17998 6556
rect 17998 6500 18054 6556
rect 18054 6500 18058 6556
rect 17994 6496 18058 6500
rect 18074 6556 18138 6560
rect 18074 6500 18078 6556
rect 18078 6500 18134 6556
rect 18134 6500 18138 6556
rect 18074 6496 18138 6500
rect 18154 6556 18218 6560
rect 18154 6500 18158 6556
rect 18158 6500 18214 6556
rect 18214 6500 18218 6556
rect 18154 6496 18218 6500
rect 18234 6556 18298 6560
rect 18234 6500 18238 6556
rect 18238 6500 18294 6556
rect 18294 6500 18298 6556
rect 18234 6496 18298 6500
rect 23675 6556 23739 6560
rect 23675 6500 23679 6556
rect 23679 6500 23735 6556
rect 23735 6500 23739 6556
rect 23675 6496 23739 6500
rect 23755 6556 23819 6560
rect 23755 6500 23759 6556
rect 23759 6500 23815 6556
rect 23815 6500 23819 6556
rect 23755 6496 23819 6500
rect 23835 6556 23899 6560
rect 23835 6500 23839 6556
rect 23839 6500 23895 6556
rect 23895 6500 23899 6556
rect 23835 6496 23899 6500
rect 23915 6556 23979 6560
rect 23915 6500 23919 6556
rect 23919 6500 23975 6556
rect 23975 6500 23979 6556
rect 23915 6496 23979 6500
rect 3792 6012 3856 6016
rect 3792 5956 3796 6012
rect 3796 5956 3852 6012
rect 3852 5956 3856 6012
rect 3792 5952 3856 5956
rect 3872 6012 3936 6016
rect 3872 5956 3876 6012
rect 3876 5956 3932 6012
rect 3932 5956 3936 6012
rect 3872 5952 3936 5956
rect 3952 6012 4016 6016
rect 3952 5956 3956 6012
rect 3956 5956 4012 6012
rect 4012 5956 4016 6012
rect 3952 5952 4016 5956
rect 4032 6012 4096 6016
rect 4032 5956 4036 6012
rect 4036 5956 4092 6012
rect 4092 5956 4096 6012
rect 4032 5952 4096 5956
rect 9473 6012 9537 6016
rect 9473 5956 9477 6012
rect 9477 5956 9533 6012
rect 9533 5956 9537 6012
rect 9473 5952 9537 5956
rect 9553 6012 9617 6016
rect 9553 5956 9557 6012
rect 9557 5956 9613 6012
rect 9613 5956 9617 6012
rect 9553 5952 9617 5956
rect 9633 6012 9697 6016
rect 9633 5956 9637 6012
rect 9637 5956 9693 6012
rect 9693 5956 9697 6012
rect 9633 5952 9697 5956
rect 9713 6012 9777 6016
rect 9713 5956 9717 6012
rect 9717 5956 9773 6012
rect 9773 5956 9777 6012
rect 9713 5952 9777 5956
rect 15154 6012 15218 6016
rect 15154 5956 15158 6012
rect 15158 5956 15214 6012
rect 15214 5956 15218 6012
rect 15154 5952 15218 5956
rect 15234 6012 15298 6016
rect 15234 5956 15238 6012
rect 15238 5956 15294 6012
rect 15294 5956 15298 6012
rect 15234 5952 15298 5956
rect 15314 6012 15378 6016
rect 15314 5956 15318 6012
rect 15318 5956 15374 6012
rect 15374 5956 15378 6012
rect 15314 5952 15378 5956
rect 15394 6012 15458 6016
rect 15394 5956 15398 6012
rect 15398 5956 15454 6012
rect 15454 5956 15458 6012
rect 15394 5952 15458 5956
rect 20835 6012 20899 6016
rect 20835 5956 20839 6012
rect 20839 5956 20895 6012
rect 20895 5956 20899 6012
rect 20835 5952 20899 5956
rect 20915 6012 20979 6016
rect 20915 5956 20919 6012
rect 20919 5956 20975 6012
rect 20975 5956 20979 6012
rect 20915 5952 20979 5956
rect 20995 6012 21059 6016
rect 20995 5956 20999 6012
rect 20999 5956 21055 6012
rect 21055 5956 21059 6012
rect 20995 5952 21059 5956
rect 21075 6012 21139 6016
rect 21075 5956 21079 6012
rect 21079 5956 21135 6012
rect 21135 5956 21139 6012
rect 21075 5952 21139 5956
rect 19932 5612 19996 5676
rect 6632 5468 6696 5472
rect 6632 5412 6636 5468
rect 6636 5412 6692 5468
rect 6692 5412 6696 5468
rect 6632 5408 6696 5412
rect 6712 5468 6776 5472
rect 6712 5412 6716 5468
rect 6716 5412 6772 5468
rect 6772 5412 6776 5468
rect 6712 5408 6776 5412
rect 6792 5468 6856 5472
rect 6792 5412 6796 5468
rect 6796 5412 6852 5468
rect 6852 5412 6856 5468
rect 6792 5408 6856 5412
rect 6872 5468 6936 5472
rect 6872 5412 6876 5468
rect 6876 5412 6932 5468
rect 6932 5412 6936 5468
rect 6872 5408 6936 5412
rect 12313 5468 12377 5472
rect 12313 5412 12317 5468
rect 12317 5412 12373 5468
rect 12373 5412 12377 5468
rect 12313 5408 12377 5412
rect 12393 5468 12457 5472
rect 12393 5412 12397 5468
rect 12397 5412 12453 5468
rect 12453 5412 12457 5468
rect 12393 5408 12457 5412
rect 12473 5468 12537 5472
rect 12473 5412 12477 5468
rect 12477 5412 12533 5468
rect 12533 5412 12537 5468
rect 12473 5408 12537 5412
rect 12553 5468 12617 5472
rect 12553 5412 12557 5468
rect 12557 5412 12613 5468
rect 12613 5412 12617 5468
rect 12553 5408 12617 5412
rect 17994 5468 18058 5472
rect 17994 5412 17998 5468
rect 17998 5412 18054 5468
rect 18054 5412 18058 5468
rect 17994 5408 18058 5412
rect 18074 5468 18138 5472
rect 18074 5412 18078 5468
rect 18078 5412 18134 5468
rect 18134 5412 18138 5468
rect 18074 5408 18138 5412
rect 18154 5468 18218 5472
rect 18154 5412 18158 5468
rect 18158 5412 18214 5468
rect 18214 5412 18218 5468
rect 18154 5408 18218 5412
rect 18234 5468 18298 5472
rect 18234 5412 18238 5468
rect 18238 5412 18294 5468
rect 18294 5412 18298 5468
rect 18234 5408 18298 5412
rect 23675 5468 23739 5472
rect 23675 5412 23679 5468
rect 23679 5412 23735 5468
rect 23735 5412 23739 5468
rect 23675 5408 23739 5412
rect 23755 5468 23819 5472
rect 23755 5412 23759 5468
rect 23759 5412 23815 5468
rect 23815 5412 23819 5468
rect 23755 5408 23819 5412
rect 23835 5468 23899 5472
rect 23835 5412 23839 5468
rect 23839 5412 23895 5468
rect 23895 5412 23899 5468
rect 23835 5408 23899 5412
rect 23915 5468 23979 5472
rect 23915 5412 23919 5468
rect 23919 5412 23975 5468
rect 23975 5412 23979 5468
rect 23915 5408 23979 5412
rect 17724 5204 17788 5268
rect 3792 4924 3856 4928
rect 3792 4868 3796 4924
rect 3796 4868 3852 4924
rect 3852 4868 3856 4924
rect 3792 4864 3856 4868
rect 3872 4924 3936 4928
rect 3872 4868 3876 4924
rect 3876 4868 3932 4924
rect 3932 4868 3936 4924
rect 3872 4864 3936 4868
rect 3952 4924 4016 4928
rect 3952 4868 3956 4924
rect 3956 4868 4012 4924
rect 4012 4868 4016 4924
rect 3952 4864 4016 4868
rect 4032 4924 4096 4928
rect 4032 4868 4036 4924
rect 4036 4868 4092 4924
rect 4092 4868 4096 4924
rect 4032 4864 4096 4868
rect 9473 4924 9537 4928
rect 9473 4868 9477 4924
rect 9477 4868 9533 4924
rect 9533 4868 9537 4924
rect 9473 4864 9537 4868
rect 9553 4924 9617 4928
rect 9553 4868 9557 4924
rect 9557 4868 9613 4924
rect 9613 4868 9617 4924
rect 9553 4864 9617 4868
rect 9633 4924 9697 4928
rect 9633 4868 9637 4924
rect 9637 4868 9693 4924
rect 9693 4868 9697 4924
rect 9633 4864 9697 4868
rect 9713 4924 9777 4928
rect 9713 4868 9717 4924
rect 9717 4868 9773 4924
rect 9773 4868 9777 4924
rect 9713 4864 9777 4868
rect 15154 4924 15218 4928
rect 15154 4868 15158 4924
rect 15158 4868 15214 4924
rect 15214 4868 15218 4924
rect 15154 4864 15218 4868
rect 15234 4924 15298 4928
rect 15234 4868 15238 4924
rect 15238 4868 15294 4924
rect 15294 4868 15298 4924
rect 15234 4864 15298 4868
rect 15314 4924 15378 4928
rect 15314 4868 15318 4924
rect 15318 4868 15374 4924
rect 15374 4868 15378 4924
rect 15314 4864 15378 4868
rect 15394 4924 15458 4928
rect 15394 4868 15398 4924
rect 15398 4868 15454 4924
rect 15454 4868 15458 4924
rect 15394 4864 15458 4868
rect 20835 4924 20899 4928
rect 20835 4868 20839 4924
rect 20839 4868 20895 4924
rect 20895 4868 20899 4924
rect 20835 4864 20899 4868
rect 20915 4924 20979 4928
rect 20915 4868 20919 4924
rect 20919 4868 20975 4924
rect 20975 4868 20979 4924
rect 20915 4864 20979 4868
rect 20995 4924 21059 4928
rect 20995 4868 20999 4924
rect 20999 4868 21055 4924
rect 21055 4868 21059 4924
rect 20995 4864 21059 4868
rect 21075 4924 21139 4928
rect 21075 4868 21079 4924
rect 21079 4868 21135 4924
rect 21135 4868 21139 4924
rect 21075 4864 21139 4868
rect 6632 4380 6696 4384
rect 6632 4324 6636 4380
rect 6636 4324 6692 4380
rect 6692 4324 6696 4380
rect 6632 4320 6696 4324
rect 6712 4380 6776 4384
rect 6712 4324 6716 4380
rect 6716 4324 6772 4380
rect 6772 4324 6776 4380
rect 6712 4320 6776 4324
rect 6792 4380 6856 4384
rect 6792 4324 6796 4380
rect 6796 4324 6852 4380
rect 6852 4324 6856 4380
rect 6792 4320 6856 4324
rect 6872 4380 6936 4384
rect 6872 4324 6876 4380
rect 6876 4324 6932 4380
rect 6932 4324 6936 4380
rect 6872 4320 6936 4324
rect 12313 4380 12377 4384
rect 12313 4324 12317 4380
rect 12317 4324 12373 4380
rect 12373 4324 12377 4380
rect 12313 4320 12377 4324
rect 12393 4380 12457 4384
rect 12393 4324 12397 4380
rect 12397 4324 12453 4380
rect 12453 4324 12457 4380
rect 12393 4320 12457 4324
rect 12473 4380 12537 4384
rect 12473 4324 12477 4380
rect 12477 4324 12533 4380
rect 12533 4324 12537 4380
rect 12473 4320 12537 4324
rect 12553 4380 12617 4384
rect 12553 4324 12557 4380
rect 12557 4324 12613 4380
rect 12613 4324 12617 4380
rect 12553 4320 12617 4324
rect 17994 4380 18058 4384
rect 17994 4324 17998 4380
rect 17998 4324 18054 4380
rect 18054 4324 18058 4380
rect 17994 4320 18058 4324
rect 18074 4380 18138 4384
rect 18074 4324 18078 4380
rect 18078 4324 18134 4380
rect 18134 4324 18138 4380
rect 18074 4320 18138 4324
rect 18154 4380 18218 4384
rect 18154 4324 18158 4380
rect 18158 4324 18214 4380
rect 18214 4324 18218 4380
rect 18154 4320 18218 4324
rect 18234 4380 18298 4384
rect 18234 4324 18238 4380
rect 18238 4324 18294 4380
rect 18294 4324 18298 4380
rect 18234 4320 18298 4324
rect 23675 4380 23739 4384
rect 23675 4324 23679 4380
rect 23679 4324 23735 4380
rect 23735 4324 23739 4380
rect 23675 4320 23739 4324
rect 23755 4380 23819 4384
rect 23755 4324 23759 4380
rect 23759 4324 23815 4380
rect 23815 4324 23819 4380
rect 23755 4320 23819 4324
rect 23835 4380 23899 4384
rect 23835 4324 23839 4380
rect 23839 4324 23895 4380
rect 23895 4324 23899 4380
rect 23835 4320 23899 4324
rect 23915 4380 23979 4384
rect 23915 4324 23919 4380
rect 23919 4324 23975 4380
rect 23975 4324 23979 4380
rect 23915 4320 23979 4324
rect 5764 3980 5828 4044
rect 3792 3836 3856 3840
rect 3792 3780 3796 3836
rect 3796 3780 3852 3836
rect 3852 3780 3856 3836
rect 3792 3776 3856 3780
rect 3872 3836 3936 3840
rect 3872 3780 3876 3836
rect 3876 3780 3932 3836
rect 3932 3780 3936 3836
rect 3872 3776 3936 3780
rect 3952 3836 4016 3840
rect 3952 3780 3956 3836
rect 3956 3780 4012 3836
rect 4012 3780 4016 3836
rect 3952 3776 4016 3780
rect 4032 3836 4096 3840
rect 4032 3780 4036 3836
rect 4036 3780 4092 3836
rect 4092 3780 4096 3836
rect 4032 3776 4096 3780
rect 9473 3836 9537 3840
rect 9473 3780 9477 3836
rect 9477 3780 9533 3836
rect 9533 3780 9537 3836
rect 9473 3776 9537 3780
rect 9553 3836 9617 3840
rect 9553 3780 9557 3836
rect 9557 3780 9613 3836
rect 9613 3780 9617 3836
rect 9553 3776 9617 3780
rect 9633 3836 9697 3840
rect 9633 3780 9637 3836
rect 9637 3780 9693 3836
rect 9693 3780 9697 3836
rect 9633 3776 9697 3780
rect 9713 3836 9777 3840
rect 9713 3780 9717 3836
rect 9717 3780 9773 3836
rect 9773 3780 9777 3836
rect 9713 3776 9777 3780
rect 15154 3836 15218 3840
rect 15154 3780 15158 3836
rect 15158 3780 15214 3836
rect 15214 3780 15218 3836
rect 15154 3776 15218 3780
rect 15234 3836 15298 3840
rect 15234 3780 15238 3836
rect 15238 3780 15294 3836
rect 15294 3780 15298 3836
rect 15234 3776 15298 3780
rect 15314 3836 15378 3840
rect 15314 3780 15318 3836
rect 15318 3780 15374 3836
rect 15374 3780 15378 3836
rect 15314 3776 15378 3780
rect 15394 3836 15458 3840
rect 15394 3780 15398 3836
rect 15398 3780 15454 3836
rect 15454 3780 15458 3836
rect 15394 3776 15458 3780
rect 20835 3836 20899 3840
rect 20835 3780 20839 3836
rect 20839 3780 20895 3836
rect 20895 3780 20899 3836
rect 20835 3776 20899 3780
rect 20915 3836 20979 3840
rect 20915 3780 20919 3836
rect 20919 3780 20975 3836
rect 20975 3780 20979 3836
rect 20915 3776 20979 3780
rect 20995 3836 21059 3840
rect 20995 3780 20999 3836
rect 20999 3780 21055 3836
rect 21055 3780 21059 3836
rect 20995 3776 21059 3780
rect 21075 3836 21139 3840
rect 21075 3780 21079 3836
rect 21079 3780 21135 3836
rect 21135 3780 21139 3836
rect 21075 3776 21139 3780
rect 6632 3292 6696 3296
rect 6632 3236 6636 3292
rect 6636 3236 6692 3292
rect 6692 3236 6696 3292
rect 6632 3232 6696 3236
rect 6712 3292 6776 3296
rect 6712 3236 6716 3292
rect 6716 3236 6772 3292
rect 6772 3236 6776 3292
rect 6712 3232 6776 3236
rect 6792 3292 6856 3296
rect 6792 3236 6796 3292
rect 6796 3236 6852 3292
rect 6852 3236 6856 3292
rect 6792 3232 6856 3236
rect 6872 3292 6936 3296
rect 6872 3236 6876 3292
rect 6876 3236 6932 3292
rect 6932 3236 6936 3292
rect 6872 3232 6936 3236
rect 12313 3292 12377 3296
rect 12313 3236 12317 3292
rect 12317 3236 12373 3292
rect 12373 3236 12377 3292
rect 12313 3232 12377 3236
rect 12393 3292 12457 3296
rect 12393 3236 12397 3292
rect 12397 3236 12453 3292
rect 12453 3236 12457 3292
rect 12393 3232 12457 3236
rect 12473 3292 12537 3296
rect 12473 3236 12477 3292
rect 12477 3236 12533 3292
rect 12533 3236 12537 3292
rect 12473 3232 12537 3236
rect 12553 3292 12617 3296
rect 12553 3236 12557 3292
rect 12557 3236 12613 3292
rect 12613 3236 12617 3292
rect 12553 3232 12617 3236
rect 17994 3292 18058 3296
rect 17994 3236 17998 3292
rect 17998 3236 18054 3292
rect 18054 3236 18058 3292
rect 17994 3232 18058 3236
rect 18074 3292 18138 3296
rect 18074 3236 18078 3292
rect 18078 3236 18134 3292
rect 18134 3236 18138 3292
rect 18074 3232 18138 3236
rect 18154 3292 18218 3296
rect 18154 3236 18158 3292
rect 18158 3236 18214 3292
rect 18214 3236 18218 3292
rect 18154 3232 18218 3236
rect 18234 3292 18298 3296
rect 18234 3236 18238 3292
rect 18238 3236 18294 3292
rect 18294 3236 18298 3292
rect 18234 3232 18298 3236
rect 23675 3292 23739 3296
rect 23675 3236 23679 3292
rect 23679 3236 23735 3292
rect 23735 3236 23739 3292
rect 23675 3232 23739 3236
rect 23755 3292 23819 3296
rect 23755 3236 23759 3292
rect 23759 3236 23815 3292
rect 23815 3236 23819 3292
rect 23755 3232 23819 3236
rect 23835 3292 23899 3296
rect 23835 3236 23839 3292
rect 23839 3236 23895 3292
rect 23895 3236 23899 3292
rect 23835 3232 23899 3236
rect 23915 3292 23979 3296
rect 23915 3236 23919 3292
rect 23919 3236 23975 3292
rect 23975 3236 23979 3292
rect 23915 3232 23979 3236
rect 4292 3028 4356 3092
rect 5396 3028 5460 3092
rect 3792 2748 3856 2752
rect 3792 2692 3796 2748
rect 3796 2692 3852 2748
rect 3852 2692 3856 2748
rect 3792 2688 3856 2692
rect 3872 2748 3936 2752
rect 3872 2692 3876 2748
rect 3876 2692 3932 2748
rect 3932 2692 3936 2748
rect 3872 2688 3936 2692
rect 3952 2748 4016 2752
rect 3952 2692 3956 2748
rect 3956 2692 4012 2748
rect 4012 2692 4016 2748
rect 3952 2688 4016 2692
rect 4032 2748 4096 2752
rect 4032 2692 4036 2748
rect 4036 2692 4092 2748
rect 4092 2692 4096 2748
rect 4032 2688 4096 2692
rect 9473 2748 9537 2752
rect 9473 2692 9477 2748
rect 9477 2692 9533 2748
rect 9533 2692 9537 2748
rect 9473 2688 9537 2692
rect 9553 2748 9617 2752
rect 9553 2692 9557 2748
rect 9557 2692 9613 2748
rect 9613 2692 9617 2748
rect 9553 2688 9617 2692
rect 9633 2748 9697 2752
rect 9633 2692 9637 2748
rect 9637 2692 9693 2748
rect 9693 2692 9697 2748
rect 9633 2688 9697 2692
rect 9713 2748 9777 2752
rect 9713 2692 9717 2748
rect 9717 2692 9773 2748
rect 9773 2692 9777 2748
rect 9713 2688 9777 2692
rect 15154 2748 15218 2752
rect 15154 2692 15158 2748
rect 15158 2692 15214 2748
rect 15214 2692 15218 2748
rect 15154 2688 15218 2692
rect 15234 2748 15298 2752
rect 15234 2692 15238 2748
rect 15238 2692 15294 2748
rect 15294 2692 15298 2748
rect 15234 2688 15298 2692
rect 15314 2748 15378 2752
rect 15314 2692 15318 2748
rect 15318 2692 15374 2748
rect 15374 2692 15378 2748
rect 15314 2688 15378 2692
rect 15394 2748 15458 2752
rect 15394 2692 15398 2748
rect 15398 2692 15454 2748
rect 15454 2692 15458 2748
rect 15394 2688 15458 2692
rect 20835 2748 20899 2752
rect 20835 2692 20839 2748
rect 20839 2692 20895 2748
rect 20895 2692 20899 2748
rect 20835 2688 20899 2692
rect 20915 2748 20979 2752
rect 20915 2692 20919 2748
rect 20919 2692 20975 2748
rect 20975 2692 20979 2748
rect 20915 2688 20979 2692
rect 20995 2748 21059 2752
rect 20995 2692 20999 2748
rect 20999 2692 21055 2748
rect 21055 2692 21059 2748
rect 20995 2688 21059 2692
rect 21075 2748 21139 2752
rect 21075 2692 21079 2748
rect 21079 2692 21135 2748
rect 21135 2692 21139 2748
rect 21075 2688 21139 2692
rect 4292 2484 4356 2548
rect 6632 2204 6696 2208
rect 6632 2148 6636 2204
rect 6636 2148 6692 2204
rect 6692 2148 6696 2204
rect 6632 2144 6696 2148
rect 6712 2204 6776 2208
rect 6712 2148 6716 2204
rect 6716 2148 6772 2204
rect 6772 2148 6776 2204
rect 6712 2144 6776 2148
rect 6792 2204 6856 2208
rect 6792 2148 6796 2204
rect 6796 2148 6852 2204
rect 6852 2148 6856 2204
rect 6792 2144 6856 2148
rect 6872 2204 6936 2208
rect 6872 2148 6876 2204
rect 6876 2148 6932 2204
rect 6932 2148 6936 2204
rect 6872 2144 6936 2148
rect 12313 2204 12377 2208
rect 12313 2148 12317 2204
rect 12317 2148 12373 2204
rect 12373 2148 12377 2204
rect 12313 2144 12377 2148
rect 12393 2204 12457 2208
rect 12393 2148 12397 2204
rect 12397 2148 12453 2204
rect 12453 2148 12457 2204
rect 12393 2144 12457 2148
rect 12473 2204 12537 2208
rect 12473 2148 12477 2204
rect 12477 2148 12533 2204
rect 12533 2148 12537 2204
rect 12473 2144 12537 2148
rect 12553 2204 12617 2208
rect 12553 2148 12557 2204
rect 12557 2148 12613 2204
rect 12613 2148 12617 2204
rect 12553 2144 12617 2148
rect 17994 2204 18058 2208
rect 17994 2148 17998 2204
rect 17998 2148 18054 2204
rect 18054 2148 18058 2204
rect 17994 2144 18058 2148
rect 18074 2204 18138 2208
rect 18074 2148 18078 2204
rect 18078 2148 18134 2204
rect 18134 2148 18138 2204
rect 18074 2144 18138 2148
rect 18154 2204 18218 2208
rect 18154 2148 18158 2204
rect 18158 2148 18214 2204
rect 18214 2148 18218 2204
rect 18154 2144 18218 2148
rect 18234 2204 18298 2208
rect 18234 2148 18238 2204
rect 18238 2148 18294 2204
rect 18294 2148 18298 2204
rect 18234 2144 18298 2148
rect 23675 2204 23739 2208
rect 23675 2148 23679 2204
rect 23679 2148 23735 2204
rect 23735 2148 23739 2204
rect 23675 2144 23739 2148
rect 23755 2204 23819 2208
rect 23755 2148 23759 2204
rect 23759 2148 23815 2204
rect 23815 2148 23819 2204
rect 23755 2144 23819 2148
rect 23835 2204 23899 2208
rect 23835 2148 23839 2204
rect 23839 2148 23895 2204
rect 23895 2148 23899 2204
rect 23835 2144 23899 2148
rect 23915 2204 23979 2208
rect 23915 2148 23919 2204
rect 23919 2148 23975 2204
rect 23975 2148 23979 2204
rect 23915 2144 23979 2148
<< metal4 >>
rect 3784 22336 4104 22352
rect 3784 22272 3792 22336
rect 3856 22272 3872 22336
rect 3936 22272 3952 22336
rect 4016 22272 4032 22336
rect 4096 22272 4104 22336
rect 3784 21248 4104 22272
rect 3784 21184 3792 21248
rect 3856 21184 3872 21248
rect 3936 21184 3952 21248
rect 4016 21184 4032 21248
rect 4096 21184 4104 21248
rect 3784 20160 4104 21184
rect 6624 21792 6944 22352
rect 6624 21728 6632 21792
rect 6696 21728 6712 21792
rect 6776 21728 6792 21792
rect 6856 21728 6872 21792
rect 6936 21728 6944 21792
rect 4659 20772 4725 20773
rect 4659 20708 4660 20772
rect 4724 20708 4725 20772
rect 4659 20707 4725 20708
rect 3784 20096 3792 20160
rect 3856 20096 3872 20160
rect 3936 20096 3952 20160
rect 4016 20096 4032 20160
rect 4096 20096 4104 20160
rect 3784 19072 4104 20096
rect 3784 19008 3792 19072
rect 3856 19008 3872 19072
rect 3936 19008 3952 19072
rect 4016 19008 4032 19072
rect 4096 19008 4104 19072
rect 3784 17984 4104 19008
rect 3784 17920 3792 17984
rect 3856 17920 3872 17984
rect 3936 17920 3952 17984
rect 4016 17920 4032 17984
rect 4096 17920 4104 17984
rect 3784 16896 4104 17920
rect 3784 16832 3792 16896
rect 3856 16832 3872 16896
rect 3936 16832 3952 16896
rect 4016 16832 4032 16896
rect 4096 16832 4104 16896
rect 3784 15808 4104 16832
rect 3784 15744 3792 15808
rect 3856 15744 3872 15808
rect 3936 15744 3952 15808
rect 4016 15744 4032 15808
rect 4096 15744 4104 15808
rect 3784 14720 4104 15744
rect 3784 14656 3792 14720
rect 3856 14656 3872 14720
rect 3936 14656 3952 14720
rect 4016 14656 4032 14720
rect 4096 14656 4104 14720
rect 3784 13632 4104 14656
rect 3784 13568 3792 13632
rect 3856 13568 3872 13632
rect 3936 13568 3952 13632
rect 4016 13568 4032 13632
rect 4096 13568 4104 13632
rect 3784 12544 4104 13568
rect 3784 12480 3792 12544
rect 3856 12480 3872 12544
rect 3936 12480 3952 12544
rect 4016 12480 4032 12544
rect 4096 12480 4104 12544
rect 3784 11456 4104 12480
rect 3784 11392 3792 11456
rect 3856 11392 3872 11456
rect 3936 11392 3952 11456
rect 4016 11392 4032 11456
rect 4096 11392 4104 11456
rect 3784 10368 4104 11392
rect 3784 10304 3792 10368
rect 3856 10304 3872 10368
rect 3936 10304 3952 10368
rect 4016 10304 4032 10368
rect 4096 10304 4104 10368
rect 3784 9280 4104 10304
rect 4662 9621 4722 20707
rect 6624 20704 6944 21728
rect 6624 20640 6632 20704
rect 6696 20640 6712 20704
rect 6776 20640 6792 20704
rect 6856 20640 6872 20704
rect 6936 20640 6944 20704
rect 6624 19616 6944 20640
rect 6624 19552 6632 19616
rect 6696 19552 6712 19616
rect 6776 19552 6792 19616
rect 6856 19552 6872 19616
rect 6936 19552 6944 19616
rect 5395 19412 5461 19413
rect 5395 19348 5396 19412
rect 5460 19348 5461 19412
rect 5395 19347 5461 19348
rect 5398 12069 5458 19347
rect 6624 18528 6944 19552
rect 6624 18464 6632 18528
rect 6696 18464 6712 18528
rect 6776 18464 6792 18528
rect 6856 18464 6872 18528
rect 6936 18464 6944 18528
rect 6624 17440 6944 18464
rect 6624 17376 6632 17440
rect 6696 17376 6712 17440
rect 6776 17376 6792 17440
rect 6856 17376 6872 17440
rect 6936 17376 6944 17440
rect 6315 16692 6381 16693
rect 6315 16628 6316 16692
rect 6380 16628 6381 16692
rect 6315 16627 6381 16628
rect 5395 12068 5461 12069
rect 5395 12004 5396 12068
rect 5460 12004 5461 12068
rect 5395 12003 5461 12004
rect 4659 9620 4725 9621
rect 4659 9556 4660 9620
rect 4724 9556 4725 9620
rect 4659 9555 4725 9556
rect 3784 9216 3792 9280
rect 3856 9216 3872 9280
rect 3936 9216 3952 9280
rect 4016 9216 4032 9280
rect 4096 9216 4104 9280
rect 3784 8192 4104 9216
rect 3784 8128 3792 8192
rect 3856 8128 3872 8192
rect 3936 8128 3952 8192
rect 4016 8128 4032 8192
rect 4096 8128 4104 8192
rect 3784 7104 4104 8128
rect 3784 7040 3792 7104
rect 3856 7040 3872 7104
rect 3936 7040 3952 7104
rect 4016 7040 4032 7104
rect 4096 7040 4104 7104
rect 3784 6016 4104 7040
rect 3784 5952 3792 6016
rect 3856 5952 3872 6016
rect 3936 5952 3952 6016
rect 4016 5952 4032 6016
rect 4096 5952 4104 6016
rect 3784 4928 4104 5952
rect 3784 4864 3792 4928
rect 3856 4864 3872 4928
rect 3936 4864 3952 4928
rect 4016 4864 4032 4928
rect 4096 4864 4104 4928
rect 3784 3840 4104 4864
rect 3784 3776 3792 3840
rect 3856 3776 3872 3840
rect 3936 3776 3952 3840
rect 4016 3776 4032 3840
rect 4096 3776 4104 3840
rect 3784 2752 4104 3776
rect 5398 3093 5458 12003
rect 6318 9757 6378 16627
rect 6624 16352 6944 17376
rect 6624 16288 6632 16352
rect 6696 16288 6712 16352
rect 6776 16288 6792 16352
rect 6856 16288 6872 16352
rect 6936 16288 6944 16352
rect 6624 15264 6944 16288
rect 6624 15200 6632 15264
rect 6696 15200 6712 15264
rect 6776 15200 6792 15264
rect 6856 15200 6872 15264
rect 6936 15200 6944 15264
rect 6624 14176 6944 15200
rect 6624 14112 6632 14176
rect 6696 14112 6712 14176
rect 6776 14112 6792 14176
rect 6856 14112 6872 14176
rect 6936 14112 6944 14176
rect 6624 13088 6944 14112
rect 6624 13024 6632 13088
rect 6696 13024 6712 13088
rect 6776 13024 6792 13088
rect 6856 13024 6872 13088
rect 6936 13024 6944 13088
rect 6624 12000 6944 13024
rect 6624 11936 6632 12000
rect 6696 11936 6712 12000
rect 6776 11936 6792 12000
rect 6856 11936 6872 12000
rect 6936 11936 6944 12000
rect 6624 10912 6944 11936
rect 6624 10848 6632 10912
rect 6696 10848 6712 10912
rect 6776 10848 6792 10912
rect 6856 10848 6872 10912
rect 6936 10848 6944 10912
rect 6624 9824 6944 10848
rect 6624 9760 6632 9824
rect 6696 9760 6712 9824
rect 6776 9760 6792 9824
rect 6856 9760 6872 9824
rect 6936 9760 6944 9824
rect 6315 9756 6381 9757
rect 6315 9692 6316 9756
rect 6380 9692 6381 9756
rect 6315 9691 6381 9692
rect 5763 9484 5829 9485
rect 5763 9420 5764 9484
rect 5828 9420 5829 9484
rect 5763 9419 5829 9420
rect 5766 4045 5826 9419
rect 6624 8736 6944 9760
rect 6624 8672 6632 8736
rect 6696 8672 6712 8736
rect 6776 8672 6792 8736
rect 6856 8672 6872 8736
rect 6936 8672 6944 8736
rect 6624 7648 6944 8672
rect 6624 7584 6632 7648
rect 6696 7584 6712 7648
rect 6776 7584 6792 7648
rect 6856 7584 6872 7648
rect 6936 7584 6944 7648
rect 6624 6560 6944 7584
rect 6624 6496 6632 6560
rect 6696 6496 6712 6560
rect 6776 6496 6792 6560
rect 6856 6496 6872 6560
rect 6936 6496 6944 6560
rect 6624 5472 6944 6496
rect 6624 5408 6632 5472
rect 6696 5408 6712 5472
rect 6776 5408 6792 5472
rect 6856 5408 6872 5472
rect 6936 5408 6944 5472
rect 6624 4384 6944 5408
rect 6624 4320 6632 4384
rect 6696 4320 6712 4384
rect 6776 4320 6792 4384
rect 6856 4320 6872 4384
rect 6936 4320 6944 4384
rect 5763 4044 5829 4045
rect 5763 3980 5764 4044
rect 5828 3980 5829 4044
rect 5763 3979 5829 3980
rect 6624 3296 6944 4320
rect 6624 3232 6632 3296
rect 6696 3232 6712 3296
rect 6776 3232 6792 3296
rect 6856 3232 6872 3296
rect 6936 3232 6944 3296
rect 4291 3092 4357 3093
rect 4291 3028 4292 3092
rect 4356 3028 4357 3092
rect 4291 3027 4357 3028
rect 5395 3092 5461 3093
rect 5395 3028 5396 3092
rect 5460 3028 5461 3092
rect 5395 3027 5461 3028
rect 3784 2688 3792 2752
rect 3856 2688 3872 2752
rect 3936 2688 3952 2752
rect 4016 2688 4032 2752
rect 4096 2688 4104 2752
rect 3784 2128 4104 2688
rect 4294 2549 4354 3027
rect 4291 2548 4357 2549
rect 4291 2484 4292 2548
rect 4356 2484 4357 2548
rect 4291 2483 4357 2484
rect 6624 2208 6944 3232
rect 6624 2144 6632 2208
rect 6696 2144 6712 2208
rect 6776 2144 6792 2208
rect 6856 2144 6872 2208
rect 6936 2144 6944 2208
rect 6624 2128 6944 2144
rect 9465 22336 9785 22352
rect 9465 22272 9473 22336
rect 9537 22272 9553 22336
rect 9617 22272 9633 22336
rect 9697 22272 9713 22336
rect 9777 22272 9785 22336
rect 9465 21248 9785 22272
rect 9465 21184 9473 21248
rect 9537 21184 9553 21248
rect 9617 21184 9633 21248
rect 9697 21184 9713 21248
rect 9777 21184 9785 21248
rect 9465 20160 9785 21184
rect 9465 20096 9473 20160
rect 9537 20096 9553 20160
rect 9617 20096 9633 20160
rect 9697 20096 9713 20160
rect 9777 20096 9785 20160
rect 9465 19072 9785 20096
rect 9465 19008 9473 19072
rect 9537 19008 9553 19072
rect 9617 19008 9633 19072
rect 9697 19008 9713 19072
rect 9777 19008 9785 19072
rect 9465 17984 9785 19008
rect 9465 17920 9473 17984
rect 9537 17920 9553 17984
rect 9617 17920 9633 17984
rect 9697 17920 9713 17984
rect 9777 17920 9785 17984
rect 9465 16896 9785 17920
rect 9465 16832 9473 16896
rect 9537 16832 9553 16896
rect 9617 16832 9633 16896
rect 9697 16832 9713 16896
rect 9777 16832 9785 16896
rect 9465 15808 9785 16832
rect 9465 15744 9473 15808
rect 9537 15744 9553 15808
rect 9617 15744 9633 15808
rect 9697 15744 9713 15808
rect 9777 15744 9785 15808
rect 9465 14720 9785 15744
rect 9465 14656 9473 14720
rect 9537 14656 9553 14720
rect 9617 14656 9633 14720
rect 9697 14656 9713 14720
rect 9777 14656 9785 14720
rect 9465 13632 9785 14656
rect 9465 13568 9473 13632
rect 9537 13568 9553 13632
rect 9617 13568 9633 13632
rect 9697 13568 9713 13632
rect 9777 13568 9785 13632
rect 9465 12544 9785 13568
rect 9465 12480 9473 12544
rect 9537 12480 9553 12544
rect 9617 12480 9633 12544
rect 9697 12480 9713 12544
rect 9777 12480 9785 12544
rect 9465 11456 9785 12480
rect 9465 11392 9473 11456
rect 9537 11392 9553 11456
rect 9617 11392 9633 11456
rect 9697 11392 9713 11456
rect 9777 11392 9785 11456
rect 9465 10368 9785 11392
rect 9465 10304 9473 10368
rect 9537 10304 9553 10368
rect 9617 10304 9633 10368
rect 9697 10304 9713 10368
rect 9777 10304 9785 10368
rect 9465 9280 9785 10304
rect 9465 9216 9473 9280
rect 9537 9216 9553 9280
rect 9617 9216 9633 9280
rect 9697 9216 9713 9280
rect 9777 9216 9785 9280
rect 9465 8192 9785 9216
rect 9465 8128 9473 8192
rect 9537 8128 9553 8192
rect 9617 8128 9633 8192
rect 9697 8128 9713 8192
rect 9777 8128 9785 8192
rect 9465 7104 9785 8128
rect 9465 7040 9473 7104
rect 9537 7040 9553 7104
rect 9617 7040 9633 7104
rect 9697 7040 9713 7104
rect 9777 7040 9785 7104
rect 9465 6016 9785 7040
rect 9465 5952 9473 6016
rect 9537 5952 9553 6016
rect 9617 5952 9633 6016
rect 9697 5952 9713 6016
rect 9777 5952 9785 6016
rect 9465 4928 9785 5952
rect 9465 4864 9473 4928
rect 9537 4864 9553 4928
rect 9617 4864 9633 4928
rect 9697 4864 9713 4928
rect 9777 4864 9785 4928
rect 9465 3840 9785 4864
rect 9465 3776 9473 3840
rect 9537 3776 9553 3840
rect 9617 3776 9633 3840
rect 9697 3776 9713 3840
rect 9777 3776 9785 3840
rect 9465 2752 9785 3776
rect 9465 2688 9473 2752
rect 9537 2688 9553 2752
rect 9617 2688 9633 2752
rect 9697 2688 9713 2752
rect 9777 2688 9785 2752
rect 9465 2128 9785 2688
rect 12305 21792 12625 22352
rect 12305 21728 12313 21792
rect 12377 21728 12393 21792
rect 12457 21728 12473 21792
rect 12537 21728 12553 21792
rect 12617 21728 12625 21792
rect 12305 20704 12625 21728
rect 15146 22336 15466 22352
rect 15146 22272 15154 22336
rect 15218 22272 15234 22336
rect 15298 22272 15314 22336
rect 15378 22272 15394 22336
rect 15458 22272 15466 22336
rect 14227 21316 14293 21317
rect 14227 21252 14228 21316
rect 14292 21252 14293 21316
rect 14227 21251 14293 21252
rect 12305 20640 12313 20704
rect 12377 20640 12393 20704
rect 12457 20640 12473 20704
rect 12537 20640 12553 20704
rect 12617 20640 12625 20704
rect 12305 19616 12625 20640
rect 12305 19552 12313 19616
rect 12377 19552 12393 19616
rect 12457 19552 12473 19616
rect 12537 19552 12553 19616
rect 12617 19552 12625 19616
rect 12305 18528 12625 19552
rect 12305 18464 12313 18528
rect 12377 18464 12393 18528
rect 12457 18464 12473 18528
rect 12537 18464 12553 18528
rect 12617 18464 12625 18528
rect 12305 17440 12625 18464
rect 12305 17376 12313 17440
rect 12377 17376 12393 17440
rect 12457 17376 12473 17440
rect 12537 17376 12553 17440
rect 12617 17376 12625 17440
rect 12305 16352 12625 17376
rect 12305 16288 12313 16352
rect 12377 16288 12393 16352
rect 12457 16288 12473 16352
rect 12537 16288 12553 16352
rect 12617 16288 12625 16352
rect 12305 15264 12625 16288
rect 12305 15200 12313 15264
rect 12377 15200 12393 15264
rect 12457 15200 12473 15264
rect 12537 15200 12553 15264
rect 12617 15200 12625 15264
rect 12305 14176 12625 15200
rect 14230 15197 14290 21251
rect 15146 21248 15466 22272
rect 15146 21184 15154 21248
rect 15218 21184 15234 21248
rect 15298 21184 15314 21248
rect 15378 21184 15394 21248
rect 15458 21184 15466 21248
rect 15146 20160 15466 21184
rect 15146 20096 15154 20160
rect 15218 20096 15234 20160
rect 15298 20096 15314 20160
rect 15378 20096 15394 20160
rect 15458 20096 15466 20160
rect 15146 19072 15466 20096
rect 15146 19008 15154 19072
rect 15218 19008 15234 19072
rect 15298 19008 15314 19072
rect 15378 19008 15394 19072
rect 15458 19008 15466 19072
rect 14963 18868 15029 18869
rect 14963 18804 14964 18868
rect 15028 18804 15029 18868
rect 14963 18803 15029 18804
rect 14227 15196 14293 15197
rect 14227 15132 14228 15196
rect 14292 15132 14293 15196
rect 14227 15131 14293 15132
rect 12305 14112 12313 14176
rect 12377 14112 12393 14176
rect 12457 14112 12473 14176
rect 12537 14112 12553 14176
rect 12617 14112 12625 14176
rect 12305 13088 12625 14112
rect 14966 13837 15026 18803
rect 15146 17984 15466 19008
rect 15146 17920 15154 17984
rect 15218 17920 15234 17984
rect 15298 17920 15314 17984
rect 15378 17920 15394 17984
rect 15458 17920 15466 17984
rect 15146 16896 15466 17920
rect 15146 16832 15154 16896
rect 15218 16832 15234 16896
rect 15298 16832 15314 16896
rect 15378 16832 15394 16896
rect 15458 16832 15466 16896
rect 15146 15808 15466 16832
rect 15146 15744 15154 15808
rect 15218 15744 15234 15808
rect 15298 15744 15314 15808
rect 15378 15744 15394 15808
rect 15458 15744 15466 15808
rect 15146 14720 15466 15744
rect 15146 14656 15154 14720
rect 15218 14656 15234 14720
rect 15298 14656 15314 14720
rect 15378 14656 15394 14720
rect 15458 14656 15466 14720
rect 14595 13836 14661 13837
rect 14595 13772 14596 13836
rect 14660 13772 14661 13836
rect 14595 13771 14661 13772
rect 14963 13836 15029 13837
rect 14963 13772 14964 13836
rect 15028 13772 15029 13836
rect 14963 13771 15029 13772
rect 12305 13024 12313 13088
rect 12377 13024 12393 13088
rect 12457 13024 12473 13088
rect 12537 13024 12553 13088
rect 12617 13024 12625 13088
rect 12305 12000 12625 13024
rect 12305 11936 12313 12000
rect 12377 11936 12393 12000
rect 12457 11936 12473 12000
rect 12537 11936 12553 12000
rect 12617 11936 12625 12000
rect 12305 10912 12625 11936
rect 12305 10848 12313 10912
rect 12377 10848 12393 10912
rect 12457 10848 12473 10912
rect 12537 10848 12553 10912
rect 12617 10848 12625 10912
rect 12305 9824 12625 10848
rect 12305 9760 12313 9824
rect 12377 9760 12393 9824
rect 12457 9760 12473 9824
rect 12537 9760 12553 9824
rect 12617 9760 12625 9824
rect 12305 8736 12625 9760
rect 12305 8672 12313 8736
rect 12377 8672 12393 8736
rect 12457 8672 12473 8736
rect 12537 8672 12553 8736
rect 12617 8672 12625 8736
rect 12305 7648 12625 8672
rect 12305 7584 12313 7648
rect 12377 7584 12393 7648
rect 12457 7584 12473 7648
rect 12537 7584 12553 7648
rect 12617 7584 12625 7648
rect 12305 6560 12625 7584
rect 14598 6901 14658 13771
rect 15146 13632 15466 14656
rect 15146 13568 15154 13632
rect 15218 13568 15234 13632
rect 15298 13568 15314 13632
rect 15378 13568 15394 13632
rect 15458 13568 15466 13632
rect 15146 12544 15466 13568
rect 15146 12480 15154 12544
rect 15218 12480 15234 12544
rect 15298 12480 15314 12544
rect 15378 12480 15394 12544
rect 15458 12480 15466 12544
rect 15146 11456 15466 12480
rect 15146 11392 15154 11456
rect 15218 11392 15234 11456
rect 15298 11392 15314 11456
rect 15378 11392 15394 11456
rect 15458 11392 15466 11456
rect 15146 10368 15466 11392
rect 17986 21792 18306 22352
rect 17986 21728 17994 21792
rect 18058 21728 18074 21792
rect 18138 21728 18154 21792
rect 18218 21728 18234 21792
rect 18298 21728 18306 21792
rect 17986 20704 18306 21728
rect 20827 22336 21147 22352
rect 20827 22272 20835 22336
rect 20899 22272 20915 22336
rect 20979 22272 20995 22336
rect 21059 22272 21075 22336
rect 21139 22272 21147 22336
rect 20827 21248 21147 22272
rect 20827 21184 20835 21248
rect 20899 21184 20915 21248
rect 20979 21184 20995 21248
rect 21059 21184 21075 21248
rect 21139 21184 21147 21248
rect 19747 20772 19813 20773
rect 19747 20708 19748 20772
rect 19812 20708 19813 20772
rect 19747 20707 19813 20708
rect 17986 20640 17994 20704
rect 18058 20640 18074 20704
rect 18138 20640 18154 20704
rect 18218 20640 18234 20704
rect 18298 20640 18306 20704
rect 17986 19616 18306 20640
rect 17986 19552 17994 19616
rect 18058 19552 18074 19616
rect 18138 19552 18154 19616
rect 18218 19552 18234 19616
rect 18298 19552 18306 19616
rect 17986 18528 18306 19552
rect 17986 18464 17994 18528
rect 18058 18464 18074 18528
rect 18138 18464 18154 18528
rect 18218 18464 18234 18528
rect 18298 18464 18306 18528
rect 17986 17440 18306 18464
rect 17986 17376 17994 17440
rect 18058 17376 18074 17440
rect 18138 17376 18154 17440
rect 18218 17376 18234 17440
rect 18298 17376 18306 17440
rect 17986 16352 18306 17376
rect 17986 16288 17994 16352
rect 18058 16288 18074 16352
rect 18138 16288 18154 16352
rect 18218 16288 18234 16352
rect 18298 16288 18306 16352
rect 17986 15264 18306 16288
rect 17986 15200 17994 15264
rect 18058 15200 18074 15264
rect 18138 15200 18154 15264
rect 18218 15200 18234 15264
rect 18298 15200 18306 15264
rect 17986 14176 18306 15200
rect 17986 14112 17994 14176
rect 18058 14112 18074 14176
rect 18138 14112 18154 14176
rect 18218 14112 18234 14176
rect 18298 14112 18306 14176
rect 17986 13088 18306 14112
rect 17986 13024 17994 13088
rect 18058 13024 18074 13088
rect 18138 13024 18154 13088
rect 18218 13024 18234 13088
rect 18298 13024 18306 13088
rect 17986 12000 18306 13024
rect 19750 12341 19810 20707
rect 20827 20160 21147 21184
rect 20827 20096 20835 20160
rect 20899 20096 20915 20160
rect 20979 20096 20995 20160
rect 21059 20096 21075 20160
rect 21139 20096 21147 20160
rect 20827 19072 21147 20096
rect 20827 19008 20835 19072
rect 20899 19008 20915 19072
rect 20979 19008 20995 19072
rect 21059 19008 21075 19072
rect 21139 19008 21147 19072
rect 19931 18052 19997 18053
rect 19931 17988 19932 18052
rect 19996 17988 19997 18052
rect 19931 17987 19997 17988
rect 19747 12340 19813 12341
rect 19747 12276 19748 12340
rect 19812 12276 19813 12340
rect 19747 12275 19813 12276
rect 17986 11936 17994 12000
rect 18058 11936 18074 12000
rect 18138 11936 18154 12000
rect 18218 11936 18234 12000
rect 18298 11936 18306 12000
rect 17723 11116 17789 11117
rect 17723 11052 17724 11116
rect 17788 11052 17789 11116
rect 17723 11051 17789 11052
rect 15146 10304 15154 10368
rect 15218 10304 15234 10368
rect 15298 10304 15314 10368
rect 15378 10304 15394 10368
rect 15458 10304 15466 10368
rect 15146 9280 15466 10304
rect 15146 9216 15154 9280
rect 15218 9216 15234 9280
rect 15298 9216 15314 9280
rect 15378 9216 15394 9280
rect 15458 9216 15466 9280
rect 15146 8192 15466 9216
rect 15146 8128 15154 8192
rect 15218 8128 15234 8192
rect 15298 8128 15314 8192
rect 15378 8128 15394 8192
rect 15458 8128 15466 8192
rect 15146 7104 15466 8128
rect 15146 7040 15154 7104
rect 15218 7040 15234 7104
rect 15298 7040 15314 7104
rect 15378 7040 15394 7104
rect 15458 7040 15466 7104
rect 14595 6900 14661 6901
rect 14595 6836 14596 6900
rect 14660 6836 14661 6900
rect 14595 6835 14661 6836
rect 12305 6496 12313 6560
rect 12377 6496 12393 6560
rect 12457 6496 12473 6560
rect 12537 6496 12553 6560
rect 12617 6496 12625 6560
rect 12305 5472 12625 6496
rect 12305 5408 12313 5472
rect 12377 5408 12393 5472
rect 12457 5408 12473 5472
rect 12537 5408 12553 5472
rect 12617 5408 12625 5472
rect 12305 4384 12625 5408
rect 12305 4320 12313 4384
rect 12377 4320 12393 4384
rect 12457 4320 12473 4384
rect 12537 4320 12553 4384
rect 12617 4320 12625 4384
rect 12305 3296 12625 4320
rect 12305 3232 12313 3296
rect 12377 3232 12393 3296
rect 12457 3232 12473 3296
rect 12537 3232 12553 3296
rect 12617 3232 12625 3296
rect 12305 2208 12625 3232
rect 12305 2144 12313 2208
rect 12377 2144 12393 2208
rect 12457 2144 12473 2208
rect 12537 2144 12553 2208
rect 12617 2144 12625 2208
rect 12305 2128 12625 2144
rect 15146 6016 15466 7040
rect 15146 5952 15154 6016
rect 15218 5952 15234 6016
rect 15298 5952 15314 6016
rect 15378 5952 15394 6016
rect 15458 5952 15466 6016
rect 15146 4928 15466 5952
rect 17726 5269 17786 11051
rect 17986 10912 18306 11936
rect 17986 10848 17994 10912
rect 18058 10848 18074 10912
rect 18138 10848 18154 10912
rect 18218 10848 18234 10912
rect 18298 10848 18306 10912
rect 17986 9824 18306 10848
rect 17986 9760 17994 9824
rect 18058 9760 18074 9824
rect 18138 9760 18154 9824
rect 18218 9760 18234 9824
rect 18298 9760 18306 9824
rect 17986 8736 18306 9760
rect 17986 8672 17994 8736
rect 18058 8672 18074 8736
rect 18138 8672 18154 8736
rect 18218 8672 18234 8736
rect 18298 8672 18306 8736
rect 17986 7648 18306 8672
rect 17986 7584 17994 7648
rect 18058 7584 18074 7648
rect 18138 7584 18154 7648
rect 18218 7584 18234 7648
rect 18298 7584 18306 7648
rect 17986 6560 18306 7584
rect 17986 6496 17994 6560
rect 18058 6496 18074 6560
rect 18138 6496 18154 6560
rect 18218 6496 18234 6560
rect 18298 6496 18306 6560
rect 17986 5472 18306 6496
rect 19934 5677 19994 17987
rect 20827 17984 21147 19008
rect 20827 17920 20835 17984
rect 20899 17920 20915 17984
rect 20979 17920 20995 17984
rect 21059 17920 21075 17984
rect 21139 17920 21147 17984
rect 20827 16896 21147 17920
rect 20827 16832 20835 16896
rect 20899 16832 20915 16896
rect 20979 16832 20995 16896
rect 21059 16832 21075 16896
rect 21139 16832 21147 16896
rect 20827 15808 21147 16832
rect 20827 15744 20835 15808
rect 20899 15744 20915 15808
rect 20979 15744 20995 15808
rect 21059 15744 21075 15808
rect 21139 15744 21147 15808
rect 20827 14720 21147 15744
rect 20827 14656 20835 14720
rect 20899 14656 20915 14720
rect 20979 14656 20995 14720
rect 21059 14656 21075 14720
rect 21139 14656 21147 14720
rect 20827 13632 21147 14656
rect 20827 13568 20835 13632
rect 20899 13568 20915 13632
rect 20979 13568 20995 13632
rect 21059 13568 21075 13632
rect 21139 13568 21147 13632
rect 20827 12544 21147 13568
rect 20827 12480 20835 12544
rect 20899 12480 20915 12544
rect 20979 12480 20995 12544
rect 21059 12480 21075 12544
rect 21139 12480 21147 12544
rect 20827 11456 21147 12480
rect 20827 11392 20835 11456
rect 20899 11392 20915 11456
rect 20979 11392 20995 11456
rect 21059 11392 21075 11456
rect 21139 11392 21147 11456
rect 20827 10368 21147 11392
rect 20827 10304 20835 10368
rect 20899 10304 20915 10368
rect 20979 10304 20995 10368
rect 21059 10304 21075 10368
rect 21139 10304 21147 10368
rect 20827 9280 21147 10304
rect 20827 9216 20835 9280
rect 20899 9216 20915 9280
rect 20979 9216 20995 9280
rect 21059 9216 21075 9280
rect 21139 9216 21147 9280
rect 20827 8192 21147 9216
rect 20827 8128 20835 8192
rect 20899 8128 20915 8192
rect 20979 8128 20995 8192
rect 21059 8128 21075 8192
rect 21139 8128 21147 8192
rect 20827 7104 21147 8128
rect 20827 7040 20835 7104
rect 20899 7040 20915 7104
rect 20979 7040 20995 7104
rect 21059 7040 21075 7104
rect 21139 7040 21147 7104
rect 20827 6016 21147 7040
rect 20827 5952 20835 6016
rect 20899 5952 20915 6016
rect 20979 5952 20995 6016
rect 21059 5952 21075 6016
rect 21139 5952 21147 6016
rect 19931 5676 19997 5677
rect 19931 5612 19932 5676
rect 19996 5612 19997 5676
rect 19931 5611 19997 5612
rect 17986 5408 17994 5472
rect 18058 5408 18074 5472
rect 18138 5408 18154 5472
rect 18218 5408 18234 5472
rect 18298 5408 18306 5472
rect 17723 5268 17789 5269
rect 17723 5204 17724 5268
rect 17788 5204 17789 5268
rect 17723 5203 17789 5204
rect 15146 4864 15154 4928
rect 15218 4864 15234 4928
rect 15298 4864 15314 4928
rect 15378 4864 15394 4928
rect 15458 4864 15466 4928
rect 15146 3840 15466 4864
rect 15146 3776 15154 3840
rect 15218 3776 15234 3840
rect 15298 3776 15314 3840
rect 15378 3776 15394 3840
rect 15458 3776 15466 3840
rect 15146 2752 15466 3776
rect 15146 2688 15154 2752
rect 15218 2688 15234 2752
rect 15298 2688 15314 2752
rect 15378 2688 15394 2752
rect 15458 2688 15466 2752
rect 15146 2128 15466 2688
rect 17986 4384 18306 5408
rect 17986 4320 17994 4384
rect 18058 4320 18074 4384
rect 18138 4320 18154 4384
rect 18218 4320 18234 4384
rect 18298 4320 18306 4384
rect 17986 3296 18306 4320
rect 17986 3232 17994 3296
rect 18058 3232 18074 3296
rect 18138 3232 18154 3296
rect 18218 3232 18234 3296
rect 18298 3232 18306 3296
rect 17986 2208 18306 3232
rect 17986 2144 17994 2208
rect 18058 2144 18074 2208
rect 18138 2144 18154 2208
rect 18218 2144 18234 2208
rect 18298 2144 18306 2208
rect 17986 2128 18306 2144
rect 20827 4928 21147 5952
rect 20827 4864 20835 4928
rect 20899 4864 20915 4928
rect 20979 4864 20995 4928
rect 21059 4864 21075 4928
rect 21139 4864 21147 4928
rect 20827 3840 21147 4864
rect 20827 3776 20835 3840
rect 20899 3776 20915 3840
rect 20979 3776 20995 3840
rect 21059 3776 21075 3840
rect 21139 3776 21147 3840
rect 20827 2752 21147 3776
rect 20827 2688 20835 2752
rect 20899 2688 20915 2752
rect 20979 2688 20995 2752
rect 21059 2688 21075 2752
rect 21139 2688 21147 2752
rect 20827 2128 21147 2688
rect 23667 21792 23987 22352
rect 23667 21728 23675 21792
rect 23739 21728 23755 21792
rect 23819 21728 23835 21792
rect 23899 21728 23915 21792
rect 23979 21728 23987 21792
rect 23667 20704 23987 21728
rect 23667 20640 23675 20704
rect 23739 20640 23755 20704
rect 23819 20640 23835 20704
rect 23899 20640 23915 20704
rect 23979 20640 23987 20704
rect 23667 19616 23987 20640
rect 23667 19552 23675 19616
rect 23739 19552 23755 19616
rect 23819 19552 23835 19616
rect 23899 19552 23915 19616
rect 23979 19552 23987 19616
rect 23667 18528 23987 19552
rect 23667 18464 23675 18528
rect 23739 18464 23755 18528
rect 23819 18464 23835 18528
rect 23899 18464 23915 18528
rect 23979 18464 23987 18528
rect 23667 17440 23987 18464
rect 23667 17376 23675 17440
rect 23739 17376 23755 17440
rect 23819 17376 23835 17440
rect 23899 17376 23915 17440
rect 23979 17376 23987 17440
rect 23667 16352 23987 17376
rect 23667 16288 23675 16352
rect 23739 16288 23755 16352
rect 23819 16288 23835 16352
rect 23899 16288 23915 16352
rect 23979 16288 23987 16352
rect 23667 15264 23987 16288
rect 23667 15200 23675 15264
rect 23739 15200 23755 15264
rect 23819 15200 23835 15264
rect 23899 15200 23915 15264
rect 23979 15200 23987 15264
rect 23667 14176 23987 15200
rect 23667 14112 23675 14176
rect 23739 14112 23755 14176
rect 23819 14112 23835 14176
rect 23899 14112 23915 14176
rect 23979 14112 23987 14176
rect 23667 13088 23987 14112
rect 23667 13024 23675 13088
rect 23739 13024 23755 13088
rect 23819 13024 23835 13088
rect 23899 13024 23915 13088
rect 23979 13024 23987 13088
rect 23667 12000 23987 13024
rect 23667 11936 23675 12000
rect 23739 11936 23755 12000
rect 23819 11936 23835 12000
rect 23899 11936 23915 12000
rect 23979 11936 23987 12000
rect 23667 10912 23987 11936
rect 23667 10848 23675 10912
rect 23739 10848 23755 10912
rect 23819 10848 23835 10912
rect 23899 10848 23915 10912
rect 23979 10848 23987 10912
rect 23667 9824 23987 10848
rect 23667 9760 23675 9824
rect 23739 9760 23755 9824
rect 23819 9760 23835 9824
rect 23899 9760 23915 9824
rect 23979 9760 23987 9824
rect 23667 8736 23987 9760
rect 23667 8672 23675 8736
rect 23739 8672 23755 8736
rect 23819 8672 23835 8736
rect 23899 8672 23915 8736
rect 23979 8672 23987 8736
rect 23667 7648 23987 8672
rect 23667 7584 23675 7648
rect 23739 7584 23755 7648
rect 23819 7584 23835 7648
rect 23899 7584 23915 7648
rect 23979 7584 23987 7648
rect 23667 6560 23987 7584
rect 23667 6496 23675 6560
rect 23739 6496 23755 6560
rect 23819 6496 23835 6560
rect 23899 6496 23915 6560
rect 23979 6496 23987 6560
rect 23667 5472 23987 6496
rect 23667 5408 23675 5472
rect 23739 5408 23755 5472
rect 23819 5408 23835 5472
rect 23899 5408 23915 5472
rect 23979 5408 23987 5472
rect 23667 4384 23987 5408
rect 23667 4320 23675 4384
rect 23739 4320 23755 4384
rect 23819 4320 23835 4384
rect 23899 4320 23915 4384
rect 23979 4320 23987 4384
rect 23667 3296 23987 4320
rect 23667 3232 23675 3296
rect 23739 3232 23755 3296
rect 23819 3232 23835 3296
rect 23899 3232 23915 3296
rect 23979 3232 23987 3296
rect 23667 2208 23987 3232
rect 23667 2144 23675 2208
rect 23739 2144 23755 2208
rect 23819 2144 23835 2208
rect 23899 2144 23915 2208
rect 23979 2144 23987 2208
rect 23667 2128 23987 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1676037725
transform -1 0 20976 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__A
timestamp 1676037725
transform 1 0 16100 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A
timestamp 1676037725
transform 1 0 5152 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__C
timestamp 1676037725
transform 1 0 3496 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__391__A
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A
timestamp 1676037725
transform -1 0 15272 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__B
timestamp 1676037725
transform 1 0 16376 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__D
timestamp 1676037725
transform 1 0 10488 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__A
timestamp 1676037725
transform -1 0 20792 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__A0
timestamp 1676037725
transform 1 0 18768 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A2
timestamp 1676037725
transform 1 0 8464 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__A2
timestamp 1676037725
transform -1 0 1748 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A2
timestamp 1676037725
transform 1 0 5704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__B1
timestamp 1676037725
transform 1 0 13616 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__A
timestamp 1676037725
transform 1 0 5888 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__A
timestamp 1676037725
transform 1 0 18768 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__B1
timestamp 1676037725
transform 1 0 17940 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__B1
timestamp 1676037725
transform 1 0 17940 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__441__A
timestamp 1676037725
transform 1 0 15088 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__A
timestamp 1676037725
transform 1 0 15916 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__A
timestamp 1676037725
transform 1 0 13156 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__449__B1
timestamp 1676037725
transform 1 0 9292 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__A1
timestamp 1676037725
transform 1 0 12972 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__B1
timestamp 1676037725
transform 1 0 11684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__A1
timestamp 1676037725
transform -1 0 14352 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__B1
timestamp 1676037725
transform 1 0 14352 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__458__A1
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__463__B1
timestamp 1676037725
transform 1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__A
timestamp 1676037725
transform -1 0 11224 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__B
timestamp 1676037725
transform -1 0 21436 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__471__A
timestamp 1676037725
transform 1 0 19504 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__B
timestamp 1676037725
transform 1 0 19412 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__A
timestamp 1676037725
transform 1 0 14812 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__A
timestamp 1676037725
transform 1 0 13616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__A
timestamp 1676037725
transform 1 0 16652 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__A
timestamp 1676037725
transform 1 0 16836 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__B
timestamp 1676037725
transform 1 0 18676 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__A1
timestamp 1676037725
transform 1 0 14996 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__A2
timestamp 1676037725
transform 1 0 15272 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__B1
timestamp 1676037725
transform 1 0 15548 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__A
timestamp 1676037725
transform 1 0 22724 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__B
timestamp 1676037725
transform 1 0 22908 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__A
timestamp 1676037725
transform 1 0 11040 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__506__A2
timestamp 1676037725
transform 1 0 20792 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__C
timestamp 1676037725
transform 1 0 19320 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__513__A1
timestamp 1676037725
transform 1 0 15364 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__514__B
timestamp 1676037725
transform 1 0 17848 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__A2
timestamp 1676037725
transform 1 0 18768 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__517__A
timestamp 1676037725
transform 1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__B1
timestamp 1676037725
transform 1 0 22724 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__C1
timestamp 1676037725
transform 1 0 21344 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__523__A
timestamp 1676037725
transform 1 0 20884 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__A
timestamp 1676037725
transform 1 0 21804 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__A2
timestamp 1676037725
transform 1 0 20976 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__529__S
timestamp 1676037725
transform 1 0 14536 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__535__A2
timestamp 1676037725
transform 1 0 20516 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__535__B2
timestamp 1676037725
transform 1 0 18768 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__537__C1
timestamp 1676037725
transform 1 0 20516 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__539__A1
timestamp 1676037725
transform 1 0 13064 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__539__B1
timestamp 1676037725
transform 1 0 15640 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__540__A3
timestamp 1676037725
transform 1 0 13432 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__541__A
timestamp 1676037725
transform 1 0 16836 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__541__B
timestamp 1676037725
transform -1 0 15732 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__C1
timestamp 1676037725
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__553__A2
timestamp 1676037725
transform 1 0 21344 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__555__B1
timestamp 1676037725
transform -1 0 23368 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__557__A1
timestamp 1676037725
transform 1 0 21344 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__557__C1
timestamp 1676037725
transform 1 0 20792 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__560__A1
timestamp 1676037725
transform 1 0 19596 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__560__C1
timestamp 1676037725
transform 1 0 19044 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__564__B
timestamp 1676037725
transform 1 0 18400 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__565__A
timestamp 1676037725
transform 1 0 16100 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__566__A
timestamp 1676037725
transform -1 0 20424 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__567__B1
timestamp 1676037725
transform 1 0 19320 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__568__A1
timestamp 1676037725
transform 1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__573__A
timestamp 1676037725
transform 1 0 13064 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__573__B
timestamp 1676037725
transform 1 0 12512 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__574__A1
timestamp 1676037725
transform 1 0 19320 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__577__A
timestamp 1676037725
transform 1 0 15824 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__579__A1
timestamp 1676037725
transform 1 0 14996 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__583__A
timestamp 1676037725
transform -1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__584__A
timestamp 1676037725
transform 1 0 18492 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__587__B1
timestamp 1676037725
transform 1 0 11684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__590__C1
timestamp 1676037725
transform 1 0 15824 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__591__A1
timestamp 1676037725
transform 1 0 17848 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__591__C1
timestamp 1676037725
transform -1 0 17572 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__593__A
timestamp 1676037725
transform 1 0 12788 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__595__A
timestamp 1676037725
transform 1 0 16100 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__598__C1
timestamp 1676037725
transform 1 0 14260 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__599__A1
timestamp 1676037725
transform 1 0 13340 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__601__C1
timestamp 1676037725
transform 1 0 19228 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__602__A1
timestamp 1676037725
transform 1 0 11408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__603__B1
timestamp 1676037725
transform -1 0 14444 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__605__B1
timestamp 1676037725
transform 1 0 12236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__608__B2
timestamp 1676037725
transform 1 0 15824 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__610__A
timestamp 1676037725
transform -1 0 15180 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__612__B2
timestamp 1676037725
transform 1 0 18952 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__617__A1
timestamp 1676037725
transform 1 0 15548 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__622__A2
timestamp 1676037725
transform -1 0 15456 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__622__B1
timestamp 1676037725
transform 1 0 15916 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__624__A1
timestamp 1676037725
transform -1 0 15548 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__624__B1
timestamp 1676037725
transform 1 0 16192 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__629__A1
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__630__S
timestamp 1676037725
transform 1 0 13156 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__641__A1_N
timestamp 1676037725
transform 1 0 14628 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__647__B1
timestamp 1676037725
transform 1 0 9108 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__660__A
timestamp 1676037725
transform 1 0 8464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__661__B2
timestamp 1676037725
transform 1 0 8004 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__662__S
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__667__A1
timestamp 1676037725
transform 1 0 16836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__667__A2
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__669__C1
timestamp 1676037725
transform -1 0 17020 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__672__A1
timestamp 1676037725
transform 1 0 10212 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__673__A1
timestamp 1676037725
transform 1 0 11040 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__674__A1
timestamp 1676037725
transform 1 0 10028 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__675__S
timestamp 1676037725
transform 1 0 11040 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__678__A
timestamp 1676037725
transform 1 0 13064 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__678__B
timestamp 1676037725
transform 1 0 13432 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__679__A1
timestamp 1676037725
transform 1 0 9384 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__680__A
timestamp 1676037725
transform 1 0 10488 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__681__C1
timestamp 1676037725
transform 1 0 7360 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__687__A1
timestamp 1676037725
transform 1 0 6808 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__693__A1
timestamp 1676037725
transform -1 0 9292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__699__A1
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__700__A1
timestamp 1676037725
transform 1 0 10948 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__702__A1
timestamp 1676037725
transform 1 0 7360 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__703__B2
timestamp 1676037725
transform 1 0 6256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__707__B1
timestamp 1676037725
transform 1 0 6716 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__712__A
timestamp 1676037725
transform 1 0 6808 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__716__A3
timestamp 1676037725
transform -1 0 5060 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__722__A3
timestamp 1676037725
transform 1 0 3772 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__729__A1
timestamp 1676037725
transform 1 0 7268 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__732__S
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__746__D
timestamp 1676037725
transform 1 0 11040 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__748__D
timestamp 1676037725
transform -1 0 8556 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__749__D
timestamp 1676037725
transform 1 0 11224 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__750__D
timestamp 1676037725
transform 1 0 10028 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__751__D
timestamp 1676037725
transform 1 0 10028 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__752__D
timestamp 1676037725
transform 1 0 8464 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__798__A
timestamp 1676037725
transform -1 0 11868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1676037725
transform 1 0 5796 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout16_A
timestamp 1676037725
transform 1 0 22816 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout17_A
timestamp 1676037725
transform -1 0 23092 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout20_A
timestamp 1676037725
transform -1 0 20792 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout24_A
timestamp 1676037725
transform -1 0 22356 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout31_A
timestamp 1676037725
transform 1 0 3956 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1676037725
transform -1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1676037725
transform -1 0 17112 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform -1 0 22448 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform -1 0 7176 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output6_A
timestamp 1676037725
transform -1 0 1748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output8_A
timestamp 1676037725
transform 1 0 4324 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output10_A
timestamp 1676037725
transform -1 0 12420 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output11_A
timestamp 1676037725
transform 1 0 11040 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output12_A
timestamp 1676037725
transform -1 0 1748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42
timestamp 1676037725
transform 1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46
timestamp 1676037725
transform 1 0 5336 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65
timestamp 1676037725
transform 1 0 7084 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71
timestamp 1676037725
transform 1 0 7636 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1676037725
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1676037725
transform 1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1676037725
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1676037725
transform 1 0 10580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1676037725
transform 1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_127
timestamp 1676037725
transform 1 0 12788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134
timestamp 1676037725
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_146 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14536 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1676037725
transform 1 0 15272 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1676037725
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1676037725
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_178
timestamp 1676037725
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_185
timestamp 1676037725
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1676037725
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1676037725
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_216
timestamp 1676037725
transform 1 0 20976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1676037725
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_237
timestamp 1676037725
transform 1 0 22908 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_243
timestamp 1676037725
transform 1 0 23460 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_8
timestamp 1676037725
transform 1 0 1840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_21
timestamp 1676037725
transform 1 0 3036 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_37
timestamp 1676037725
transform 1 0 4508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_50
timestamp 1676037725
transform 1 0 5704 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_72
timestamp 1676037725
transform 1 0 7728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_80
timestamp 1676037725
transform 1 0 8464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_99
timestamp 1676037725
transform 1 0 10212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106
timestamp 1676037725
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_124
timestamp 1676037725
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_128
timestamp 1676037725
transform 1 0 12880 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_135
timestamp 1676037725
transform 1 0 13524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_141
timestamp 1676037725
transform 1 0 14076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1676037725
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_179
timestamp 1676037725
transform 1 0 17572 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_183
timestamp 1676037725
transform 1 0 17940 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_206
timestamp 1676037725
transform 1 0 20056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1676037725
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_230
timestamp 1676037725
transform 1 0 22264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1676037725
transform 1 0 23460 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1676037725
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_17
timestamp 1676037725
transform 1 0 2668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1676037725
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_37
timestamp 1676037725
transform 1 0 4508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_55
timestamp 1676037725
transform 1 0 6164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_76
timestamp 1676037725
transform 1 0 8096 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1676037725
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_92
timestamp 1676037725
transform 1 0 9568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_102
timestamp 1676037725
transform 1 0 10488 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_114
timestamp 1676037725
transform 1 0 11592 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_122
timestamp 1676037725
transform 1 0 12328 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_131
timestamp 1676037725
transform 1 0 13156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_146
timestamp 1676037725
transform 1 0 14536 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_160
timestamp 1676037725
transform 1 0 15824 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_167
timestamp 1676037725
transform 1 0 16468 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_173
timestamp 1676037725
transform 1 0 17020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_179
timestamp 1676037725
transform 1 0 17572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_185
timestamp 1676037725
transform 1 0 18124 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_191
timestamp 1676037725
transform 1 0 18676 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1676037725
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_208
timestamp 1676037725
transform 1 0 20240 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_214 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20792 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_226
timestamp 1676037725
transform 1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_232
timestamp 1676037725
transform 1 0 22448 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_239
timestamp 1676037725
transform 1 0 23092 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_243
timestamp 1676037725
transform 1 0 23460 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1676037725
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_24
timestamp 1676037725
transform 1 0 3312 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_32
timestamp 1676037725
transform 1 0 4048 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_43
timestamp 1676037725
transform 1 0 5060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1676037725
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_75
timestamp 1676037725
transform 1 0 8004 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_79
timestamp 1676037725
transform 1 0 8372 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_89
timestamp 1676037725
transform 1 0 9292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_96
timestamp 1676037725
transform 1 0 9936 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_103
timestamp 1676037725
transform 1 0 10580 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1676037725
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_117
timestamp 1676037725
transform 1 0 11868 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_123
timestamp 1676037725
transform 1 0 12420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_135
timestamp 1676037725
transform 1 0 13524 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_138
timestamp 1676037725
transform 1 0 13800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_144
timestamp 1676037725
transform 1 0 14352 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_154
timestamp 1676037725
transform 1 0 15272 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_173
timestamp 1676037725
transform 1 0 17020 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_185
timestamp 1676037725
transform 1 0 18124 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_206
timestamp 1676037725
transform 1 0 20056 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_218
timestamp 1676037725
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_236
timestamp 1676037725
transform 1 0 22816 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1676037725
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_52
timestamp 1676037725
transform 1 0 5888 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_70
timestamp 1676037725
transform 1 0 7544 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_89
timestamp 1676037725
transform 1 0 9292 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_98
timestamp 1676037725
transform 1 0 10120 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_104
timestamp 1676037725
transform 1 0 10672 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_110
timestamp 1676037725
transform 1 0 11224 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_118
timestamp 1676037725
transform 1 0 11960 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_125
timestamp 1676037725
transform 1 0 12604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1676037725
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1676037725
transform 1 0 14444 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_162
timestamp 1676037725
transform 1 0 16008 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_168
timestamp 1676037725
transform 1 0 16560 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_183
timestamp 1676037725
transform 1 0 17940 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_191
timestamp 1676037725
transform 1 0 18676 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1676037725
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_204
timestamp 1676037725
transform 1 0 19872 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_210
timestamp 1676037725
transform 1 0 20424 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_216
timestamp 1676037725
transform 1 0 20976 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_228
timestamp 1676037725
transform 1 0 22080 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_239
timestamp 1676037725
transform 1 0 23092 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_243
timestamp 1676037725
transform 1 0 23460 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_9
timestamp 1676037725
transform 1 0 1932 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_17
timestamp 1676037725
transform 1 0 2668 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_29
timestamp 1676037725
transform 1 0 3772 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_44
timestamp 1676037725
transform 1 0 5152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1676037725
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_62
timestamp 1676037725
transform 1 0 6808 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_70
timestamp 1676037725
transform 1 0 7544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_84
timestamp 1676037725
transform 1 0 8832 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_97
timestamp 1676037725
transform 1 0 10028 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1676037725
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_121
timestamp 1676037725
transform 1 0 12236 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_130
timestamp 1676037725
transform 1 0 13064 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_136
timestamp 1676037725
transform 1 0 13616 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_146
timestamp 1676037725
transform 1 0 14536 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_150
timestamp 1676037725
transform 1 0 14904 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_159
timestamp 1676037725
transform 1 0 15732 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1676037725
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_173
timestamp 1676037725
transform 1 0 17020 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_179
timestamp 1676037725
transform 1 0 17572 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_192
timestamp 1676037725
transform 1 0 18768 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_196
timestamp 1676037725
transform 1 0 19136 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_204
timestamp 1676037725
transform 1 0 19872 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_208
timestamp 1676037725
transform 1 0 20240 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_212
timestamp 1676037725
transform 1 0 20608 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_216
timestamp 1676037725
transform 1 0 20976 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1676037725
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_231
timestamp 1676037725
transform 1 0 22356 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_241
timestamp 1676037725
transform 1 0 23276 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_7
timestamp 1676037725
transform 1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_18
timestamp 1676037725
transform 1 0 2760 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_22
timestamp 1676037725
transform 1 0 3128 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1676037725
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_36
timestamp 1676037725
transform 1 0 4416 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_56
timestamp 1676037725
transform 1 0 6256 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_67
timestamp 1676037725
transform 1 0 7268 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1676037725
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_89
timestamp 1676037725
transform 1 0 9292 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_104
timestamp 1676037725
transform 1 0 10672 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_116
timestamp 1676037725
transform 1 0 11776 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_129
timestamp 1676037725
transform 1 0 12972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1676037725
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_158
timestamp 1676037725
transform 1 0 15640 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_164
timestamp 1676037725
transform 1 0 16192 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_169
timestamp 1676037725
transform 1 0 16652 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_187
timestamp 1676037725
transform 1 0 18308 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_202
timestamp 1676037725
transform 1 0 19688 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1676037725
transform 1 0 20884 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_231
timestamp 1676037725
transform 1 0 22356 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_241
timestamp 1676037725
transform 1 0 23276 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_9
timestamp 1676037725
transform 1 0 1932 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_34
timestamp 1676037725
transform 1 0 4232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_47
timestamp 1676037725
transform 1 0 5428 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1676037725
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_62
timestamp 1676037725
transform 1 0 6808 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_89
timestamp 1676037725
transform 1 0 9292 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_101
timestamp 1676037725
transform 1 0 10396 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 1676037725
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_117
timestamp 1676037725
transform 1 0 11868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_126
timestamp 1676037725
transform 1 0 12696 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_132
timestamp 1676037725
transform 1 0 13248 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_142
timestamp 1676037725
transform 1 0 14168 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_146
timestamp 1676037725
transform 1 0 14536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_185
timestamp 1676037725
transform 1 0 18124 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_198
timestamp 1676037725
transform 1 0 19320 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_211
timestamp 1676037725
transform 1 0 20516 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_215
timestamp 1676037725
transform 1 0 20884 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1676037725
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_233
timestamp 1676037725
transform 1 0 22540 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_242
timestamp 1676037725
transform 1 0 23368 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_16
timestamp 1676037725
transform 1 0 2576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 1676037725
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_63
timestamp 1676037725
transform 1 0 6900 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_67
timestamp 1676037725
transform 1 0 7268 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_70
timestamp 1676037725
transform 1 0 7544 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1676037725
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_89
timestamp 1676037725
transform 1 0 9292 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_92
timestamp 1676037725
transform 1 0 9568 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_103
timestamp 1676037725
transform 1 0 10580 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_111
timestamp 1676037725
transform 1 0 11316 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_118
timestamp 1676037725
transform 1 0 11960 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_130
timestamp 1676037725
transform 1 0 13064 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1676037725
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_149
timestamp 1676037725
transform 1 0 14812 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_155
timestamp 1676037725
transform 1 0 15364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_167
timestamp 1676037725
transform 1 0 16468 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_171
timestamp 1676037725
transform 1 0 16836 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_175
timestamp 1676037725
transform 1 0 17204 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_188
timestamp 1676037725
transform 1 0 18400 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1676037725
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_213
timestamp 1676037725
transform 1 0 20700 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_225
timestamp 1676037725
transform 1 0 21804 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_236
timestamp 1676037725
transform 1 0 22816 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_11
timestamp 1676037725
transform 1 0 2116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_21
timestamp 1676037725
transform 1 0 3036 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_31
timestamp 1676037725
transform 1 0 3956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_41
timestamp 1676037725
transform 1 0 4876 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1676037725
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_65
timestamp 1676037725
transform 1 0 7084 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_73
timestamp 1676037725
transform 1 0 7820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_80
timestamp 1676037725
transform 1 0 8464 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_92
timestamp 1676037725
transform 1 0 9568 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_101
timestamp 1676037725
transform 1 0 10396 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_107
timestamp 1676037725
transform 1 0 10948 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1676037725
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_117
timestamp 1676037725
transform 1 0 11868 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_121
timestamp 1676037725
transform 1 0 12236 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_127
timestamp 1676037725
transform 1 0 12788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_139
timestamp 1676037725
transform 1 0 13892 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_146
timestamp 1676037725
transform 1 0 14536 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_157
timestamp 1676037725
transform 1 0 15548 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1676037725
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_180
timestamp 1676037725
transform 1 0 17664 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_188
timestamp 1676037725
transform 1 0 18400 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_207
timestamp 1676037725
transform 1 0 20148 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_219
timestamp 1676037725
transform 1 0 21252 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_239
timestamp 1676037725
transform 1 0 23092 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_243
timestamp 1676037725
transform 1 0 23460 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_14
timestamp 1676037725
transform 1 0 2392 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1676037725
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_33
timestamp 1676037725
transform 1 0 4140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_51
timestamp 1676037725
transform 1 0 5796 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_55
timestamp 1676037725
transform 1 0 6164 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_67
timestamp 1676037725
transform 1 0 7268 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_71
timestamp 1676037725
transform 1 0 7636 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_94
timestamp 1676037725
transform 1 0 9752 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_113
timestamp 1676037725
transform 1 0 11500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_131
timestamp 1676037725
transform 1 0 13156 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_135
timestamp 1676037725
transform 1 0 13524 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_148
timestamp 1676037725
transform 1 0 14720 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1676037725
transform 1 0 15272 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_163
timestamp 1676037725
transform 1 0 16100 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_184
timestamp 1676037725
transform 1 0 18032 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1676037725
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_208
timestamp 1676037725
transform 1 0 20240 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_218
timestamp 1676037725
transform 1 0 21160 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_226
timestamp 1676037725
transform 1 0 21896 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_231
timestamp 1676037725
transform 1 0 22356 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_237
timestamp 1676037725
transform 1 0 22908 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_243
timestamp 1676037725
transform 1 0 23460 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1676037725
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_17
timestamp 1676037725
transform 1 0 2668 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_28
timestamp 1676037725
transform 1 0 3680 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_40
timestamp 1676037725
transform 1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_46
timestamp 1676037725
transform 1 0 5336 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1676037725
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_68
timestamp 1676037725
transform 1 0 7360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_80
timestamp 1676037725
transform 1 0 8464 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_88
timestamp 1676037725
transform 1 0 9200 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_91
timestamp 1676037725
transform 1 0 9476 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_102
timestamp 1676037725
transform 1 0 10488 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_106
timestamp 1676037725
transform 1 0 10856 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1676037725
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1676037725
transform 1 0 11868 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_131
timestamp 1676037725
transform 1 0 13156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_160
timestamp 1676037725
transform 1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_173
timestamp 1676037725
transform 1 0 17020 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_200
timestamp 1676037725
transform 1 0 19504 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_212
timestamp 1676037725
transform 1 0 20608 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_218
timestamp 1676037725
transform 1 0 21160 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_235
timestamp 1676037725
transform 1 0 22724 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_243
timestamp 1676037725
transform 1 0 23460 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1676037725
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_11
timestamp 1676037725
transform 1 0 2116 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1676037725
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_37
timestamp 1676037725
transform 1 0 4508 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_47
timestamp 1676037725
transform 1 0 5428 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_55
timestamp 1676037725
transform 1 0 6164 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_98
timestamp 1676037725
transform 1 0 10120 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_106
timestamp 1676037725
transform 1 0 10856 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_120
timestamp 1676037725
transform 1 0 12144 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_127
timestamp 1676037725
transform 1 0 12788 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1676037725
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_157
timestamp 1676037725
transform 1 0 15548 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_163
timestamp 1676037725
transform 1 0 16100 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_176
timestamp 1676037725
transform 1 0 17296 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_187
timestamp 1676037725
transform 1 0 18308 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_193
timestamp 1676037725
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_201
timestamp 1676037725
transform 1 0 19596 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_205
timestamp 1676037725
transform 1 0 19964 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_213
timestamp 1676037725
transform 1 0 20700 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_224
timestamp 1676037725
transform 1 0 21712 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_236
timestamp 1676037725
transform 1 0 22816 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_242
timestamp 1676037725
transform 1 0 23368 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_7
timestamp 1676037725
transform 1 0 1748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_17
timestamp 1676037725
transform 1 0 2668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_24
timestamp 1676037725
transform 1 0 3312 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_28
timestamp 1676037725
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_31
timestamp 1676037725
transform 1 0 3956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_37
timestamp 1676037725
transform 1 0 4508 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_49
timestamp 1676037725
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_63
timestamp 1676037725
transform 1 0 6900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_70
timestamp 1676037725
transform 1 0 7544 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_83
timestamp 1676037725
transform 1 0 8740 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_95
timestamp 1676037725
transform 1 0 9844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_104
timestamp 1676037725
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_118
timestamp 1676037725
transform 1 0 11960 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_138
timestamp 1676037725
transform 1 0 13800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_147
timestamp 1676037725
transform 1 0 14628 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_156
timestamp 1676037725
transform 1 0 15456 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_162
timestamp 1676037725
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_180
timestamp 1676037725
transform 1 0 17664 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_189
timestamp 1676037725
transform 1 0 18492 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_201
timestamp 1676037725
transform 1 0 19596 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_210
timestamp 1676037725
transform 1 0 20424 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_216
timestamp 1676037725
transform 1 0 20976 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_233
timestamp 1676037725
transform 1 0 22540 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_241
timestamp 1676037725
transform 1 0 23276 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1676037725
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_13
timestamp 1676037725
transform 1 0 2300 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_19
timestamp 1676037725
transform 1 0 2852 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1676037725
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_38
timestamp 1676037725
transform 1 0 4600 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_49
timestamp 1676037725
transform 1 0 5612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_58
timestamp 1676037725
transform 1 0 6440 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_64
timestamp 1676037725
transform 1 0 6992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_70
timestamp 1676037725
transform 1 0 7544 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_78
timestamp 1676037725
transform 1 0 8280 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1676037725
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_95
timestamp 1676037725
transform 1 0 9844 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_101
timestamp 1676037725
transform 1 0 10396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_127
timestamp 1676037725
transform 1 0 12788 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_152
timestamp 1676037725
transform 1 0 15088 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_161
timestamp 1676037725
transform 1 0 15916 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_173
timestamp 1676037725
transform 1 0 17020 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_179
timestamp 1676037725
transform 1 0 17572 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_183
timestamp 1676037725
transform 1 0 17940 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1676037725
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_212
timestamp 1676037725
transform 1 0 20608 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_224
timestamp 1676037725
transform 1 0 21712 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_236
timestamp 1676037725
transform 1 0 22816 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_13
timestamp 1676037725
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_22
timestamp 1676037725
transform 1 0 3128 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_28
timestamp 1676037725
transform 1 0 3680 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_38
timestamp 1676037725
transform 1 0 4600 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_46
timestamp 1676037725
transform 1 0 5336 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1676037725
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_68
timestamp 1676037725
transform 1 0 7360 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_75
timestamp 1676037725
transform 1 0 8004 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_83
timestamp 1676037725
transform 1 0 8740 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_89
timestamp 1676037725
transform 1 0 9292 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_98
timestamp 1676037725
transform 1 0 10120 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_104
timestamp 1676037725
transform 1 0 10672 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1676037725
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_122
timestamp 1676037725
transform 1 0 12328 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_162
timestamp 1676037725
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_179
timestamp 1676037725
transform 1 0 17572 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_194
timestamp 1676037725
transform 1 0 18952 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_200
timestamp 1676037725
transform 1 0 19504 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_212
timestamp 1676037725
transform 1 0 20608 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_234
timestamp 1676037725
transform 1 0 22632 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_242
timestamp 1676037725
transform 1 0 23368 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1676037725
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_38
timestamp 1676037725
transform 1 0 4600 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_50
timestamp 1676037725
transform 1 0 5704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1676037725
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_93
timestamp 1676037725
transform 1 0 9660 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_99
timestamp 1676037725
transform 1 0 10212 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_111
timestamp 1676037725
transform 1 0 11316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_120
timestamp 1676037725
transform 1 0 12144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_126
timestamp 1676037725
transform 1 0 12696 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_132
timestamp 1676037725
transform 1 0 13248 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1676037725
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_145
timestamp 1676037725
transform 1 0 14444 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_157
timestamp 1676037725
transform 1 0 15548 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1676037725
transform 1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_170
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_178
timestamp 1676037725
transform 1 0 17480 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_184
timestamp 1676037725
transform 1 0 18032 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1676037725
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_207
timestamp 1676037725
transform 1 0 20148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_219
timestamp 1676037725
transform 1 0 21252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_227
timestamp 1676037725
transform 1 0 21988 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_238
timestamp 1676037725
transform 1 0 23000 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_36
timestamp 1676037725
transform 1 0 4416 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1676037725
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_67
timestamp 1676037725
transform 1 0 7268 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_77
timestamp 1676037725
transform 1 0 8188 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_89
timestamp 1676037725
transform 1 0 9292 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1676037725
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_127
timestamp 1676037725
transform 1 0 12788 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_145
timestamp 1676037725
transform 1 0 14444 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_159
timestamp 1676037725
transform 1 0 15732 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 1676037725
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_178
timestamp 1676037725
transform 1 0 17480 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_184
timestamp 1676037725
transform 1 0 18032 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_190
timestamp 1676037725
transform 1 0 18584 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_200
timestamp 1676037725
transform 1 0 19504 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_212
timestamp 1676037725
transform 1 0 20608 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_218
timestamp 1676037725
transform 1 0 21160 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_231
timestamp 1676037725
transform 1 0 22356 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_237
timestamp 1676037725
transform 1 0 22908 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_243
timestamp 1676037725
transform 1 0 23460 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_10
timestamp 1676037725
transform 1 0 2024 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_19
timestamp 1676037725
transform 1 0 2852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_37
timestamp 1676037725
transform 1 0 4508 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_43
timestamp 1676037725
transform 1 0 5060 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_55
timestamp 1676037725
transform 1 0 6164 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_58
timestamp 1676037725
transform 1 0 6440 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_64
timestamp 1676037725
transform 1 0 6992 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_71
timestamp 1676037725
transform 1 0 7636 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1676037725
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_96
timestamp 1676037725
transform 1 0 9936 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_107
timestamp 1676037725
transform 1 0 10948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_113
timestamp 1676037725
transform 1 0 11500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_126
timestamp 1676037725
transform 1 0 12696 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp 1676037725
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_150
timestamp 1676037725
transform 1 0 14904 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_163
timestamp 1676037725
transform 1 0 16100 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_175
timestamp 1676037725
transform 1 0 17204 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_186
timestamp 1676037725
transform 1 0 18216 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_201
timestamp 1676037725
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_210
timestamp 1676037725
transform 1 0 20424 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_216
timestamp 1676037725
transform 1 0 20976 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_225
timestamp 1676037725
transform 1 0 21804 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_234
timestamp 1676037725
transform 1 0 22632 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_241
timestamp 1676037725
transform 1 0 23276 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1676037725
transform 1 0 1748 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_14
timestamp 1676037725
transform 1 0 2392 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_22
timestamp 1676037725
transform 1 0 3128 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_34
timestamp 1676037725
transform 1 0 4232 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_40
timestamp 1676037725
transform 1 0 4784 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1676037725
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_65
timestamp 1676037725
transform 1 0 7084 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_77
timestamp 1676037725
transform 1 0 8188 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_85
timestamp 1676037725
transform 1 0 8924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_91
timestamp 1676037725
transform 1 0 9476 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1676037725
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_122
timestamp 1676037725
transform 1 0 12328 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_131
timestamp 1676037725
transform 1 0 13156 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_144
timestamp 1676037725
transform 1 0 14352 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_151
timestamp 1676037725
transform 1 0 14996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_155
timestamp 1676037725
transform 1 0 15364 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1676037725
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_179
timestamp 1676037725
transform 1 0 17572 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_194
timestamp 1676037725
transform 1 0 18952 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_200
timestamp 1676037725
transform 1 0 19504 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_212
timestamp 1676037725
transform 1 0 20608 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_233
timestamp 1676037725
transform 1 0 22540 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_239
timestamp 1676037725
transform 1 0 23092 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_243
timestamp 1676037725
transform 1 0 23460 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_11
timestamp 1676037725
transform 1 0 2116 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_19
timestamp 1676037725
transform 1 0 2852 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1676037725
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_35
timestamp 1676037725
transform 1 0 4324 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_48
timestamp 1676037725
transform 1 0 5520 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_57
timestamp 1676037725
transform 1 0 6348 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_63
timestamp 1676037725
transform 1 0 6900 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_67
timestamp 1676037725
transform 1 0 7268 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_71
timestamp 1676037725
transform 1 0 7636 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1676037725
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_98
timestamp 1676037725
transform 1 0 10120 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_107
timestamp 1676037725
transform 1 0 10948 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_119
timestamp 1676037725
transform 1 0 12052 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_123
timestamp 1676037725
transform 1 0 12420 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_128
timestamp 1676037725
transform 1 0 12880 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_150
timestamp 1676037725
transform 1 0 14904 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_156
timestamp 1676037725
transform 1 0 15456 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_162
timestamp 1676037725
transform 1 0 16008 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_172
timestamp 1676037725
transform 1 0 16928 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_184
timestamp 1676037725
transform 1 0 18032 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_206
timestamp 1676037725
transform 1 0 20056 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_214
timestamp 1676037725
transform 1 0 20792 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_222
timestamp 1676037725
transform 1 0 21528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_232
timestamp 1676037725
transform 1 0 22448 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_238
timestamp 1676037725
transform 1 0 23000 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_35
timestamp 1676037725
transform 1 0 4324 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_41
timestamp 1676037725
transform 1 0 4876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1676037725
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_67
timestamp 1676037725
transform 1 0 7268 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_75
timestamp 1676037725
transform 1 0 8004 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_92
timestamp 1676037725
transform 1 0 9568 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_104
timestamp 1676037725
transform 1 0 10672 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_118
timestamp 1676037725
transform 1 0 11960 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_126
timestamp 1676037725
transform 1 0 12696 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_129
timestamp 1676037725
transform 1 0 12972 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_147
timestamp 1676037725
transform 1 0 14628 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1676037725
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_159
timestamp 1676037725
transform 1 0 15732 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1676037725
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_178
timestamp 1676037725
transform 1 0 17480 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_190
timestamp 1676037725
transform 1 0 18584 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_202
timestamp 1676037725
transform 1 0 19688 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_211
timestamp 1676037725
transform 1 0 20516 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_236
timestamp 1676037725
transform 1 0 22816 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_14
timestamp 1676037725
transform 1 0 2392 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1676037725
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_38
timestamp 1676037725
transform 1 0 4600 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_42
timestamp 1676037725
transform 1 0 4968 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_50
timestamp 1676037725
transform 1 0 5704 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_61
timestamp 1676037725
transform 1 0 6716 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_69
timestamp 1676037725
transform 1 0 7452 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_78
timestamp 1676037725
transform 1 0 8280 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_94
timestamp 1676037725
transform 1 0 9752 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_109
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_127
timestamp 1676037725
transform 1 0 12788 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_135
timestamp 1676037725
transform 1 0 13524 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_145
timestamp 1676037725
transform 1 0 14444 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_151
timestamp 1676037725
transform 1 0 14996 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_157
timestamp 1676037725
transform 1 0 15548 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_162
timestamp 1676037725
transform 1 0 16008 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_174
timestamp 1676037725
transform 1 0 17112 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_186
timestamp 1676037725
transform 1 0 18216 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_191
timestamp 1676037725
transform 1 0 18676 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_207
timestamp 1676037725
transform 1 0 20148 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_217
timestamp 1676037725
transform 1 0 21068 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_231
timestamp 1676037725
transform 1 0 22356 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_238
timestamp 1676037725
transform 1 0 23000 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1676037725
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_40
timestamp 1676037725
transform 1 0 4784 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1676037725
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_63
timestamp 1676037725
transform 1 0 6900 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_103
timestamp 1676037725
transform 1 0 10580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_124
timestamp 1676037725
transform 1 0 12512 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_136
timestamp 1676037725
transform 1 0 13616 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_142
timestamp 1676037725
transform 1 0 14168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_150
timestamp 1676037725
transform 1 0 14904 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_158
timestamp 1676037725
transform 1 0 15640 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_178
timestamp 1676037725
transform 1 0 17480 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_189
timestamp 1676037725
transform 1 0 18492 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_202
timestamp 1676037725
transform 1 0 19688 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_216
timestamp 1676037725
transform 1 0 20976 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1676037725
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_237
timestamp 1676037725
transform 1 0 22908 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_243
timestamp 1676037725
transform 1 0 23460 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_51
timestamp 1676037725
transform 1 0 5796 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_59
timestamp 1676037725
transform 1 0 6532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_104
timestamp 1676037725
transform 1 0 10672 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_110
timestamp 1676037725
transform 1 0 11224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_114
timestamp 1676037725
transform 1 0 11592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_117
timestamp 1676037725
transform 1 0 11868 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_127
timestamp 1676037725
transform 1 0 12788 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_154
timestamp 1676037725
transform 1 0 15272 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_164
timestamp 1676037725
transform 1 0 16192 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_172
timestamp 1676037725
transform 1 0 16928 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_181
timestamp 1676037725
transform 1 0 17756 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_206
timestamp 1676037725
transform 1 0 20056 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_214
timestamp 1676037725
transform 1 0 20792 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_221
timestamp 1676037725
transform 1 0 21436 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_231
timestamp 1676037725
transform 1 0 22356 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_243
timestamp 1676037725
transform 1 0 23460 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_36
timestamp 1676037725
transform 1 0 4416 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_48
timestamp 1676037725
transform 1 0 5520 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1676037725
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_142
timestamp 1676037725
transform 1 0 14168 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_148
timestamp 1676037725
transform 1 0 14720 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_154
timestamp 1676037725
transform 1 0 15272 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_162
timestamp 1676037725
transform 1 0 16008 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_175
timestamp 1676037725
transform 1 0 17204 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_182
timestamp 1676037725
transform 1 0 17848 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_190
timestamp 1676037725
transform 1 0 18584 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_194
timestamp 1676037725
transform 1 0 18952 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_197
timestamp 1676037725
transform 1 0 19228 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_203
timestamp 1676037725
transform 1 0 19780 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_214
timestamp 1676037725
transform 1 0 20792 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_233
timestamp 1676037725
transform 1 0 22540 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_239
timestamp 1676037725
transform 1 0 23092 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_243
timestamp 1676037725
transform 1 0 23460 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_9
timestamp 1676037725
transform 1 0 1932 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1676037725
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_47
timestamp 1676037725
transform 1 0 5428 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_59
timestamp 1676037725
transform 1 0 6532 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp 1676037725
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_106
timestamp 1676037725
transform 1 0 10856 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_112
timestamp 1676037725
transform 1 0 11408 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_120
timestamp 1676037725
transform 1 0 12144 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_129
timestamp 1676037725
transform 1 0 12972 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_135
timestamp 1676037725
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_145
timestamp 1676037725
transform 1 0 14444 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_151
timestamp 1676037725
transform 1 0 14996 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_157
timestamp 1676037725
transform 1 0 15548 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_163
timestamp 1676037725
transform 1 0 16100 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_171
timestamp 1676037725
transform 1 0 16836 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_179
timestamp 1676037725
transform 1 0 17572 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_186
timestamp 1676037725
transform 1 0 18216 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_207
timestamp 1676037725
transform 1 0 20148 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_213
timestamp 1676037725
transform 1 0 20700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_225
timestamp 1676037725
transform 1 0 21804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_231
timestamp 1676037725
transform 1 0 22356 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_243
timestamp 1676037725
transform 1 0 23460 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_19
timestamp 1676037725
transform 1 0 2852 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_75
timestamp 1676037725
transform 1 0 8004 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_79
timestamp 1676037725
transform 1 0 8372 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_96
timestamp 1676037725
transform 1 0 9936 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1676037725
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_123
timestamp 1676037725
transform 1 0 12420 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_134
timestamp 1676037725
transform 1 0 13432 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_141
timestamp 1676037725
transform 1 0 14076 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_145
timestamp 1676037725
transform 1 0 14444 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_154
timestamp 1676037725
transform 1 0 15272 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_160
timestamp 1676037725
transform 1 0 15824 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_176
timestamp 1676037725
transform 1 0 17296 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_188
timestamp 1676037725
transform 1 0 18400 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_196
timestamp 1676037725
transform 1 0 19136 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_206
timestamp 1676037725
transform 1 0 20056 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_216
timestamp 1676037725
transform 1 0 20976 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_233
timestamp 1676037725
transform 1 0 22540 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_241
timestamp 1676037725
transform 1 0 23276 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_66
timestamp 1676037725
transform 1 0 7176 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_78
timestamp 1676037725
transform 1 0 8280 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_81
timestamp 1676037725
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_103
timestamp 1676037725
transform 1 0 10580 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_107
timestamp 1676037725
transform 1 0 10948 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_110
timestamp 1676037725
transform 1 0 11224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_117
timestamp 1676037725
transform 1 0 11868 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_127
timestamp 1676037725
transform 1 0 12788 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_145
timestamp 1676037725
transform 1 0 14444 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_152
timestamp 1676037725
transform 1 0 15088 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_162
timestamp 1676037725
transform 1 0 16008 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_172
timestamp 1676037725
transform 1 0 16928 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_181
timestamp 1676037725
transform 1 0 17756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1676037725
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1676037725
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_223
timestamp 1676037725
transform 1 0 21620 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_235
timestamp 1676037725
transform 1 0 22724 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_243
timestamp 1676037725
transform 1 0 23460 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_37
timestamp 1676037725
transform 1 0 4508 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_49
timestamp 1676037725
transform 1 0 5612 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_126
timestamp 1676037725
transform 1 0 12696 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_132
timestamp 1676037725
transform 1 0 13248 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_142
timestamp 1676037725
transform 1 0 14168 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_154
timestamp 1676037725
transform 1 0 15272 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_160
timestamp 1676037725
transform 1 0 15824 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1676037725
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_178
timestamp 1676037725
transform 1 0 17480 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_188
timestamp 1676037725
transform 1 0 18400 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_196
timestamp 1676037725
transform 1 0 19136 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_206
timestamp 1676037725
transform 1 0 20056 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_218
timestamp 1676037725
transform 1 0 21160 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_243
timestamp 1676037725
transform 1 0 23460 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_9
timestamp 1676037725
transform 1 0 1932 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1676037725
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_49
timestamp 1676037725
transform 1 0 5612 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_103
timestamp 1676037725
transform 1 0 10580 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_115
timestamp 1676037725
transform 1 0 11684 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_123
timestamp 1676037725
transform 1 0 12420 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_151
timestamp 1676037725
transform 1 0 14996 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_157
timestamp 1676037725
transform 1 0 15548 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_172
timestamp 1676037725
transform 1 0 16928 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_184
timestamp 1676037725
transform 1 0 18032 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_207
timestamp 1676037725
transform 1 0 20148 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_213
timestamp 1676037725
transform 1 0 20700 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_225
timestamp 1676037725
transform 1 0 21804 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_237
timestamp 1676037725
transform 1 0 22908 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_243
timestamp 1676037725
transform 1 0 23460 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_19
timestamp 1676037725
transform 1 0 2852 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_93
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_99
timestamp 1676037725
transform 1 0 10212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_121
timestamp 1676037725
transform 1 0 12236 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_130
timestamp 1676037725
transform 1 0 13064 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_136
timestamp 1676037725
transform 1 0 13616 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_144
timestamp 1676037725
transform 1 0 14352 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_149
timestamp 1676037725
transform 1 0 14812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_153
timestamp 1676037725
transform 1 0 15180 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_156
timestamp 1676037725
transform 1 0 15456 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_162
timestamp 1676037725
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_180
timestamp 1676037725
transform 1 0 17664 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_190
timestamp 1676037725
transform 1 0 18584 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_204
timestamp 1676037725
transform 1 0 19872 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_216
timestamp 1676037725
transform 1 0 20976 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_232
timestamp 1676037725
transform 1 0 22448 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_9
timestamp 1676037725
transform 1 0 1932 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1676037725
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_45
timestamp 1676037725
transform 1 0 5244 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_62
timestamp 1676037725
transform 1 0 6808 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1676037725
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_106
timestamp 1676037725
transform 1 0 10856 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_114
timestamp 1676037725
transform 1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_126
timestamp 1676037725
transform 1 0 12696 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_130
timestamp 1676037725
transform 1 0 13064 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_135
timestamp 1676037725
transform 1 0 13524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1676037725
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_147
timestamp 1676037725
transform 1 0 14628 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_153
timestamp 1676037725
transform 1 0 15180 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_159
timestamp 1676037725
transform 1 0 15732 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_171
timestamp 1676037725
transform 1 0 16836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_183
timestamp 1676037725
transform 1 0 17940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1676037725
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_205
timestamp 1676037725
transform 1 0 19964 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_217
timestamp 1676037725
transform 1 0 21068 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_229
timestamp 1676037725
transform 1 0 22172 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_241
timestamp 1676037725
transform 1 0 23276 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_36
timestamp 1676037725
transform 1 0 4416 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_48
timestamp 1676037725
transform 1 0 5520 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_93
timestamp 1676037725
transform 1 0 9660 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_99
timestamp 1676037725
transform 1 0 10212 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_107
timestamp 1676037725
transform 1 0 10948 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_119
timestamp 1676037725
transform 1 0 12052 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_129
timestamp 1676037725
transform 1 0 12972 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_139
timestamp 1676037725
transform 1 0 13892 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_146
timestamp 1676037725
transform 1 0 14536 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_157
timestamp 1676037725
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1676037725
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1676037725
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_193
timestamp 1676037725
transform 1 0 18860 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_199
timestamp 1676037725
transform 1 0 19412 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_208
timestamp 1676037725
transform 1 0 20240 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_214
timestamp 1676037725
transform 1 0 20792 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_230
timestamp 1676037725
transform 1 0 22264 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_237
timestamp 1676037725
transform 1 0 22908 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_243
timestamp 1676037725
transform 1 0 23460 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1676037725
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_49
timestamp 1676037725
transform 1 0 5612 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_67
timestamp 1676037725
transform 1 0 7268 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_79
timestamp 1676037725
transform 1 0 8372 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1676037725
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_103
timestamp 1676037725
transform 1 0 10580 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_114
timestamp 1676037725
transform 1 0 11592 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_121
timestamp 1676037725
transform 1 0 12236 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_135
timestamp 1676037725
transform 1 0 13524 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1676037725
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1676037725
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_151
timestamp 1676037725
transform 1 0 14996 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_165
timestamp 1676037725
transform 1 0 16284 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_173
timestamp 1676037725
transform 1 0 17020 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_182
timestamp 1676037725
transform 1 0 17848 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_191
timestamp 1676037725
transform 1 0 18676 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1676037725
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_206
timestamp 1676037725
transform 1 0 20056 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_216
timestamp 1676037725
transform 1 0 20976 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_224
timestamp 1676037725
transform 1 0 21712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_239
timestamp 1676037725
transform 1 0 23092 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_243
timestamp 1676037725
transform 1 0 23460 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_34
timestamp 1676037725
transform 1 0 4232 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1676037725
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_75
timestamp 1676037725
transform 1 0 8004 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_95
timestamp 1676037725
transform 1 0 9844 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_107
timestamp 1676037725
transform 1 0 10948 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1676037725
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_119
timestamp 1676037725
transform 1 0 12052 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_127
timestamp 1676037725
transform 1 0 12788 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_133
timestamp 1676037725
transform 1 0 13340 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_143
timestamp 1676037725
transform 1 0 14260 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_150
timestamp 1676037725
transform 1 0 14904 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_158
timestamp 1676037725
transform 1 0 15640 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_173
timestamp 1676037725
transform 1 0 17020 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_177
timestamp 1676037725
transform 1 0 17388 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_186
timestamp 1676037725
transform 1 0 18216 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_198
timestamp 1676037725
transform 1 0 19320 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_202
timestamp 1676037725
transform 1 0 19688 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_209
timestamp 1676037725
transform 1 0 20332 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_218
timestamp 1676037725
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_229
timestamp 1676037725
transform 1 0 22172 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_232
timestamp 1676037725
transform 1 0 22448 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_9
timestamp 1676037725
transform 1 0 1932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1676037725
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_57
timestamp 1676037725
transform 1 0 6348 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_63
timestamp 1676037725
transform 1 0 6900 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_66
timestamp 1676037725
transform 1 0 7176 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_76
timestamp 1676037725
transform 1 0 8096 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_109
timestamp 1676037725
transform 1 0 11132 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_113
timestamp 1676037725
transform 1 0 11500 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_117
timestamp 1676037725
transform 1 0 11868 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_124
timestamp 1676037725
transform 1 0 12512 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_132
timestamp 1676037725
transform 1 0 13248 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1676037725
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_145
timestamp 1676037725
transform 1 0 14444 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_153
timestamp 1676037725
transform 1 0 15180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_159
timestamp 1676037725
transform 1 0 15732 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_167
timestamp 1676037725
transform 1 0 16468 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_169
timestamp 1676037725
transform 1 0 16652 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_174
timestamp 1676037725
transform 1 0 17112 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_182
timestamp 1676037725
transform 1 0 17848 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1676037725
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_209
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_213
timestamp 1676037725
transform 1 0 20700 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_221
timestamp 1676037725
transform 1 0 21436 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_225
timestamp 1676037725
transform 1 0 21804 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_231
timestamp 1676037725
transform 1 0 22356 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_236
timestamp 1676037725
transform 1 0 22816 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 23828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 23828 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 23828 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 23828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 23828 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 23828 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 23828 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 23828 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 23828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 23828 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 23828 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 23828 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 23828 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 23828 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 23828 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 23828 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 23828 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 23828 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 23828 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 23828 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 23828 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 23828 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 23828 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 23828 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 23828 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 23828 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 23828 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 23828 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 23828 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 23828 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 23828 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 23828 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 23828 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 23828 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 6256 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 11408 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 16560 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 21712 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__inv_6  _369_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4968 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _370_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4232 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1676037725
transform 1 0 3220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1676037725
transform 1 0 10948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1676037725
transform 1 0 14260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1676037725
transform -1 0 20608 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _375_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16652 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_8  _376_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8096 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_4  _377_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5428 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _378_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2944 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _379_
timestamp 1676037725
transform 1 0 4416 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _380_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2668 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_4  _381_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__or3_4  _382_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4600 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _383_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4416 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _384_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5428 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _385_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2300 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _386_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3036 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_4  _387_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4784 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_4  _388_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_2  _389_
timestamp 1676037725
transform 1 0 1840 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand4b_4  _390_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 10880
box -38 -48 1786 592
use sky130_fd_sc_hd__nor3_4  _391_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10948 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _392_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _393_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9016 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _394_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3496 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _395_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2392 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _396_
timestamp 1676037725
transform -1 0 2116 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _397_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _398_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3588 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_1  _399_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16008 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_4  _400_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2668 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_1  _401_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2300 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _402_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_4  _403_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _404_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4048 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _405_
timestamp 1676037725
transform 1 0 20424 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _406_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _407_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2668 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _408_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_4  _409_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4784 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _410_
timestamp 1676037725
transform 1 0 11960 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_4  _411_
timestamp 1676037725
transform 1 0 9108 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_4  _412_
timestamp 1676037725
transform 1 0 6256 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__xor2_4  _413_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8464 0 1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _414_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _415_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7084 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _416_
timestamp 1676037725
transform 1 0 4508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _417_
timestamp 1676037725
transform 1 0 6532 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _418_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5980 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_4  _419_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6900 0 1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _420_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6256 0 1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__a31o_4  _421_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1326 592
use sky130_fd_sc_hd__o221a_2  _422_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2208 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _423_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8832 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _424_
timestamp 1676037725
transform -1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _425_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4508 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_2  _426_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7452 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__o311ai_4  _427_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14168 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__nor3_4  _428_
timestamp 1676037725
transform 1 0 6532 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__or4_2  _429_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _430_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _431_
timestamp 1676037725
transform 1 0 6532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _432_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4968 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _433_
timestamp 1676037725
transform 1 0 8096 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_4  _434_
timestamp 1676037725
transform -1 0 5704 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _435_
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _436_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18768 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a41oi_4  _437_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18032 0 -1 3264
box -38 -48 2062 592
use sky130_fd_sc_hd__a41o_4  _438_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18492 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _439_
timestamp 1676037725
transform 1 0 14260 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _440_
timestamp 1676037725
transform 1 0 15088 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _441_
timestamp 1676037725
transform -1 0 14720 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _442_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15640 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _443_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14996 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _444_
timestamp 1676037725
transform 1 0 14168 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _445_
timestamp 1676037725
transform -1 0 17572 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_4  _446_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13708 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__nor3_2  _447_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11316 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _448_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7268 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _449_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10488 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _450_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12604 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _451_
timestamp 1676037725
transform -1 0 15180 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _452_
timestamp 1676037725
transform 1 0 14812 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _453_
timestamp 1676037725
transform 1 0 14260 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _454_
timestamp 1676037725
transform -1 0 12788 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _455_
timestamp 1676037725
transform 1 0 12880 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _456_
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_4  _457_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14812 0 -1 8704
box -38 -48 1326 592
use sky130_fd_sc_hd__a31o_2  _458_
timestamp 1676037725
transform -1 0 15548 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _459_
timestamp 1676037725
transform -1 0 13800 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_4  _460_
timestamp 1676037725
transform -1 0 18124 0 -1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _461_
timestamp 1676037725
transform -1 0 20240 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_4  _462_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17664 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_4  _463_
timestamp 1676037725
transform -1 0 15548 0 1 8704
box -38 -48 1326 592
use sky130_fd_sc_hd__o211a_4  _464_
timestamp 1676037725
transform -1 0 18308 0 1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_8  _465_
timestamp 1676037725
transform 1 0 18676 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _466_
timestamp 1676037725
transform 1 0 11592 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _467_
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _468_
timestamp 1676037725
transform 1 0 19688 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_4  _469_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16468 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__and3_1  _470_
timestamp 1676037725
transform -1 0 18860 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _471_
timestamp 1676037725
transform 1 0 20056 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_4  _472_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20700 0 1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__a2bb2o_4  _473_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17388 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_2  _474_
timestamp 1676037725
transform -1 0 18492 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _475_
timestamp 1676037725
transform 1 0 15180 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _476_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13800 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _477_
timestamp 1676037725
transform 1 0 22080 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _478_
timestamp 1676037725
transform 1 0 10764 0 1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _479_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12144 0 -1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _480_
timestamp 1676037725
transform 1 0 19228 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _481_
timestamp 1676037725
transform -1 0 23000 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_4  _482_
timestamp 1676037725
transform 1 0 13156 0 -1 11968
box -38 -48 1326 592
use sky130_fd_sc_hd__a21oi_2  _483_
timestamp 1676037725
transform -1 0 17480 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _484_
timestamp 1676037725
transform 1 0 13800 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _485_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _486_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _487_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19780 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o211ai_1  _488_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17572 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _489_
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _490_
timestamp 1676037725
transform -1 0 10948 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _491_
timestamp 1676037725
transform 1 0 12696 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _492_
timestamp 1676037725
transform -1 0 12236 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _493_
timestamp 1676037725
transform 1 0 16836 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _494_
timestamp 1676037725
transform 1 0 16376 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _495_
timestamp 1676037725
transform 1 0 18492 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _496_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16100 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_4  _497_
timestamp 1676037725
transform 1 0 13340 0 -1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_2  _498_
timestamp 1676037725
transform 1 0 22172 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _499_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20056 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _500_
timestamp 1676037725
transform -1 0 16928 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _501_
timestamp 1676037725
transform -1 0 11960 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _502_
timestamp 1676037725
transform -1 0 12788 0 1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _503_
timestamp 1676037725
transform 1 0 11316 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_2  _504_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18860 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _505_
timestamp 1676037725
transform 1 0 21804 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _506_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 21712 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _507_
timestamp 1676037725
transform -1 0 23000 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _508_
timestamp 1676037725
transform 1 0 23000 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _509_
timestamp 1676037725
transform 1 0 17020 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _510_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19504 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _511_
timestamp 1676037725
transform 1 0 19688 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _512_
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _513_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15272 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and4_2  _514_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14996 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _515_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18400 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_1  _516_
timestamp 1676037725
transform 1 0 15732 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _517_
timestamp 1676037725
transform -1 0 14996 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _518_
timestamp 1676037725
transform -1 0 22816 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _519_
timestamp 1676037725
transform -1 0 22356 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _520_
timestamp 1676037725
transform -1 0 23092 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _521_
timestamp 1676037725
transform -1 0 23092 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _522_
timestamp 1676037725
transform -1 0 22540 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _523_
timestamp 1676037725
transform -1 0 21528 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _524_
timestamp 1676037725
transform 1 0 22080 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _525_
timestamp 1676037725
transform -1 0 21804 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _526_
timestamp 1676037725
transform -1 0 21712 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _527_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22172 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _528_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _529_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14444 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _530_
timestamp 1676037725
transform 1 0 21896 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _531_
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _532_
timestamp 1676037725
transform -1 0 20976 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _533_
timestamp 1676037725
transform -1 0 17756 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _534_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20148 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _535_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _536_
timestamp 1676037725
transform -1 0 18676 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _537_
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _538_
timestamp 1676037725
transform 1 0 17020 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _539_
timestamp 1676037725
transform 1 0 13156 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _540_
timestamp 1676037725
transform -1 0 13064 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _541_
timestamp 1676037725
transform -1 0 14904 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_2  _542_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12604 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _543_
timestamp 1676037725
transform 1 0 21620 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _544_
timestamp 1676037725
transform 1 0 19228 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _545_
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _546_
timestamp 1676037725
transform -1 0 22724 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _547_
timestamp 1676037725
transform -1 0 20240 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_2  _548_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15364 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _549_
timestamp 1676037725
transform -1 0 19596 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _550_
timestamp 1676037725
transform -1 0 21528 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _551_
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _552_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _553_
timestamp 1676037725
transform -1 0 22632 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _554_
timestamp 1676037725
transform 1 0 21988 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _555_
timestamp 1676037725
transform 1 0 22080 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _556_
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _557_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 22908 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _558_
timestamp 1676037725
transform -1 0 21160 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _559_
timestamp 1676037725
transform -1 0 20516 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _560_
timestamp 1676037725
transform -1 0 20792 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _561_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _562_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _563_
timestamp 1676037725
transform -1 0 17480 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _564_
timestamp 1676037725
transform -1 0 16376 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _565_
timestamp 1676037725
transform 1 0 15456 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _566_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 19872 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _567_
timestamp 1676037725
transform 1 0 18308 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _568_
timestamp 1676037725
transform 1 0 13064 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _569_
timestamp 1676037725
transform 1 0 16836 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _570_
timestamp 1676037725
transform -1 0 17204 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _571_
timestamp 1676037725
transform -1 0 18216 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _572_
timestamp 1676037725
transform 1 0 17848 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _573_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11592 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _574_
timestamp 1676037725
transform 1 0 18308 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _575_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16376 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _576_
timestamp 1676037725
transform -1 0 20056 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _577_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _578_
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _579_
timestamp 1676037725
transform 1 0 14444 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _580_
timestamp 1676037725
transform 1 0 20792 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _581_
timestamp 1676037725
transform 1 0 20056 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _582_
timestamp 1676037725
transform 1 0 15364 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _583_
timestamp 1676037725
transform -1 0 15916 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _584_
timestamp 1676037725
transform -1 0 18492 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _585_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16008 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _586_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 22816 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _587_
timestamp 1676037725
transform 1 0 13156 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _588_
timestamp 1676037725
transform 1 0 12052 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _589_
timestamp 1676037725
transform -1 0 16376 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _590_
timestamp 1676037725
transform 1 0 14076 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _591_
timestamp 1676037725
transform 1 0 14812 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_1  _592_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13524 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _593_
timestamp 1676037725
transform -1 0 12880 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _594_
timestamp 1676037725
transform -1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _595_
timestamp 1676037725
transform -1 0 14996 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _596_
timestamp 1676037725
transform -1 0 18584 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _597_
timestamp 1676037725
transform -1 0 18216 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _598_
timestamp 1676037725
transform 1 0 12788 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _599_
timestamp 1676037725
transform 1 0 12328 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _600_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21068 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _601_
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _602_
timestamp 1676037725
transform 1 0 11960 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _603_
timestamp 1676037725
transform 1 0 11960 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _604_
timestamp 1676037725
transform -1 0 12788 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _605_
timestamp 1676037725
transform -1 0 12788 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _606_
timestamp 1676037725
transform -1 0 13340 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _607_
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _608_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15272 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _609_
timestamp 1676037725
transform -1 0 14536 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _610_
timestamp 1676037725
transform 1 0 14536 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _611_
timestamp 1676037725
transform -1 0 20056 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _612_
timestamp 1676037725
transform 1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _613_
timestamp 1676037725
transform 1 0 19320 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _614_
timestamp 1676037725
transform 1 0 19504 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _615_
timestamp 1676037725
transform 1 0 17112 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _616_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16376 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _617_
timestamp 1676037725
transform 1 0 14904 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _618_
timestamp 1676037725
transform -1 0 18952 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _619_
timestamp 1676037725
transform -1 0 17848 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _620_
timestamp 1676037725
transform 1 0 17020 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _621_
timestamp 1676037725
transform 1 0 16376 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _622_
timestamp 1676037725
transform 1 0 15456 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _623_
timestamp 1676037725
transform 1 0 15364 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _624_
timestamp 1676037725
transform -1 0 14168 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _625_
timestamp 1676037725
transform 1 0 14352 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _626_
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _627_
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _628_
timestamp 1676037725
transform 1 0 17480 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _629_
timestamp 1676037725
transform 1 0 13524 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _630_
timestamp 1676037725
transform 1 0 12144 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _631_
timestamp 1676037725
transform 1 0 20700 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _632_
timestamp 1676037725
transform -1 0 20700 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _633_
timestamp 1676037725
transform -1 0 22908 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _634_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 23092 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_1  _635_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 19320 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_4  _636_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9844 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _637_
timestamp 1676037725
transform -1 0 13800 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _638_
timestamp 1676037725
transform 1 0 7820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _639_
timestamp 1676037725
transform -1 0 17940 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _640_
timestamp 1676037725
transform -1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _641_
timestamp 1676037725
transform 1 0 15180 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _642_
timestamp 1676037725
transform -1 0 15732 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _643_
timestamp 1676037725
transform -1 0 8648 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _644_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10028 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _645_
timestamp 1676037725
transform 1 0 7728 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _646_
timestamp 1676037725
transform -1 0 9292 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _647_
timestamp 1676037725
transform -1 0 8464 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _648_
timestamp 1676037725
transform -1 0 10396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _649_
timestamp 1676037725
transform -1 0 11040 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _650_
timestamp 1676037725
transform 1 0 13616 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _651_
timestamp 1676037725
transform 1 0 12328 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _652_
timestamp 1676037725
transform -1 0 10948 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _653_
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _654_
timestamp 1676037725
transform -1 0 2668 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _655_
timestamp 1676037725
transform 1 0 3036 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _656_
timestamp 1676037725
transform -1 0 8464 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _657_
timestamp 1676037725
transform 1 0 7728 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _658_
timestamp 1676037725
transform -1 0 7544 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _659_
timestamp 1676037725
transform -1 0 8740 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _660_
timestamp 1676037725
transform 1 0 8832 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _661_
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_4  _662_
timestamp 1676037725
transform 1 0 11592 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_2  _663_
timestamp 1676037725
transform -1 0 5888 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _664_
timestamp 1676037725
transform 1 0 8004 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _665_
timestamp 1676037725
transform 1 0 9108 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _666_
timestamp 1676037725
transform -1 0 11132 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _667_
timestamp 1676037725
transform 1 0 16928 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _668_
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _669_
timestamp 1676037725
transform 1 0 15640 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _670_
timestamp 1676037725
transform 1 0 13248 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _671_
timestamp 1676037725
transform -1 0 13156 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _672_
timestamp 1676037725
transform -1 0 9844 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _673_
timestamp 1676037725
transform -1 0 12328 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _674_
timestamp 1676037725
transform -1 0 10488 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _675_
timestamp 1676037725
transform 1 0 10304 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _676_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10856 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _677_
timestamp 1676037725
transform 1 0 9384 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _678_
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _679_
timestamp 1676037725
transform 1 0 9936 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _680_
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _681_
timestamp 1676037725
transform 1 0 7912 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _682_
timestamp 1676037725
transform -1 0 9568 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _683_
timestamp 1676037725
transform 1 0 10212 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _684_
timestamp 1676037725
transform 1 0 2668 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _685_
timestamp 1676037725
transform 1 0 3956 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _686_
timestamp 1676037725
transform -1 0 7084 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _687_
timestamp 1676037725
transform 1 0 5428 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _688_
timestamp 1676037725
transform 1 0 5152 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _689_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12972 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _690_
timestamp 1676037725
transform 1 0 11684 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _691_
timestamp 1676037725
transform 1 0 12512 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _692_
timestamp 1676037725
transform 1 0 11684 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _693_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 9660 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _694_
timestamp 1676037725
transform 1 0 12420 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _695_
timestamp 1676037725
transform -1 0 13064 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _696_
timestamp 1676037725
transform 1 0 11408 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _697_
timestamp 1676037725
transform 1 0 10120 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _698_
timestamp 1676037725
transform -1 0 11776 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _699_
timestamp 1676037725
transform 1 0 11592 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _700_
timestamp 1676037725
transform 1 0 11500 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _701_
timestamp 1676037725
transform 1 0 4048 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _702_
timestamp 1676037725
transform 1 0 6716 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _703_
timestamp 1676037725
transform 1 0 6532 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _704_
timestamp 1676037725
transform 1 0 2944 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _705_
timestamp 1676037725
transform -1 0 2852 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _706_
timestamp 1676037725
transform -1 0 6348 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _707_
timestamp 1676037725
transform -1 0 7084 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _708_
timestamp 1676037725
transform 1 0 7636 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _709_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6716 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _710_
timestamp 1676037725
transform 1 0 5244 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _711_
timestamp 1676037725
transform -1 0 6716 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _712_
timestamp 1676037725
transform -1 0 7636 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _713_
timestamp 1676037725
transform -1 0 8648 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _714_
timestamp 1676037725
transform 1 0 7360 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _715_
timestamp 1676037725
transform -1 0 9752 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _716_
timestamp 1676037725
transform -1 0 4416 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _717_
timestamp 1676037725
transform -1 0 4600 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _718_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2116 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _719_
timestamp 1676037725
transform 1 0 1656 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _720_
timestamp 1676037725
transform 1 0 1748 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _721_
timestamp 1676037725
transform -1 0 3312 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _722_
timestamp 1676037725
transform -1 0 4600 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _723_
timestamp 1676037725
transform -1 0 4324 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _724_
timestamp 1676037725
transform -1 0 5704 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _725_
timestamp 1676037725
transform 1 0 2760 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _726_
timestamp 1676037725
transform -1 0 2484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _727_
timestamp 1676037725
transform 1 0 1840 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _728_
timestamp 1676037725
transform 1 0 5152 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _729_
timestamp 1676037725
transform 1 0 6532 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _730_
timestamp 1676037725
transform -1 0 3496 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _731_
timestamp 1676037725
transform -1 0 4784 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _732_
timestamp 1676037725
transform 1 0 4692 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _733_
timestamp 1676037725
transform 1 0 12052 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o221ai_4  _734_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 9292 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__a32o_1  _735_
timestamp 1676037725
transform 1 0 11960 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _736_
timestamp 1676037725
transform 1 0 4876 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _737_
timestamp 1676037725
transform 1 0 7728 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _738_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7268 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _739_
timestamp 1676037725
transform -1 0 7176 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _740_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3036 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _741_
timestamp 1676037725
transform -1 0 6808 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _742_
timestamp 1676037725
transform -1 0 10580 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _743_
timestamp 1676037725
transform 1 0 6532 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _744_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2944 0 -1 19584
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _745_
timestamp 1676037725
transform 1 0 3036 0 -1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _746_
timestamp 1676037725
transform 1 0 9108 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _747_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _748_
timestamp 1676037725
transform -1 0 8372 0 1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _749_
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _750_
timestamp 1676037725
transform 1 0 8188 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _751_
timestamp 1676037725
transform 1 0 8188 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _752_
timestamp 1676037725
transform 1 0 7176 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _753_
timestamp 1676037725
transform -1 0 6072 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _754_
timestamp 1676037725
transform 1 0 2944 0 -1 17408
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _755_
timestamp 1676037725
transform 1 0 8464 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _756_
timestamp 1676037725
transform 1 0 8372 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _757_
timestamp 1676037725
transform 1 0 9108 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _758_
timestamp 1676037725
transform 1 0 9108 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _759_
timestamp 1676037725
transform 1 0 4508 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _760_
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _761_
timestamp 1676037725
transform 1 0 6716 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _762_
timestamp 1676037725
transform 1 0 6532 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _763_
timestamp 1676037725
transform -1 0 5428 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _764_
timestamp 1676037725
transform -1 0 4324 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _765_
timestamp 1676037725
transform 1 0 1932 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _766_
timestamp 1676037725
transform 1 0 2024 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _767_
timestamp 1676037725
transform -1 0 3496 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _768_
timestamp 1676037725
transform 1 0 2024 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _769_
timestamp 1676037725
transform -1 0 4232 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _770_
timestamp 1676037725
transform -1 0 3496 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  _798_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4048 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6348 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1676037725
transform -1 0 4416 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1676037725
transform -1 0 4416 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1676037725
transform 1 0 7820 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1676037725
transform 1 0 7820 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14260 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout14
timestamp 1676037725
transform 1 0 15640 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout16
timestamp 1676037725
transform 1 0 20976 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout18
timestamp 1676037725
transform -1 0 22448 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout19
timestamp 1676037725
transform -1 0 21436 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout20
timestamp 1676037725
transform 1 0 20424 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout21
timestamp 1676037725
transform -1 0 20332 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout22
timestamp 1676037725
transform 1 0 21988 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout23
timestamp 1676037725
transform -1 0 18584 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout24
timestamp 1676037725
transform 1 0 22724 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout25
timestamp 1676037725
transform 1 0 22724 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout26
timestamp 1676037725
transform -1 0 15088 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout27
timestamp 1676037725
transform 1 0 13248 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16468 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout29
timestamp 1676037725
transform -1 0 9660 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout30
timestamp 1676037725
transform 1 0 3220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout31
timestamp 1676037725
transform -1 0 3956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4140 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout33
timestamp 1676037725
transform -1 0 3312 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout34
timestamp 1676037725
transform 1 0 5520 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout35
timestamp 1676037725
transform 1 0 5244 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 1676037725
transform -1 0 2484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout37
timestamp 1676037725
transform -1 0 4876 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout38
timestamp 1676037725
transform 1 0 5520 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout39
timestamp 1676037725
transform 1 0 3956 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout40
timestamp 1676037725
transform -1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout41
timestamp 1676037725
transform -1 0 3496 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout42
timestamp 1676037725
transform -1 0 4600 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout43
timestamp 1676037725
transform -1 0 2392 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout44
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  fanout45
timestamp 1676037725
transform 1 0 9108 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout46
timestamp 1676037725
transform -1 0 5796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1676037725
transform 1 0 12880 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1676037725
transform 1 0 17480 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1676037725
transform -1 0 22816 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1676037725
transform 1 0 7544 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output5
timestamp 1676037725
transform 1 0 6532 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output6
timestamp 1676037725
transform -1 0 2484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output7
timestamp 1676037725
transform -1 0 3404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output8
timestamp 1676037725
transform -1 0 2576 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output9
timestamp 1676037725
transform -1 0 4508 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output10
timestamp 1676037725
transform -1 0 3496 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output11
timestamp 1676037725
transform -1 0 5980 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output12
timestamp 1676037725
transform -1 0 7084 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_47 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_48
timestamp 1676037725
transform -1 0 11224 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_49
timestamp 1676037725
transform -1 0 10580 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_50
timestamp 1676037725
transform -1 0 9936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_51
timestamp 1676037725
transform -1 0 9568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_52
timestamp 1676037725
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_53
timestamp 1676037725
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_54
timestamp 1676037725
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_55
timestamp 1676037725
transform 1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_56
timestamp 1676037725
transform -1 0 12788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_57
timestamp 1676037725
transform -1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_58
timestamp 1676037725
transform -1 0 14536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_59
timestamp 1676037725
transform -1 0 15180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_60
timestamp 1676037725
transform -1 0 15824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_61
timestamp 1676037725
transform -1 0 16468 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_62
timestamp 1676037725
transform -1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_63
timestamp 1676037725
transform -1 0 18768 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_64
timestamp 1676037725
transform -1 0 19688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_65
timestamp 1676037725
transform -1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_66
timestamp 1676037725
transform -1 0 20976 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_67
timestamp 1676037725
transform -1 0 21528 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_68
timestamp 1676037725
transform -1 0 22264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_69
timestamp 1676037725
transform -1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_70
timestamp 1676037725
transform -1 0 22264 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_71
timestamp 1676037725
transform -1 0 22908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_72
timestamp 1676037725
transform -1 0 23092 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt2_tholin_namebadge_73
timestamp 1676037725
transform 1 0 22172 0 1 3264
box -38 -48 314 592
<< labels >>
flabel metal2 s 2502 24200 2558 25000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 12438 24200 12494 25000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 17406 24200 17462 25000 0 FreeSans 224 90 0 0 io_in[1]
port 2 nsew signal input
flabel metal2 s 22374 24200 22430 25000 0 FreeSans 224 90 0 0 io_in[2]
port 3 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 4 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 io_oeb[10]
port 5 nsew signal tristate
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 io_oeb[11]
port 6 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 io_oeb[12]
port 7 nsew signal tristate
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 io_oeb[13]
port 8 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 io_oeb[14]
port 9 nsew signal tristate
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 io_oeb[15]
port 10 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 io_oeb[16]
port 11 nsew signal tristate
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 io_oeb[17]
port 12 nsew signal tristate
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 io_oeb[18]
port 13 nsew signal tristate
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 io_oeb[19]
port 14 nsew signal tristate
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 io_oeb[1]
port 15 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 io_oeb[20]
port 16 nsew signal tristate
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 io_oeb[21]
port 17 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 io_oeb[22]
port 18 nsew signal tristate
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 io_oeb[23]
port 19 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 io_oeb[24]
port 20 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 io_oeb[25]
port 21 nsew signal tristate
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 io_oeb[26]
port 22 nsew signal tristate
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 io_oeb[2]
port 23 nsew signal tristate
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 io_oeb[3]
port 24 nsew signal tristate
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 io_oeb[4]
port 25 nsew signal tristate
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 io_oeb[5]
port 26 nsew signal tristate
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 27 nsew signal tristate
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 io_oeb[7]
port 28 nsew signal tristate
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 io_oeb[8]
port 29 nsew signal tristate
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 io_oeb[9]
port 30 nsew signal tristate
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 io_out[0]
port 31 nsew signal tristate
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 io_out[1]
port 32 nsew signal tristate
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 io_out[2]
port 33 nsew signal tristate
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 io_out[3]
port 34 nsew signal tristate
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 io_out[4]
port 35 nsew signal tristate
flabel metal2 s 4710 0 4766 800 0 FreeSans 224 90 0 0 io_out[5]
port 36 nsew signal tristate
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 io_out[6]
port 37 nsew signal tristate
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 io_out[7]
port 38 nsew signal tristate
flabel metal2 s 7470 24200 7526 25000 0 FreeSans 224 90 0 0 rst
port 39 nsew signal input
flabel metal4 s 3784 2128 4104 22352 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 9465 2128 9785 22352 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 15146 2128 15466 22352 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 20827 2128 21147 22352 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 6624 2128 6944 22352 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 12305 2128 12625 22352 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 17986 2128 18306 22352 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 23667 2128 23987 22352 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 25000 25000
<< end >>
