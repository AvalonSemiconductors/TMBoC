* NGSPICE file created from wrapped_MC14500.ext - technology: sky130B

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

.subckt wrapped_MC14500 clk io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_oeb io_out[0]
+ io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8]
+ rst vccd1 vssd1
XFILLER_23_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_062_ mc14500.instr\[0\] io_out[3] vssd1 vssd1 vccd1 vccd1 _027_ sky130_fd_sc_hd__and2b_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_045_ _013_ mc14500.instr\[2\] vssd1 vssd1 vccd1 vccd1 _014_ sky130_fd_sc_hd__or2_1
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_061_ io_out[3] mc14500.instr\[1\] vssd1 vssd1 vccd1 vccd1 _026_ sky130_fd_sc_hd__and2b_1
X_044_ mc14500.instr\[3\] vssd1 vssd1 vccd1 vccd1 _013_ sky130_fd_sc_hd__inv_2
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_060_ mc14500.instr\[0\] mc14500.instr\[1\] vssd1 vssd1 vccd1 vccd1 _025_ sky130_fd_sc_hd__and2b_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_091__4 clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__inv_2
X_043_ mc14500.instr\[1\] vssd1 vssd1 vccd1 vccd1 _012_ sky130_fd_sc_hd__inv_2
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_099_ net11 _011_ vssd1 vssd1 vccd1 vccd1 mc14500.IEN_l sky130_fd_sc_hd__dfxtp_1
XFILLER_1_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapped_MC14500_7 vssd1 vssd1 vccd1 vccd1 wrapped_MC14500_7/HI io_out[8] sky130_fd_sc_hd__conb_1
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input6_A rst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_098_ net10 _000_ vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__dfxtp_4
XFILLER_1_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_16_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_097_ clknet_1_1__leaf_clk _004_ vssd1 vssd1 vccd1 vccd1 mc14500.instr\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_096_ clknet_1_1__leaf_clk _003_ vssd1 vssd1 vccd1 vccd1 mc14500.instr\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_079_ _037_ vssd1 vssd1 vccd1 vccd1 _003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input4_A io_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_095_ clknet_1_0__leaf_clk _002_ vssd1 vssd1 vccd1 vccd1 mc14500.instr\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_078_ _021_ net3 vssd1 vssd1 vccd1 vccd1 _037_ sky130_fd_sc_hd__and2_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_094_ clknet_1_0__leaf_clk _001_ vssd1 vssd1 vccd1 vccd1 mc14500.instr\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_077_ _036_ vssd1 vssd1 vccd1 vccd1 _002_ sky130_fd_sc_hd__clkbuf_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_093_ net8 _010_ vssd1 vssd1 vccd1 vccd1 mc14500.OEN_l sky130_fd_sc_hd__dfxtp_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput1 io_in[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_1
X_076_ _021_ net2 vssd1 vssd1 vccd1 vccd1 _036_ sky130_fd_sc_hd__and2_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_059_ _024_ vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__buf_2
XFILLER_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input2_A io_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput2 io_in[1] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XTAP_80 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_075_ _035_ vssd1 vssd1 vccd1 vccd1 _001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_058_ _013_ _021_ _023_ vssd1 vssd1 vccd1 vccd1 _024_ sky130_fd_sc_hd__and3_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput3 io_in[2] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XTAP_70 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_074_ _021_ net1 vssd1 vssd1 vccd1 vccd1 _035_ sky130_fd_sc_hd__and2_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_057_ mc14500.instr\[2\] _022_ vssd1 vssd1 vccd1 vccd1 _023_ sky130_fd_sc_hd__nor2_1
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_60 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_092__5 clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__inv_2
Xinput4 io_in[3] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XTAP_82 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_073_ net9 io_oeb vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__nor2_2
XFILLER_24_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_056_ mc14500.instr\[0\] mc14500.instr\[1\] vssd1 vssd1 vccd1 vccd1 _022_ sky130_fd_sc_hd__or2_2
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput5 io_in[4] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_83 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_50 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_72 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_055_ mc14500.skip vssd1 vssd1 vccd1 vccd1 _021_ sky130_fd_sc_hd__inv_2
XFILLER_23_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput6 rst vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XTAP_84 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_51 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_73 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_071_ mc14500.instr\[3\] mc14500.instr\[2\] _034_ _025_ net6 vssd1 vssd1 vccd1 vccd1
+ _005_ sky130_fd_sc_hd__a41o_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_054_ _020_ vssd1 vssd1 vccd1 vccd1 io_oeb sky130_fd_sc_hd__clkbuf_4
XFILLER_7_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_85 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_070_ io_out[3] vssd1 vssd1 vccd1 vccd1 _034_ sky130_fd_sc_hd__inv_2
XFILLER_19_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_053_ mc14500.instr\[1\] _014_ mc14500.OEN_l vssd1 vssd1 vccd1 vccd1 _020_ sky130_fd_sc_hd__or3b_1
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_86 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_052_ _019_ vssd1 vssd1 vccd1 vccd1 _010_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_8_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_87 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_76 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_051_ mc14500.OEN_l net5 _018_ vssd1 vssd1 vccd1 vccd1 _019_ sky130_fd_sc_hd__mux2_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_88 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_050_ _014_ _017_ vssd1 vssd1 vccd1 vccd1 _018_ sky130_fd_sc_hd__nor2_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_102_ clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__buf_2
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_89 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_57 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_100_ net12 _005_ vssd1 vssd1 vccd1 vccd1 mc14500.skip sky130_fd_sc_hd__dfxtp_1
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_58 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_090__3 clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__inv_2
XFILLER_12_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_59 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_089_ _042_ vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__buf_2
XFILLER_17_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_input5_A io_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_088_ mc14500.instr\[0\] _012_ mc14500.instr\[3\] mc14500.instr\[2\] vssd1 vssd1
+ vccd1 vccd1 _042_ sky130_fd_sc_hd__and4b_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_087_ _041_ vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__buf_2
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_086_ mc14500.instr\[3\] mc14500.instr\[2\] mc14500.instr\[0\] _012_ vssd1 vssd1
+ vccd1 vccd1 _041_ sky130_fd_sc_hd__and4_1
XFILLER_8_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_069_ _031_ _033_ net6 vssd1 vssd1 vccd1 vccd1 _000_ sky130_fd_sc_hd__o21ba_1
XFILLER_10_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input3_A io_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_085_ _040_ vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__buf_2
X_068_ mc14500.instr\[3\] _023_ _032_ io_out[3] vssd1 vssd1 vccd1 vccd1 _033_ sky130_fd_sc_hd__o31a_1
XFILLER_0_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_084_ mc14500.instr\[3\] mc14500.instr\[2\] mc14500.instr\[0\] mc14500.instr\[1\]
+ vssd1 vssd1 vccd1 vccd1 _040_ sky130_fd_sc_hd__and4_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_067_ mc14500.instr\[2\] _017_ _022_ vssd1 vssd1 vccd1 vccd1 _032_ sky130_fd_sc_hd__and3_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_083_ io_out[3] _022_ _039_ vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__a21oi_4
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_066_ mc14500.instr\[2\] _022_ _029_ _030_ _013_ vssd1 vssd1 vccd1 vccd1 _031_ sky130_fd_sc_hd__o221a_1
X_049_ mc14500.instr\[0\] mc14500.instr\[1\] vssd1 vssd1 vccd1 vccd1 _017_ sky130_fd_sc_hd__nand2_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input1_A io_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_082_ io_out[3] _022_ mc14500.OEN_l vssd1 vssd1 vccd1 vccd1 _039_ sky130_fd_sc_hd__o21ai_1
XFILLER_17_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_065_ _026_ mc14500.instr\[0\] net5 mc14500.IEN_l vssd1 vssd1 vccd1 vccd1 _030_ sky130_fd_sc_hd__and4b_1
XFILLER_9_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_048_ _016_ vssd1 vssd1 vccd1 vccd1 _011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_072__1 clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__inv_2
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_081_ _038_ vssd1 vssd1 vccd1 vccd1 _004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_064_ mc14500.instr\[2\] _025_ _026_ _027_ _028_ vssd1 vssd1 vccd1 vccd1 _029_ sky130_fd_sc_hd__o221a_1
XFILLER_9_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_047_ net5 mc14500.IEN_l _015_ vssd1 vssd1 vccd1 vccd1 _016_ sky130_fd_sc_hd__mux2_1
X_072__2 clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__inv_2
XFILLER_6_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_080_ _021_ net4 vssd1 vssd1 vccd1 vccd1 _038_ sky130_fd_sc_hd__and2_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_063_ mc14500.IEN_l net5 vssd1 vssd1 vccd1 vccd1 _028_ sky130_fd_sc_hd__nand2_1
XFILLER_9_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_046_ mc14500.instr\[0\] _012_ _014_ vssd1 vssd1 vccd1 vccd1 _015_ sky130_fd_sc_hd__or3_1
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
.ends

