magic
tech sky130B
magscale 1 2
timestamp 1680008150
<< nwell >>
rect 1066 66629 68854 67195
rect 1066 65541 68854 66107
rect 1066 64453 68854 65019
rect 1066 63365 68854 63931
rect 1066 62277 68854 62843
rect 1066 61189 68854 61755
rect 1066 60101 68854 60667
rect 1066 59013 68854 59579
rect 1066 57925 68854 58491
rect 1066 56837 68854 57403
rect 1066 55749 68854 56315
rect 1066 54661 68854 55227
rect 1066 53573 68854 54139
rect 1066 52485 68854 53051
rect 1066 51397 68854 51963
rect 1066 50309 68854 50875
rect 1066 49221 68854 49787
rect 1066 48133 68854 48699
rect 1066 47045 68854 47611
rect 1066 45957 68854 46523
rect 1066 44869 68854 45435
rect 1066 43781 68854 44347
rect 1066 42693 68854 43259
rect 1066 41605 68854 42171
rect 1066 40517 68854 41083
rect 1066 39429 68854 39995
rect 1066 38341 68854 38907
rect 1066 37253 68854 37819
rect 1066 36165 68854 36731
rect 1066 35077 68854 35643
rect 1066 33989 68854 34555
rect 1066 32901 68854 33467
rect 1066 31813 68854 32379
rect 1066 30725 68854 31291
rect 1066 29637 68854 30203
rect 1066 28549 68854 29115
rect 1066 27461 68854 28027
rect 1066 26373 68854 26939
rect 1066 25285 68854 25851
rect 1066 24197 68854 24763
rect 1066 23109 68854 23675
rect 1066 22021 68854 22587
rect 1066 20933 68854 21499
rect 1066 19845 68854 20411
rect 1066 18757 68854 19323
rect 1066 17669 68854 18235
rect 1066 16581 68854 17147
rect 1066 15493 68854 16059
rect 1066 14405 68854 14971
rect 1066 13317 68854 13883
rect 1066 12229 68854 12795
rect 1066 11141 68854 11707
rect 1066 10053 68854 10619
rect 1066 8965 68854 9531
rect 1066 7877 68854 8443
rect 1066 6789 68854 7355
rect 1066 5701 68854 6267
rect 1066 4613 68854 5179
rect 1066 3525 68854 4091
rect 1066 2437 68854 3003
<< obsli1 >>
rect 1104 2159 68816 67473
<< obsm1 >>
rect 1104 2128 69078 69148
<< metal2 >>
rect 2778 69200 2834 70000
rect 7378 69200 7434 70000
rect 11978 69200 12034 70000
rect 16578 69200 16634 70000
rect 21178 69200 21234 70000
rect 25778 69200 25834 70000
rect 30378 69200 30434 70000
rect 34978 69200 35034 70000
rect 39578 69200 39634 70000
rect 44178 69200 44234 70000
rect 48778 69200 48834 70000
rect 53378 69200 53434 70000
rect 57978 69200 58034 70000
rect 62578 69200 62634 70000
rect 67178 69200 67234 70000
<< obsm2 >>
rect 2890 69144 7322 69306
rect 7490 69144 11922 69306
rect 12090 69144 16522 69306
rect 16690 69144 21122 69306
rect 21290 69144 25722 69306
rect 25890 69144 30322 69306
rect 30490 69144 34922 69306
rect 35090 69144 39522 69306
rect 39690 69144 44122 69306
rect 44290 69144 48722 69306
rect 48890 69144 53322 69306
rect 53490 69144 57922 69306
rect 58090 69144 62522 69306
rect 62690 69144 67122 69306
rect 67290 69144 69074 69306
rect 2834 1799 69074 69144
<< metal3 >>
rect 69200 67872 70000 67992
rect 69200 65424 70000 65544
rect 69200 62976 70000 63096
rect 69200 60528 70000 60648
rect 69200 58080 70000 58200
rect 69200 55632 70000 55752
rect 69200 53184 70000 53304
rect 69200 50736 70000 50856
rect 69200 48288 70000 48408
rect 69200 45840 70000 45960
rect 69200 43392 70000 43512
rect 69200 40944 70000 41064
rect 69200 38496 70000 38616
rect 69200 36048 70000 36168
rect 69200 33600 70000 33720
rect 69200 31152 70000 31272
rect 69200 28704 70000 28824
rect 69200 26256 70000 26376
rect 69200 23808 70000 23928
rect 69200 21360 70000 21480
rect 69200 18912 70000 19032
rect 69200 16464 70000 16584
rect 69200 14016 70000 14136
rect 69200 11568 70000 11688
rect 69200 9120 70000 9240
rect 69200 6672 70000 6792
rect 69200 4224 70000 4344
rect 69200 1776 70000 1896
<< obsm3 >>
rect 4210 67792 69120 67965
rect 4210 65624 69200 67792
rect 4210 65344 69120 65624
rect 4210 63176 69200 65344
rect 4210 62896 69120 63176
rect 4210 60728 69200 62896
rect 4210 60448 69120 60728
rect 4210 58280 69200 60448
rect 4210 58000 69120 58280
rect 4210 55832 69200 58000
rect 4210 55552 69120 55832
rect 4210 53384 69200 55552
rect 4210 53104 69120 53384
rect 4210 50936 69200 53104
rect 4210 50656 69120 50936
rect 4210 48488 69200 50656
rect 4210 48208 69120 48488
rect 4210 46040 69200 48208
rect 4210 45760 69120 46040
rect 4210 43592 69200 45760
rect 4210 43312 69120 43592
rect 4210 41144 69200 43312
rect 4210 40864 69120 41144
rect 4210 38696 69200 40864
rect 4210 38416 69120 38696
rect 4210 36248 69200 38416
rect 4210 35968 69120 36248
rect 4210 33800 69200 35968
rect 4210 33520 69120 33800
rect 4210 31352 69200 33520
rect 4210 31072 69120 31352
rect 4210 28904 69200 31072
rect 4210 28624 69120 28904
rect 4210 26456 69200 28624
rect 4210 26176 69120 26456
rect 4210 24008 69200 26176
rect 4210 23728 69120 24008
rect 4210 21560 69200 23728
rect 4210 21280 69120 21560
rect 4210 19112 69200 21280
rect 4210 18832 69120 19112
rect 4210 16664 69200 18832
rect 4210 16384 69120 16664
rect 4210 14216 69200 16384
rect 4210 13936 69120 14216
rect 4210 11768 69200 13936
rect 4210 11488 69120 11768
rect 4210 9320 69200 11488
rect 4210 9040 69120 9320
rect 4210 6872 69200 9040
rect 4210 6592 69120 6872
rect 4210 4424 69200 6592
rect 4210 4144 69120 4424
rect 4210 1976 69200 4144
rect 4210 1803 69120 1976
<< metal4 >>
rect 4208 2128 4528 67504
rect 19568 2128 19888 67504
rect 34928 2128 35248 67504
rect 50288 2128 50608 67504
rect 65648 2128 65968 67504
<< obsm4 >>
rect 18459 9555 19488 64973
rect 19968 9555 34848 64973
rect 35328 9555 50208 64973
rect 50688 9555 59557 64973
<< labels >>
rlabel metal2 s 62578 69200 62634 70000 6 clk
port 1 nsew signal input
rlabel metal2 s 2778 69200 2834 70000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 48778 69200 48834 70000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 53378 69200 53434 70000 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 57978 69200 58034 70000 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 7378 69200 7434 70000 6 io_in[1]
port 6 nsew signal input
rlabel metal2 s 11978 69200 12034 70000 6 io_in[2]
port 7 nsew signal input
rlabel metal2 s 16578 69200 16634 70000 6 io_in[3]
port 8 nsew signal input
rlabel metal2 s 21178 69200 21234 70000 6 io_in[4]
port 9 nsew signal input
rlabel metal2 s 25778 69200 25834 70000 6 io_in[5]
port 10 nsew signal input
rlabel metal2 s 30378 69200 30434 70000 6 io_in[6]
port 11 nsew signal input
rlabel metal2 s 34978 69200 35034 70000 6 io_in[7]
port 12 nsew signal input
rlabel metal2 s 39578 69200 39634 70000 6 io_in[8]
port 13 nsew signal input
rlabel metal2 s 44178 69200 44234 70000 6 io_in[9]
port 14 nsew signal input
rlabel metal3 s 69200 67872 70000 67992 6 io_oeb
port 15 nsew signal output
rlabel metal3 s 69200 1776 70000 1896 6 io_out[0]
port 16 nsew signal output
rlabel metal3 s 69200 26256 70000 26376 6 io_out[10]
port 17 nsew signal output
rlabel metal3 s 69200 28704 70000 28824 6 io_out[11]
port 18 nsew signal output
rlabel metal3 s 69200 31152 70000 31272 6 io_out[12]
port 19 nsew signal output
rlabel metal3 s 69200 33600 70000 33720 6 io_out[13]
port 20 nsew signal output
rlabel metal3 s 69200 36048 70000 36168 6 io_out[14]
port 21 nsew signal output
rlabel metal3 s 69200 38496 70000 38616 6 io_out[15]
port 22 nsew signal output
rlabel metal3 s 69200 40944 70000 41064 6 io_out[16]
port 23 nsew signal output
rlabel metal3 s 69200 43392 70000 43512 6 io_out[17]
port 24 nsew signal output
rlabel metal3 s 69200 45840 70000 45960 6 io_out[18]
port 25 nsew signal output
rlabel metal3 s 69200 48288 70000 48408 6 io_out[19]
port 26 nsew signal output
rlabel metal3 s 69200 4224 70000 4344 6 io_out[1]
port 27 nsew signal output
rlabel metal3 s 69200 50736 70000 50856 6 io_out[20]
port 28 nsew signal output
rlabel metal3 s 69200 53184 70000 53304 6 io_out[21]
port 29 nsew signal output
rlabel metal3 s 69200 55632 70000 55752 6 io_out[22]
port 30 nsew signal output
rlabel metal3 s 69200 58080 70000 58200 6 io_out[23]
port 31 nsew signal output
rlabel metal3 s 69200 60528 70000 60648 6 io_out[24]
port 32 nsew signal output
rlabel metal3 s 69200 62976 70000 63096 6 io_out[25]
port 33 nsew signal output
rlabel metal3 s 69200 65424 70000 65544 6 io_out[26]
port 34 nsew signal output
rlabel metal3 s 69200 6672 70000 6792 6 io_out[2]
port 35 nsew signal output
rlabel metal3 s 69200 9120 70000 9240 6 io_out[3]
port 36 nsew signal output
rlabel metal3 s 69200 11568 70000 11688 6 io_out[4]
port 37 nsew signal output
rlabel metal3 s 69200 14016 70000 14136 6 io_out[5]
port 38 nsew signal output
rlabel metal3 s 69200 16464 70000 16584 6 io_out[6]
port 39 nsew signal output
rlabel metal3 s 69200 18912 70000 19032 6 io_out[7]
port 40 nsew signal output
rlabel metal3 s 69200 21360 70000 21480 6 io_out[8]
port 41 nsew signal output
rlabel metal3 s 69200 23808 70000 23928 6 io_out[9]
port 42 nsew signal output
rlabel metal2 s 67178 69200 67234 70000 6 rst
port 43 nsew signal input
rlabel metal4 s 4208 2128 4528 67504 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 67504 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 67504 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 67504 6 vssd1
port 45 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 67504 6 vssd1
port 45 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 70000 70000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9688640
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/AS1802/runs/23_03_28_14_51/results/signoff/wrapped_as1802.magic.gds
string GDS_START 1222116
<< end >>

