magic
tech sky130B
magscale 1 2
timestamp 1680007868
<< viali >>
rect 1777 19805 1811 19839
rect 2053 19805 2087 19839
rect 8861 18241 8895 18275
rect 9045 18241 9079 18275
rect 8953 18037 8987 18071
rect 5365 17697 5399 17731
rect 8033 17697 8067 17731
rect 10701 17697 10735 17731
rect 7021 17629 7055 17663
rect 7113 17629 7147 17663
rect 7205 17629 7239 17663
rect 8217 17629 8251 17663
rect 8309 17629 8343 17663
rect 9321 17629 9355 17663
rect 9505 17629 9539 17663
rect 10425 17629 10459 17663
rect 10517 17629 10551 17663
rect 5181 17561 5215 17595
rect 8033 17561 8067 17595
rect 4721 17493 4755 17527
rect 5089 17493 5123 17527
rect 6837 17493 6871 17527
rect 9413 17493 9447 17527
rect 10701 17493 10735 17527
rect 5273 17289 5307 17323
rect 6929 17289 6963 17323
rect 9413 17289 9447 17323
rect 7297 17221 7331 17255
rect 7941 17221 7975 17255
rect 3065 17153 3099 17187
rect 5181 17153 5215 17187
rect 7113 17153 7147 17187
rect 7205 17153 7239 17187
rect 7481 17153 7515 17187
rect 8125 17153 8159 17187
rect 8309 17153 8343 17187
rect 9597 17153 9631 17187
rect 9689 17153 9723 17187
rect 9873 17153 9907 17187
rect 9965 17153 9999 17187
rect 10609 17153 10643 17187
rect 3157 17085 3191 17119
rect 3249 17085 3283 17119
rect 5365 17085 5399 17119
rect 10425 17085 10459 17119
rect 10793 17085 10827 17119
rect 2697 16949 2731 16983
rect 4813 16949 4847 16983
rect 9321 16745 9355 16779
rect 10609 16745 10643 16779
rect 6837 16677 6871 16711
rect 3065 16609 3099 16643
rect 3249 16609 3283 16643
rect 5733 16609 5767 16643
rect 7941 16609 7975 16643
rect 9137 16609 9171 16643
rect 4997 16541 5031 16575
rect 5273 16541 5307 16575
rect 5641 16541 5675 16575
rect 6377 16541 6411 16575
rect 7021 16541 7055 16575
rect 7323 16541 7357 16575
rect 7481 16541 7515 16575
rect 8125 16541 8159 16575
rect 9413 16541 9447 16575
rect 10609 16541 10643 16575
rect 10885 16541 10919 16575
rect 7113 16473 7147 16507
rect 7205 16473 7239 16507
rect 8309 16473 8343 16507
rect 10701 16473 10735 16507
rect 2605 16405 2639 16439
rect 2973 16405 3007 16439
rect 9137 16405 9171 16439
rect 2605 16201 2639 16235
rect 4905 16201 4939 16235
rect 10057 16133 10091 16167
rect 10609 16133 10643 16167
rect 11805 16133 11839 16167
rect 2513 16065 2547 16099
rect 4813 16065 4847 16099
rect 8309 16065 8343 16099
rect 11713 16065 11747 16099
rect 11897 16065 11931 16099
rect 2697 15997 2731 16031
rect 5089 15997 5123 16031
rect 8401 15997 8435 16031
rect 8493 15997 8527 16031
rect 8585 15997 8619 16031
rect 9873 15997 9907 16031
rect 10149 15997 10183 16031
rect 10609 15929 10643 15963
rect 2145 15861 2179 15895
rect 4445 15861 4479 15895
rect 8125 15861 8159 15895
rect 10425 15657 10459 15691
rect 10977 15589 11011 15623
rect 4813 15521 4847 15555
rect 4997 15521 5031 15555
rect 7021 15453 7055 15487
rect 7205 15453 7239 15487
rect 9321 15453 9355 15487
rect 10333 15453 10367 15487
rect 10517 15453 10551 15487
rect 11345 15453 11379 15487
rect 11161 15385 11195 15419
rect 4353 15317 4387 15351
rect 4721 15317 4755 15351
rect 7021 15317 7055 15351
rect 9229 15317 9263 15351
rect 8033 15113 8067 15147
rect 8677 15113 8711 15147
rect 2053 15045 2087 15079
rect 4721 15045 4755 15079
rect 7021 15045 7055 15079
rect 9965 15045 9999 15079
rect 10977 15045 11011 15079
rect 1869 14977 1903 15011
rect 2145 14977 2179 15011
rect 2973 14977 3007 15011
rect 3157 14977 3191 15011
rect 4537 14977 4571 15011
rect 4813 14977 4847 15011
rect 4905 14977 4939 15011
rect 6929 14977 6963 15011
rect 8125 14977 8159 15011
rect 8953 14977 8987 15011
rect 10149 14977 10183 15011
rect 10425 14977 10459 15011
rect 10885 14977 10919 15011
rect 11069 14977 11103 15011
rect 7113 14909 7147 14943
rect 8861 14909 8895 14943
rect 9321 14909 9355 14943
rect 10057 14909 10091 14943
rect 10333 14909 10367 14943
rect 1869 14773 1903 14807
rect 3065 14773 3099 14807
rect 5089 14773 5123 14807
rect 6561 14773 6595 14807
rect 1777 14569 1811 14603
rect 3985 14569 4019 14603
rect 5089 14569 5123 14603
rect 9505 14569 9539 14603
rect 3341 14501 3375 14535
rect 4353 14433 4387 14467
rect 6561 14433 6595 14467
rect 6653 14433 6687 14467
rect 9413 14433 9447 14467
rect 9597 14433 9631 14467
rect 1961 14365 1995 14399
rect 2145 14365 2179 14399
rect 4169 14365 4203 14399
rect 4445 14365 4479 14399
rect 4997 14365 5031 14399
rect 5181 14365 5215 14399
rect 5549 14365 5583 14399
rect 9321 14365 9355 14399
rect 11345 14365 11379 14399
rect 2973 14297 3007 14331
rect 3157 14297 3191 14331
rect 6745 14297 6779 14331
rect 10793 14297 10827 14331
rect 5365 14229 5399 14263
rect 7113 14229 7147 14263
rect 2329 14025 2363 14059
rect 3610 14025 3644 14059
rect 5273 14025 5307 14059
rect 7205 14025 7239 14059
rect 3709 13957 3743 13991
rect 6837 13957 6871 13991
rect 6929 13957 6963 13991
rect 9229 13957 9263 13991
rect 9597 13957 9631 13991
rect 2053 13889 2087 13923
rect 2145 13889 2179 13923
rect 3433 13889 3467 13923
rect 3525 13889 3559 13923
rect 4629 13889 4663 13923
rect 6561 13889 6595 13923
rect 6653 13889 6687 13923
rect 7021 13889 7055 13923
rect 8309 13889 8343 13923
rect 8585 13889 8619 13923
rect 8769 13889 8803 13923
rect 9413 13889 9447 13923
rect 9689 13889 9723 13923
rect 10793 13889 10827 13923
rect 13093 13889 13127 13923
rect 13277 13889 13311 13923
rect 15301 13889 15335 13923
rect 2329 13821 2363 13855
rect 4813 13821 4847 13855
rect 4905 13821 4939 13855
rect 8125 13821 8159 13855
rect 13645 13821 13679 13855
rect 15209 13821 15243 13855
rect 15669 13753 15703 13787
rect 10609 13685 10643 13719
rect 13277 13481 13311 13515
rect 14381 13481 14415 13515
rect 17693 13481 17727 13515
rect 19533 13481 19567 13515
rect 17877 13413 17911 13447
rect 18613 13413 18647 13447
rect 2513 13345 2547 13379
rect 12081 13345 12115 13379
rect 12817 13345 12851 13379
rect 15577 13345 15611 13379
rect 2237 13277 2271 13311
rect 3157 13277 3191 13311
rect 3249 13277 3283 13311
rect 9137 13277 9171 13311
rect 9321 13277 9355 13311
rect 10517 13277 10551 13311
rect 10701 13277 10735 13311
rect 10793 13277 10827 13311
rect 10885 13277 10919 13311
rect 11621 13277 11655 13311
rect 11805 13277 11839 13311
rect 12173 13277 12207 13311
rect 13461 13277 13495 13311
rect 13553 13277 13587 13311
rect 14381 13277 14415 13311
rect 15485 13277 15519 13311
rect 16037 13277 16071 13311
rect 16497 13277 16531 13311
rect 16590 13277 16624 13311
rect 17417 13277 17451 13311
rect 17785 13277 17819 13311
rect 18797 13277 18831 13311
rect 18889 13277 18923 13311
rect 19533 13277 19567 13311
rect 3433 13209 3467 13243
rect 13277 13209 13311 13243
rect 18613 13209 18647 13243
rect 3157 13141 3191 13175
rect 9229 13141 9263 13175
rect 11161 13141 11195 13175
rect 15853 13141 15887 13175
rect 16865 13141 16899 13175
rect 17509 13141 17543 13175
rect 18153 13141 18187 13175
rect 3617 12937 3651 12971
rect 9137 12937 9171 12971
rect 11805 12937 11839 12971
rect 12449 12937 12483 12971
rect 13553 12937 13587 12971
rect 15669 12937 15703 12971
rect 20085 12937 20119 12971
rect 20269 12937 20303 12971
rect 3249 12869 3283 12903
rect 3449 12869 3483 12903
rect 5733 12869 5767 12903
rect 9289 12869 9323 12903
rect 9505 12869 9539 12903
rect 16865 12869 16899 12903
rect 2697 12801 2731 12835
rect 4629 12801 4663 12835
rect 4813 12801 4847 12835
rect 5549 12801 5583 12835
rect 5825 12801 5859 12835
rect 6561 12801 6595 12835
rect 6837 12801 6871 12835
rect 7481 12801 7515 12835
rect 8401 12801 8435 12835
rect 10333 12801 10367 12835
rect 10517 12801 10551 12835
rect 10885 12801 10919 12835
rect 10977 12801 11011 12835
rect 11161 12801 11195 12835
rect 11713 12801 11747 12835
rect 12357 12801 12391 12835
rect 13461 12801 13495 12835
rect 13645 12801 13679 12835
rect 15485 12801 15519 12835
rect 17049 12801 17083 12835
rect 18153 12801 18187 12835
rect 18245 12801 18279 12835
rect 18337 12801 18371 12835
rect 18521 12801 18555 12835
rect 19349 12801 19383 12835
rect 19441 12801 19475 12835
rect 20210 12801 20244 12835
rect 20637 12801 20671 12835
rect 22201 12801 22235 12835
rect 2421 12733 2455 12767
rect 7297 12733 7331 12767
rect 8677 12733 8711 12767
rect 13277 12733 13311 12767
rect 15209 12733 15243 12767
rect 15301 12733 15335 12767
rect 15393 12733 15427 12767
rect 19625 12733 19659 12767
rect 20729 12733 20763 12767
rect 22109 12733 22143 12767
rect 6745 12665 6779 12699
rect 8585 12665 8619 12699
rect 3433 12597 3467 12631
rect 4629 12597 4663 12631
rect 5549 12597 5583 12631
rect 6837 12597 6871 12631
rect 7665 12597 7699 12631
rect 8217 12597 8251 12631
rect 9321 12597 9355 12631
rect 13829 12597 13863 12631
rect 17141 12597 17175 12631
rect 17877 12597 17911 12631
rect 19533 12597 19567 12631
rect 3157 12393 3191 12427
rect 7021 12393 7055 12427
rect 7757 12393 7791 12427
rect 10977 12393 11011 12427
rect 13093 12393 13127 12427
rect 5825 12325 5859 12359
rect 11437 12325 11471 12359
rect 17141 12325 17175 12359
rect 2329 12257 2363 12291
rect 3985 12257 4019 12291
rect 4721 12257 4755 12291
rect 5917 12257 5951 12291
rect 8125 12257 8159 12291
rect 10333 12257 10367 12291
rect 12081 12257 12115 12291
rect 13277 12257 13311 12291
rect 15301 12257 15335 12291
rect 20453 12257 20487 12291
rect 2145 12189 2179 12223
rect 2421 12189 2455 12223
rect 2881 12189 2915 12223
rect 5641 12189 5675 12223
rect 6745 12189 6779 12223
rect 7941 12189 7975 12223
rect 10701 12189 10735 12223
rect 10793 12189 10827 12223
rect 11805 12189 11839 12223
rect 13369 12189 13403 12223
rect 13461 12189 13495 12223
rect 13553 12189 13587 12223
rect 15025 12189 15059 12223
rect 15209 12189 15243 12223
rect 15393 12189 15427 12223
rect 15577 12189 15611 12223
rect 16405 12189 16439 12223
rect 16589 12189 16623 12223
rect 17233 12189 17267 12223
rect 17693 12189 17727 12223
rect 17877 12189 17911 12223
rect 20269 12189 20303 12223
rect 20361 12189 20395 12223
rect 20545 12189 20579 12223
rect 21557 12189 21591 12223
rect 21741 12189 21775 12223
rect 2973 12121 3007 12155
rect 3157 12121 3191 12155
rect 4353 12121 4387 12155
rect 7021 12121 7055 12155
rect 10425 12121 10459 12155
rect 21649 12121 21683 12155
rect 1961 12053 1995 12087
rect 4169 12053 4203 12087
rect 4261 12053 4295 12087
rect 5457 12053 5491 12087
rect 6837 12053 6871 12087
rect 10517 12053 10551 12087
rect 11897 12053 11931 12087
rect 15761 12053 15795 12087
rect 16497 12053 16531 12087
rect 17785 12053 17819 12087
rect 20085 12053 20119 12087
rect 2329 11781 2363 11815
rect 19993 11781 20027 11815
rect 20085 11781 20119 11815
rect 2145 11713 2179 11747
rect 2421 11713 2455 11747
rect 4445 11713 4479 11747
rect 4629 11713 4663 11747
rect 15577 11713 15611 11747
rect 17141 11713 17175 11747
rect 17234 11713 17268 11747
rect 17417 11713 17451 11747
rect 17509 11713 17543 11747
rect 17647 11713 17681 11747
rect 19717 11713 19751 11747
rect 21189 11713 21223 11747
rect 21373 11713 21407 11747
rect 4353 11645 4387 11679
rect 15393 11645 15427 11679
rect 19625 11645 19659 11679
rect 2145 11577 2179 11611
rect 4813 11509 4847 11543
rect 17785 11509 17819 11543
rect 19441 11509 19475 11543
rect 21189 11509 21223 11543
rect 6469 11305 6503 11339
rect 8309 11305 8343 11339
rect 18797 11305 18831 11339
rect 21281 11305 21315 11339
rect 1869 11237 1903 11271
rect 14749 11237 14783 11271
rect 21189 11237 21223 11271
rect 17693 11169 17727 11203
rect 17877 11169 17911 11203
rect 18153 11169 18187 11203
rect 21373 11169 21407 11203
rect 1685 11101 1719 11135
rect 5089 11101 5123 11135
rect 5356 11101 5390 11135
rect 6929 11101 6963 11135
rect 7196 11101 7230 11135
rect 13369 11101 13403 11135
rect 13461 11101 13495 11135
rect 13645 11101 13679 11135
rect 13737 11101 13771 11135
rect 14473 11101 14507 11135
rect 14565 11101 14599 11135
rect 14841 11101 14875 11135
rect 15485 11101 15519 11135
rect 15577 11101 15611 11135
rect 15761 11101 15795 11135
rect 15853 11101 15887 11135
rect 16773 11101 16807 11135
rect 17969 11101 18003 11135
rect 18061 11101 18095 11135
rect 18705 11101 18739 11135
rect 18889 11101 18923 11135
rect 19625 11101 19659 11135
rect 19717 11101 19751 11135
rect 19993 11101 20027 11135
rect 20821 11101 20855 11135
rect 21097 11101 21131 11135
rect 21557 11101 21591 11135
rect 15301 11033 15335 11067
rect 16497 11033 16531 11067
rect 19809 11033 19843 11067
rect 13185 10965 13219 10999
rect 14289 10965 14323 10999
rect 19441 10965 19475 10999
rect 3065 10761 3099 10795
rect 4537 10761 4571 10795
rect 8585 10761 8619 10795
rect 10885 10761 10919 10795
rect 13829 10761 13863 10795
rect 15577 10761 15611 10795
rect 18797 10761 18831 10795
rect 21005 10761 21039 10795
rect 1952 10693 1986 10727
rect 5650 10693 5684 10727
rect 7472 10693 7506 10727
rect 9772 10693 9806 10727
rect 13277 10693 13311 10727
rect 15209 10693 15243 10727
rect 19257 10693 19291 10727
rect 7205 10625 7239 10659
rect 11989 10625 12023 10659
rect 12173 10625 12207 10659
rect 12265 10625 12299 10659
rect 13001 10625 13035 10659
rect 14105 10625 14139 10659
rect 16221 10625 16255 10659
rect 16865 10625 16899 10659
rect 17049 10625 17083 10659
rect 17141 10625 17175 10659
rect 17233 10625 17267 10659
rect 18521 10625 18555 10659
rect 19441 10625 19475 10659
rect 19533 10625 19567 10659
rect 19717 10625 19751 10659
rect 19809 10625 19843 10659
rect 22017 10625 22051 10659
rect 22201 10625 22235 10659
rect 1685 10557 1719 10591
rect 5917 10557 5951 10591
rect 9505 10557 9539 10591
rect 12909 10557 12943 10591
rect 13369 10557 13403 10591
rect 13829 10557 13863 10591
rect 14013 10557 14047 10591
rect 15025 10557 15059 10591
rect 15117 10557 15151 10591
rect 18337 10557 18371 10591
rect 18429 10557 18463 10591
rect 18613 10557 18647 10591
rect 21465 10557 21499 10591
rect 11989 10489 12023 10523
rect 21097 10489 21131 10523
rect 12725 10421 12759 10455
rect 16129 10421 16163 10455
rect 17509 10421 17543 10455
rect 22017 10421 22051 10455
rect 3065 10217 3099 10251
rect 5549 10217 5583 10251
rect 8493 10217 8527 10251
rect 10885 10217 10919 10251
rect 13461 10217 13495 10251
rect 15669 10217 15703 10251
rect 16957 10217 16991 10251
rect 19625 10217 19659 10251
rect 19993 10217 20027 10251
rect 20637 10217 20671 10251
rect 20453 10149 20487 10183
rect 4169 10081 4203 10115
rect 7113 10081 7147 10115
rect 13553 10081 13587 10115
rect 16313 10081 16347 10115
rect 19717 10081 19751 10115
rect 1685 10013 1719 10047
rect 1941 10013 1975 10047
rect 4436 10013 4470 10047
rect 9505 10013 9539 10047
rect 9772 10013 9806 10047
rect 13090 10013 13124 10047
rect 17049 10013 17083 10047
rect 19441 10013 19475 10047
rect 7380 9945 7414 9979
rect 20821 9945 20855 9979
rect 12909 9877 12943 9911
rect 13093 9877 13127 9911
rect 16037 9877 16071 9911
rect 16129 9877 16163 9911
rect 20611 9877 20645 9911
rect 15853 9673 15887 9707
rect 16957 9673 16991 9707
rect 9864 9605 9898 9639
rect 18061 9605 18095 9639
rect 21189 9605 21223 9639
rect 1777 9537 1811 9571
rect 2044 9537 2078 9571
rect 4261 9537 4295 9571
rect 4528 9537 4562 9571
rect 9597 9537 9631 9571
rect 15761 9537 15795 9571
rect 15945 9537 15979 9571
rect 16865 9537 16899 9571
rect 17141 9537 17175 9571
rect 17785 9537 17819 9571
rect 18521 9537 18555 9571
rect 18705 9537 18739 9571
rect 18797 9537 18831 9571
rect 20821 9537 20855 9571
rect 20914 9537 20948 9571
rect 21097 9537 21131 9571
rect 21286 9537 21320 9571
rect 22017 9537 22051 9571
rect 22201 9537 22235 9571
rect 18061 9469 18095 9503
rect 3157 9401 3191 9435
rect 5641 9401 5675 9435
rect 10977 9401 11011 9435
rect 17877 9401 17911 9435
rect 18521 9401 18555 9435
rect 17141 9333 17175 9367
rect 21465 9333 21499 9367
rect 22017 9333 22051 9367
rect 3433 9129 3467 9163
rect 10885 9129 10919 9163
rect 13093 9129 13127 9163
rect 14933 9129 14967 9163
rect 17325 9061 17359 9095
rect 21005 9061 21039 9095
rect 2053 8993 2087 9027
rect 9505 8993 9539 9027
rect 14565 8993 14599 9027
rect 15669 8993 15703 9027
rect 18061 8993 18095 9027
rect 2320 8925 2354 8959
rect 9772 8925 9806 8959
rect 13001 8925 13035 8959
rect 13185 8925 13219 8959
rect 14749 8925 14783 8959
rect 15761 8925 15795 8959
rect 16405 8925 16439 8959
rect 16681 8925 16715 8959
rect 17417 8925 17451 8959
rect 17601 8925 17635 8959
rect 18429 8925 18463 8959
rect 20821 8925 20855 8959
rect 20913 8925 20947 8959
rect 21097 8925 21131 8959
rect 21281 8925 21315 8959
rect 15485 8857 15519 8891
rect 18613 8857 18647 8891
rect 15761 8789 15795 8823
rect 16221 8789 16255 8823
rect 16589 8789 16623 8823
rect 20637 8789 20671 8823
rect 4353 8585 4387 8619
rect 8033 8585 8067 8619
rect 10885 8585 10919 8619
rect 12817 8585 12851 8619
rect 13369 8585 13403 8619
rect 17877 8585 17911 8619
rect 19533 8585 19567 8619
rect 20453 8585 20487 8619
rect 5466 8517 5500 8551
rect 6920 8517 6954 8551
rect 20621 8517 20655 8551
rect 20821 8517 20855 8551
rect 5733 8449 5767 8483
rect 6653 8449 6687 8483
rect 9505 8449 9539 8483
rect 9781 8449 9815 8483
rect 12725 8449 12759 8483
rect 13645 8449 13679 8483
rect 14657 8449 14691 8483
rect 14842 8449 14876 8483
rect 14933 8449 14967 8483
rect 15209 8449 15243 8483
rect 15853 8449 15887 8483
rect 15945 8449 15979 8483
rect 16865 8449 16899 8483
rect 17049 8449 17083 8483
rect 17509 8449 17543 8483
rect 18889 8449 18923 8483
rect 19073 8449 19107 8483
rect 19165 8449 19199 8483
rect 19257 8449 19291 8483
rect 13553 8381 13587 8415
rect 13921 8381 13955 8415
rect 14013 8381 14047 8415
rect 16957 8381 16991 8415
rect 17601 8381 17635 8415
rect 15117 8245 15151 8279
rect 15945 8245 15979 8279
rect 17601 8245 17635 8279
rect 20637 8245 20671 8279
rect 10977 8041 11011 8075
rect 14933 8041 14967 8075
rect 17417 8041 17451 8075
rect 19809 8041 19843 8075
rect 17049 7973 17083 8007
rect 9597 7905 9631 7939
rect 15301 7905 15335 7939
rect 20637 7905 20671 7939
rect 2329 7837 2363 7871
rect 2513 7837 2547 7871
rect 12909 7837 12943 7871
rect 13277 7837 13311 7871
rect 13369 7837 13403 7871
rect 15117 7837 15151 7871
rect 20085 7837 20119 7871
rect 20545 7837 20579 7871
rect 20729 7837 20763 7871
rect 5733 7769 5767 7803
rect 7481 7769 7515 7803
rect 9864 7769 9898 7803
rect 13093 7769 13127 7803
rect 19809 7769 19843 7803
rect 2421 7701 2455 7735
rect 12633 7701 12667 7735
rect 13001 7701 13035 7735
rect 17417 7701 17451 7735
rect 17601 7701 17635 7735
rect 19993 7701 20027 7735
rect 2881 7497 2915 7531
rect 17601 7497 17635 7531
rect 19809 7497 19843 7531
rect 4353 7429 4387 7463
rect 9505 7429 9539 7463
rect 17877 7429 17911 7463
rect 7849 7361 7883 7395
rect 12725 7361 12759 7395
rect 12909 7361 12943 7395
rect 13001 7361 13035 7395
rect 15117 7361 15151 7395
rect 17693 7361 17727 7395
rect 19717 7361 19751 7395
rect 20361 7361 20395 7395
rect 20545 7361 20579 7395
rect 12817 7293 12851 7327
rect 12541 7157 12575 7191
rect 15209 7157 15243 7191
rect 20361 7157 20395 7191
rect 17509 6953 17543 6987
rect 18429 6953 18463 6987
rect 18797 6885 18831 6919
rect 13553 6817 13587 6851
rect 14289 6817 14323 6851
rect 15209 6817 15243 6851
rect 16313 6817 16347 6851
rect 17601 6817 17635 6851
rect 17693 6817 17727 6851
rect 18521 6817 18555 6851
rect 19809 6817 19843 6851
rect 19901 6817 19935 6851
rect 1685 6749 1719 6783
rect 1952 6749 1986 6783
rect 5733 6749 5767 6783
rect 6929 6749 6963 6783
rect 9505 6749 9539 6783
rect 11437 6749 11471 6783
rect 11704 6749 11738 6783
rect 13277 6749 13311 6783
rect 13369 6749 13403 6783
rect 15117 6749 15151 6783
rect 16589 6749 16623 6783
rect 17380 6749 17414 6783
rect 18429 6749 18463 6783
rect 19625 6749 19659 6783
rect 19717 6749 19751 6783
rect 5466 6681 5500 6715
rect 7196 6681 7230 6715
rect 9772 6681 9806 6715
rect 16773 6681 16807 6715
rect 17233 6681 17267 6715
rect 3065 6613 3099 6647
rect 4353 6613 4387 6647
rect 8309 6613 8343 6647
rect 10885 6613 10919 6647
rect 12817 6613 12851 6647
rect 13277 6613 13311 6647
rect 19441 6613 19475 6647
rect 3157 6409 3191 6443
rect 17417 6409 17451 6443
rect 18521 6409 18555 6443
rect 19717 6409 19751 6443
rect 10977 6341 11011 6375
rect 1777 6273 1811 6307
rect 2044 6273 2078 6307
rect 3985 6273 4019 6307
rect 6828 6273 6862 6307
rect 9321 6273 9355 6307
rect 9597 6273 9631 6307
rect 12817 6273 12851 6307
rect 13093 6273 13127 6307
rect 13277 6273 13311 6307
rect 13829 6273 13863 6307
rect 14105 6273 14139 6307
rect 15669 6273 15703 6307
rect 15853 6273 15887 6307
rect 16129 6273 16163 6307
rect 16957 6273 16991 6307
rect 17233 6273 17267 6307
rect 18153 6273 18187 6307
rect 18245 6273 18279 6307
rect 19349 6273 19383 6307
rect 19487 6273 19521 6307
rect 19809 6273 19843 6307
rect 4261 6205 4295 6239
rect 6561 6205 6595 6239
rect 12633 6205 12667 6239
rect 16221 6205 16255 6239
rect 19625 6205 19659 6239
rect 13829 6137 13863 6171
rect 17049 6137 17083 6171
rect 5549 6069 5583 6103
rect 7941 6069 7975 6103
rect 18153 6069 18187 6103
rect 4353 5865 4387 5899
rect 14473 5865 14507 5899
rect 15945 5865 15979 5899
rect 16129 5865 16163 5899
rect 10977 5797 11011 5831
rect 3157 5729 3191 5763
rect 5733 5729 5767 5763
rect 14657 5729 14691 5763
rect 5477 5661 5511 5695
rect 9413 5661 9447 5695
rect 9689 5661 9723 5695
rect 13001 5661 13035 5695
rect 13185 5661 13219 5695
rect 14749 5661 14783 5695
rect 14841 5661 14875 5695
rect 14933 5661 14967 5695
rect 2912 5593 2946 5627
rect 15761 5593 15795 5627
rect 1777 5525 1811 5559
rect 12817 5525 12851 5559
rect 15961 5525 15995 5559
rect 3065 5321 3099 5355
rect 13645 5321 13679 5355
rect 18153 5321 18187 5355
rect 4353 5253 4387 5287
rect 7849 5253 7883 5287
rect 9505 5253 9539 5287
rect 13553 5185 13587 5219
rect 13749 5185 13783 5219
rect 14933 5185 14967 5219
rect 16865 5185 16899 5219
rect 17233 5185 17267 5219
rect 17509 5185 17543 5219
rect 14565 5117 14599 5151
rect 14657 5049 14691 5083
rect 14768 5049 14802 5083
rect 14289 4981 14323 5015
rect 8401 4777 8435 4811
rect 15761 4777 15795 4811
rect 17325 4777 17359 4811
rect 13093 4709 13127 4743
rect 17141 4709 17175 4743
rect 5181 4641 5215 4675
rect 9597 4641 9631 4675
rect 15209 4641 15243 4675
rect 16865 4641 16899 4675
rect 1869 4573 1903 4607
rect 7021 4573 7055 4607
rect 12817 4573 12851 4607
rect 12909 4573 12943 4607
rect 13185 4573 13219 4607
rect 14473 4573 14507 4607
rect 14841 4573 14875 4607
rect 14933 4573 14967 4607
rect 15301 4573 15335 4607
rect 2136 4505 2170 4539
rect 5448 4505 5482 4539
rect 7288 4505 7322 4539
rect 9864 4505 9898 4539
rect 3249 4437 3283 4471
rect 6561 4437 6595 4471
rect 10977 4437 11011 4471
rect 12633 4437 12667 4471
rect 12265 4233 12299 4267
rect 12725 4233 12759 4267
rect 9956 4165 9990 4199
rect 1685 4097 1719 4131
rect 1952 4097 1986 4131
rect 4261 4097 4295 4131
rect 4528 4097 4562 4131
rect 7113 4097 7147 4131
rect 7380 4097 7414 4131
rect 9689 4097 9723 4131
rect 12633 4097 12667 4131
rect 14749 4097 14783 4131
rect 14841 4097 14875 4131
rect 15025 4097 15059 4131
rect 15117 4097 15151 4131
rect 15209 4097 15243 4131
rect 12817 4029 12851 4063
rect 11069 3961 11103 3995
rect 15393 3961 15427 3995
rect 3065 3893 3099 3927
rect 5641 3893 5675 3927
rect 8493 3893 8527 3927
rect 4813 3689 4847 3723
rect 14565 3689 14599 3723
rect 15209 3689 15243 3723
rect 11621 3621 11655 3655
rect 2329 3553 2363 3587
rect 2605 3553 2639 3587
rect 4997 3553 5031 3587
rect 6009 3553 6043 3587
rect 8125 3553 8159 3587
rect 2237 3485 2271 3519
rect 5089 3485 5123 3519
rect 5917 3485 5951 3519
rect 7941 3485 7975 3519
rect 10885 3485 10919 3519
rect 11345 3485 11379 3519
rect 11621 3485 11655 3519
rect 13277 3485 13311 3519
rect 14473 3485 14507 3519
rect 14657 3485 14691 3519
rect 15117 3485 15151 3519
rect 5365 3417 5399 3451
rect 5457 3417 5491 3451
rect 7757 3417 7791 3451
rect 10640 3417 10674 3451
rect 13093 3417 13127 3451
rect 9505 3349 9539 3383
rect 11437 3349 11471 3383
rect 13461 3349 13495 3383
rect 2513 3145 2547 3179
rect 7665 3145 7699 3179
rect 8033 3145 8067 3179
rect 8125 3145 8159 3179
rect 10057 3145 10091 3179
rect 15301 3145 15335 3179
rect 5733 3077 5767 3111
rect 10701 3077 10735 3111
rect 2697 3009 2731 3043
rect 2789 3009 2823 3043
rect 3065 3009 3099 3043
rect 4169 3009 4203 3043
rect 4353 3009 4387 3043
rect 9045 3009 9079 3043
rect 10333 3009 10367 3043
rect 12081 3009 12115 3043
rect 12173 3009 12207 3043
rect 12909 3009 12943 3043
rect 13093 3009 13127 3043
rect 13185 3009 13219 3043
rect 13277 3009 13311 3043
rect 13395 3009 13429 3043
rect 13553 3009 13587 3043
rect 14473 3009 14507 3043
rect 14657 3009 14691 3043
rect 15209 3009 15243 3043
rect 4813 2941 4847 2975
rect 5365 2941 5399 2975
rect 8217 2941 8251 2975
rect 9321 2941 9355 2975
rect 10241 2941 10275 2975
rect 10609 2941 10643 2975
rect 12357 2941 12391 2975
rect 5181 2873 5215 2907
rect 11713 2873 11747 2907
rect 14657 2873 14691 2907
rect 2973 2805 3007 2839
rect 4353 2805 4387 2839
rect 5273 2805 5307 2839
rect 8861 2805 8895 2839
rect 9229 2805 9263 2839
rect 2329 2601 2363 2635
rect 4353 2601 4387 2635
rect 5733 2601 5767 2635
rect 7205 2601 7239 2635
rect 9229 2601 9263 2635
rect 12541 2601 12575 2635
rect 13461 2601 13495 2635
rect 2789 2533 2823 2567
rect 4813 2465 4847 2499
rect 4997 2465 5031 2499
rect 7849 2465 7883 2499
rect 10793 2465 10827 2499
rect 13461 2465 13495 2499
rect 2513 2397 2547 2431
rect 2605 2397 2639 2431
rect 2881 2397 2915 2431
rect 4721 2397 4755 2431
rect 5825 2397 5859 2431
rect 7573 2397 7607 2431
rect 7665 2397 7699 2431
rect 9137 2397 9171 2431
rect 9321 2397 9355 2431
rect 10977 2397 11011 2431
rect 12449 2397 12483 2431
rect 12633 2397 12667 2431
rect 13093 2397 13127 2431
rect 11161 2329 11195 2363
rect 13277 2261 13311 2295
<< metal1 >>
rect 1104 21786 22976 21808
rect 1104 21734 6378 21786
rect 6430 21734 6442 21786
rect 6494 21734 6506 21786
rect 6558 21734 6570 21786
rect 6622 21734 6634 21786
rect 6686 21734 11806 21786
rect 11858 21734 11870 21786
rect 11922 21734 11934 21786
rect 11986 21734 11998 21786
rect 12050 21734 12062 21786
rect 12114 21734 17234 21786
rect 17286 21734 17298 21786
rect 17350 21734 17362 21786
rect 17414 21734 17426 21786
rect 17478 21734 17490 21786
rect 17542 21734 22662 21786
rect 22714 21734 22726 21786
rect 22778 21734 22790 21786
rect 22842 21734 22854 21786
rect 22906 21734 22918 21786
rect 22970 21734 22976 21786
rect 1104 21712 22976 21734
rect 1104 21242 22816 21264
rect 1104 21190 3664 21242
rect 3716 21190 3728 21242
rect 3780 21190 3792 21242
rect 3844 21190 3856 21242
rect 3908 21190 3920 21242
rect 3972 21190 9092 21242
rect 9144 21190 9156 21242
rect 9208 21190 9220 21242
rect 9272 21190 9284 21242
rect 9336 21190 9348 21242
rect 9400 21190 14520 21242
rect 14572 21190 14584 21242
rect 14636 21190 14648 21242
rect 14700 21190 14712 21242
rect 14764 21190 14776 21242
rect 14828 21190 19948 21242
rect 20000 21190 20012 21242
rect 20064 21190 20076 21242
rect 20128 21190 20140 21242
rect 20192 21190 20204 21242
rect 20256 21190 22816 21242
rect 1104 21168 22816 21190
rect 1104 20698 22976 20720
rect 1104 20646 6378 20698
rect 6430 20646 6442 20698
rect 6494 20646 6506 20698
rect 6558 20646 6570 20698
rect 6622 20646 6634 20698
rect 6686 20646 11806 20698
rect 11858 20646 11870 20698
rect 11922 20646 11934 20698
rect 11986 20646 11998 20698
rect 12050 20646 12062 20698
rect 12114 20646 17234 20698
rect 17286 20646 17298 20698
rect 17350 20646 17362 20698
rect 17414 20646 17426 20698
rect 17478 20646 17490 20698
rect 17542 20646 22662 20698
rect 22714 20646 22726 20698
rect 22778 20646 22790 20698
rect 22842 20646 22854 20698
rect 22906 20646 22918 20698
rect 22970 20646 22976 20698
rect 1104 20624 22976 20646
rect 1104 20154 22816 20176
rect 1104 20102 3664 20154
rect 3716 20102 3728 20154
rect 3780 20102 3792 20154
rect 3844 20102 3856 20154
rect 3908 20102 3920 20154
rect 3972 20102 9092 20154
rect 9144 20102 9156 20154
rect 9208 20102 9220 20154
rect 9272 20102 9284 20154
rect 9336 20102 9348 20154
rect 9400 20102 14520 20154
rect 14572 20102 14584 20154
rect 14636 20102 14648 20154
rect 14700 20102 14712 20154
rect 14764 20102 14776 20154
rect 14828 20102 19948 20154
rect 20000 20102 20012 20154
rect 20064 20102 20076 20154
rect 20128 20102 20140 20154
rect 20192 20102 20204 20154
rect 20256 20102 22816 20154
rect 1104 20080 22816 20102
rect 934 19796 940 19848
rect 992 19836 998 19848
rect 1765 19839 1823 19845
rect 1765 19836 1777 19839
rect 992 19808 1777 19836
rect 992 19796 998 19808
rect 1765 19805 1777 19808
rect 1811 19805 1823 19839
rect 1765 19799 1823 19805
rect 2041 19839 2099 19845
rect 2041 19805 2053 19839
rect 2087 19805 2099 19839
rect 2041 19799 2099 19805
rect 1578 19728 1584 19780
rect 1636 19768 1642 19780
rect 2056 19768 2084 19799
rect 1636 19740 2084 19768
rect 1636 19728 1642 19740
rect 1104 19610 22976 19632
rect 1104 19558 6378 19610
rect 6430 19558 6442 19610
rect 6494 19558 6506 19610
rect 6558 19558 6570 19610
rect 6622 19558 6634 19610
rect 6686 19558 11806 19610
rect 11858 19558 11870 19610
rect 11922 19558 11934 19610
rect 11986 19558 11998 19610
rect 12050 19558 12062 19610
rect 12114 19558 17234 19610
rect 17286 19558 17298 19610
rect 17350 19558 17362 19610
rect 17414 19558 17426 19610
rect 17478 19558 17490 19610
rect 17542 19558 22662 19610
rect 22714 19558 22726 19610
rect 22778 19558 22790 19610
rect 22842 19558 22854 19610
rect 22906 19558 22918 19610
rect 22970 19558 22976 19610
rect 1104 19536 22976 19558
rect 1104 19066 22816 19088
rect 1104 19014 3664 19066
rect 3716 19014 3728 19066
rect 3780 19014 3792 19066
rect 3844 19014 3856 19066
rect 3908 19014 3920 19066
rect 3972 19014 9092 19066
rect 9144 19014 9156 19066
rect 9208 19014 9220 19066
rect 9272 19014 9284 19066
rect 9336 19014 9348 19066
rect 9400 19014 14520 19066
rect 14572 19014 14584 19066
rect 14636 19014 14648 19066
rect 14700 19014 14712 19066
rect 14764 19014 14776 19066
rect 14828 19014 19948 19066
rect 20000 19014 20012 19066
rect 20064 19014 20076 19066
rect 20128 19014 20140 19066
rect 20192 19014 20204 19066
rect 20256 19014 22816 19066
rect 1104 18992 22816 19014
rect 1104 18522 22976 18544
rect 1104 18470 6378 18522
rect 6430 18470 6442 18522
rect 6494 18470 6506 18522
rect 6558 18470 6570 18522
rect 6622 18470 6634 18522
rect 6686 18470 11806 18522
rect 11858 18470 11870 18522
rect 11922 18470 11934 18522
rect 11986 18470 11998 18522
rect 12050 18470 12062 18522
rect 12114 18470 17234 18522
rect 17286 18470 17298 18522
rect 17350 18470 17362 18522
rect 17414 18470 17426 18522
rect 17478 18470 17490 18522
rect 17542 18470 22662 18522
rect 22714 18470 22726 18522
rect 22778 18470 22790 18522
rect 22842 18470 22854 18522
rect 22906 18470 22918 18522
rect 22970 18470 22976 18522
rect 1104 18448 22976 18470
rect 8846 18232 8852 18284
rect 8904 18232 8910 18284
rect 9033 18275 9091 18281
rect 9033 18241 9045 18275
rect 9079 18241 9091 18275
rect 9033 18235 9091 18241
rect 8386 18164 8392 18216
rect 8444 18204 8450 18216
rect 9048 18204 9076 18235
rect 8444 18176 9076 18204
rect 8444 18164 8450 18176
rect 8938 18028 8944 18080
rect 8996 18028 9002 18080
rect 1104 17978 22816 18000
rect 1104 17926 3664 17978
rect 3716 17926 3728 17978
rect 3780 17926 3792 17978
rect 3844 17926 3856 17978
rect 3908 17926 3920 17978
rect 3972 17926 9092 17978
rect 9144 17926 9156 17978
rect 9208 17926 9220 17978
rect 9272 17926 9284 17978
rect 9336 17926 9348 17978
rect 9400 17926 14520 17978
rect 14572 17926 14584 17978
rect 14636 17926 14648 17978
rect 14700 17926 14712 17978
rect 14764 17926 14776 17978
rect 14828 17926 19948 17978
rect 20000 17926 20012 17978
rect 20064 17926 20076 17978
rect 20128 17926 20140 17978
rect 20192 17926 20204 17978
rect 20256 17926 22816 17978
rect 1104 17904 22816 17926
rect 8938 17796 8944 17808
rect 7116 17768 8944 17796
rect 5353 17731 5411 17737
rect 5353 17697 5365 17731
rect 5399 17728 5411 17731
rect 5718 17728 5724 17740
rect 5399 17700 5724 17728
rect 5399 17697 5411 17700
rect 5353 17691 5411 17697
rect 5718 17688 5724 17700
rect 5776 17688 5782 17740
rect 7006 17620 7012 17672
rect 7064 17620 7070 17672
rect 7116 17669 7144 17768
rect 8938 17756 8944 17768
rect 8996 17756 9002 17808
rect 9306 17756 9312 17808
rect 9364 17796 9370 17808
rect 9364 17768 10732 17796
rect 9364 17756 9370 17768
rect 8021 17731 8079 17737
rect 8021 17697 8033 17731
rect 8067 17728 8079 17731
rect 9398 17728 9404 17740
rect 8067 17700 9404 17728
rect 8067 17697 8079 17700
rect 8021 17691 8079 17697
rect 9398 17688 9404 17700
rect 9456 17688 9462 17740
rect 10704 17737 10732 17768
rect 10689 17731 10747 17737
rect 10689 17697 10701 17731
rect 10735 17728 10747 17731
rect 10870 17728 10876 17740
rect 10735 17700 10876 17728
rect 10735 17697 10747 17700
rect 10689 17691 10747 17697
rect 10870 17688 10876 17700
rect 10928 17688 10934 17740
rect 7101 17663 7159 17669
rect 7101 17629 7113 17663
rect 7147 17629 7159 17663
rect 7101 17623 7159 17629
rect 7190 17620 7196 17672
rect 7248 17620 7254 17672
rect 8202 17620 8208 17672
rect 8260 17620 8266 17672
rect 8294 17620 8300 17672
rect 8352 17620 8358 17672
rect 8846 17620 8852 17672
rect 8904 17660 8910 17672
rect 9306 17660 9312 17672
rect 8904 17632 9312 17660
rect 8904 17620 8910 17632
rect 9306 17620 9312 17632
rect 9364 17620 9370 17672
rect 9493 17663 9551 17669
rect 9493 17629 9505 17663
rect 9539 17629 9551 17663
rect 9493 17623 9551 17629
rect 5169 17595 5227 17601
rect 5169 17561 5181 17595
rect 5215 17592 5227 17595
rect 8021 17595 8079 17601
rect 8021 17592 8033 17595
rect 5215 17564 8033 17592
rect 5215 17561 5227 17564
rect 5169 17555 5227 17561
rect 8021 17561 8033 17564
rect 8067 17561 8079 17595
rect 9508 17592 9536 17623
rect 9950 17620 9956 17672
rect 10008 17660 10014 17672
rect 10413 17663 10471 17669
rect 10413 17660 10425 17663
rect 10008 17632 10425 17660
rect 10008 17620 10014 17632
rect 10413 17629 10425 17632
rect 10459 17629 10471 17663
rect 10413 17623 10471 17629
rect 10505 17663 10563 17669
rect 10505 17629 10517 17663
rect 10551 17660 10563 17663
rect 10594 17660 10600 17672
rect 10551 17632 10600 17660
rect 10551 17629 10563 17632
rect 10505 17623 10563 17629
rect 10520 17592 10548 17623
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 9508 17564 10548 17592
rect 8021 17555 8079 17561
rect 4706 17484 4712 17536
rect 4764 17484 4770 17536
rect 4890 17484 4896 17536
rect 4948 17524 4954 17536
rect 5077 17527 5135 17533
rect 5077 17524 5089 17527
rect 4948 17496 5089 17524
rect 4948 17484 4954 17496
rect 5077 17493 5089 17496
rect 5123 17493 5135 17527
rect 5077 17487 5135 17493
rect 6825 17527 6883 17533
rect 6825 17493 6837 17527
rect 6871 17524 6883 17527
rect 7098 17524 7104 17536
rect 6871 17496 7104 17524
rect 6871 17493 6883 17496
rect 6825 17487 6883 17493
rect 7098 17484 7104 17496
rect 7156 17484 7162 17536
rect 9401 17527 9459 17533
rect 9401 17493 9413 17527
rect 9447 17524 9459 17527
rect 9490 17524 9496 17536
rect 9447 17496 9496 17524
rect 9447 17493 9459 17496
rect 9401 17487 9459 17493
rect 9490 17484 9496 17496
rect 9548 17484 9554 17536
rect 10594 17484 10600 17536
rect 10652 17524 10658 17536
rect 10689 17527 10747 17533
rect 10689 17524 10701 17527
rect 10652 17496 10701 17524
rect 10652 17484 10658 17496
rect 10689 17493 10701 17496
rect 10735 17493 10747 17527
rect 10689 17487 10747 17493
rect 1104 17434 22976 17456
rect 1104 17382 6378 17434
rect 6430 17382 6442 17434
rect 6494 17382 6506 17434
rect 6558 17382 6570 17434
rect 6622 17382 6634 17434
rect 6686 17382 11806 17434
rect 11858 17382 11870 17434
rect 11922 17382 11934 17434
rect 11986 17382 11998 17434
rect 12050 17382 12062 17434
rect 12114 17382 17234 17434
rect 17286 17382 17298 17434
rect 17350 17382 17362 17434
rect 17414 17382 17426 17434
rect 17478 17382 17490 17434
rect 17542 17382 22662 17434
rect 22714 17382 22726 17434
rect 22778 17382 22790 17434
rect 22842 17382 22854 17434
rect 22906 17382 22918 17434
rect 22970 17382 22976 17434
rect 1104 17360 22976 17382
rect 5261 17323 5319 17329
rect 5261 17289 5273 17323
rect 5307 17320 5319 17323
rect 6917 17323 6975 17329
rect 6917 17320 6929 17323
rect 5307 17292 6929 17320
rect 5307 17289 5319 17292
rect 5261 17283 5319 17289
rect 6917 17289 6929 17292
rect 6963 17289 6975 17323
rect 6917 17283 6975 17289
rect 8110 17280 8116 17332
rect 8168 17320 8174 17332
rect 8846 17320 8852 17332
rect 8168 17292 8852 17320
rect 8168 17280 8174 17292
rect 8846 17280 8852 17292
rect 8904 17280 8910 17332
rect 9398 17280 9404 17332
rect 9456 17280 9462 17332
rect 7006 17212 7012 17264
rect 7064 17252 7070 17264
rect 7285 17255 7343 17261
rect 7285 17252 7297 17255
rect 7064 17224 7297 17252
rect 7064 17212 7070 17224
rect 7285 17221 7297 17224
rect 7331 17252 7343 17255
rect 7929 17255 7987 17261
rect 7929 17252 7941 17255
rect 7331 17224 7941 17252
rect 7331 17221 7343 17224
rect 7285 17215 7343 17221
rect 7929 17221 7941 17224
rect 7975 17221 7987 17255
rect 7929 17215 7987 17221
rect 8036 17224 8984 17252
rect 3053 17187 3111 17193
rect 3053 17153 3065 17187
rect 3099 17184 3111 17187
rect 3326 17184 3332 17196
rect 3099 17156 3332 17184
rect 3099 17153 3111 17156
rect 3053 17147 3111 17153
rect 3326 17144 3332 17156
rect 3384 17144 3390 17196
rect 5074 17144 5080 17196
rect 5132 17184 5138 17196
rect 5169 17187 5227 17193
rect 5169 17184 5181 17187
rect 5132 17156 5181 17184
rect 5132 17144 5138 17156
rect 5169 17153 5181 17156
rect 5215 17153 5227 17187
rect 5169 17147 5227 17153
rect 7101 17187 7159 17193
rect 7101 17153 7113 17187
rect 7147 17153 7159 17187
rect 7101 17147 7159 17153
rect 3145 17119 3203 17125
rect 3145 17085 3157 17119
rect 3191 17085 3203 17119
rect 3145 17079 3203 17085
rect 3160 17048 3188 17079
rect 3234 17076 3240 17128
rect 3292 17116 3298 17128
rect 5353 17119 5411 17125
rect 5353 17116 5365 17119
rect 3292 17088 5365 17116
rect 3292 17076 3298 17088
rect 5353 17085 5365 17088
rect 5399 17116 5411 17119
rect 5718 17116 5724 17128
rect 5399 17088 5724 17116
rect 5399 17085 5411 17088
rect 5353 17079 5411 17085
rect 5718 17076 5724 17088
rect 5776 17076 5782 17128
rect 7116 17116 7144 17147
rect 7190 17144 7196 17196
rect 7248 17144 7254 17196
rect 7469 17187 7527 17193
rect 7469 17153 7481 17187
rect 7515 17184 7527 17187
rect 8036 17184 8064 17224
rect 8956 17196 8984 17224
rect 7515 17156 8064 17184
rect 7515 17153 7527 17156
rect 7469 17147 7527 17153
rect 8110 17144 8116 17196
rect 8168 17144 8174 17196
rect 8297 17187 8355 17193
rect 8297 17184 8309 17187
rect 8220 17156 8309 17184
rect 8220 17116 8248 17156
rect 8297 17153 8309 17156
rect 8343 17184 8355 17187
rect 8386 17184 8392 17196
rect 8343 17156 8392 17184
rect 8343 17153 8355 17156
rect 8297 17147 8355 17153
rect 8386 17144 8392 17156
rect 8444 17144 8450 17196
rect 8938 17144 8944 17196
rect 8996 17184 9002 17196
rect 9585 17187 9643 17193
rect 9585 17184 9597 17187
rect 8996 17156 9597 17184
rect 8996 17144 9002 17156
rect 9585 17153 9597 17156
rect 9631 17153 9643 17187
rect 9585 17147 9643 17153
rect 9674 17144 9680 17196
rect 9732 17144 9738 17196
rect 9861 17187 9919 17193
rect 9861 17153 9873 17187
rect 9907 17153 9919 17187
rect 9861 17147 9919 17153
rect 9876 17116 9904 17147
rect 9950 17144 9956 17196
rect 10008 17144 10014 17196
rect 10597 17187 10655 17193
rect 10597 17153 10609 17187
rect 10643 17184 10655 17187
rect 10686 17184 10692 17196
rect 10643 17156 10692 17184
rect 10643 17153 10655 17156
rect 10597 17147 10655 17153
rect 10686 17144 10692 17156
rect 10744 17144 10750 17196
rect 10413 17119 10471 17125
rect 10413 17116 10425 17119
rect 7116 17088 8248 17116
rect 8312 17088 10425 17116
rect 8312 17060 8340 17088
rect 10413 17085 10425 17088
rect 10459 17085 10471 17119
rect 10413 17079 10471 17085
rect 10781 17119 10839 17125
rect 10781 17085 10793 17119
rect 10827 17116 10839 17119
rect 10870 17116 10876 17128
rect 10827 17088 10876 17116
rect 10827 17085 10839 17088
rect 10781 17079 10839 17085
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 3160 17020 8156 17048
rect 2682 16940 2688 16992
rect 2740 16940 2746 16992
rect 4798 16940 4804 16992
rect 4856 16940 4862 16992
rect 8128 16980 8156 17020
rect 8294 17008 8300 17060
rect 8352 17008 8358 17060
rect 10502 16980 10508 16992
rect 8128 16952 10508 16980
rect 10502 16940 10508 16952
rect 10560 16940 10566 16992
rect 1104 16890 22816 16912
rect 1104 16838 3664 16890
rect 3716 16838 3728 16890
rect 3780 16838 3792 16890
rect 3844 16838 3856 16890
rect 3908 16838 3920 16890
rect 3972 16838 9092 16890
rect 9144 16838 9156 16890
rect 9208 16838 9220 16890
rect 9272 16838 9284 16890
rect 9336 16838 9348 16890
rect 9400 16838 14520 16890
rect 14572 16838 14584 16890
rect 14636 16838 14648 16890
rect 14700 16838 14712 16890
rect 14764 16838 14776 16890
rect 14828 16838 19948 16890
rect 20000 16838 20012 16890
rect 20064 16838 20076 16890
rect 20128 16838 20140 16890
rect 20192 16838 20204 16890
rect 20256 16838 22816 16890
rect 1104 16816 22816 16838
rect 7466 16776 7472 16788
rect 6932 16748 7472 16776
rect 6825 16711 6883 16717
rect 6825 16708 6837 16711
rect 3068 16680 6837 16708
rect 3068 16649 3096 16680
rect 6825 16677 6837 16680
rect 6871 16677 6883 16711
rect 6825 16671 6883 16677
rect 3053 16643 3111 16649
rect 3053 16609 3065 16643
rect 3099 16609 3111 16643
rect 3053 16603 3111 16609
rect 3237 16643 3295 16649
rect 3237 16609 3249 16643
rect 3283 16640 3295 16643
rect 3283 16612 4844 16640
rect 3283 16609 3295 16612
rect 3237 16603 3295 16609
rect 4816 16504 4844 16612
rect 4890 16600 4896 16652
rect 4948 16640 4954 16652
rect 4948 16612 5028 16640
rect 4948 16600 4954 16612
rect 5000 16581 5028 16612
rect 5718 16600 5724 16652
rect 5776 16640 5782 16652
rect 6730 16640 6736 16652
rect 5776 16612 6736 16640
rect 5776 16600 5782 16612
rect 6730 16600 6736 16612
rect 6788 16600 6794 16652
rect 4985 16575 5043 16581
rect 4985 16541 4997 16575
rect 5031 16541 5043 16575
rect 4985 16535 5043 16541
rect 5074 16532 5080 16584
rect 5132 16572 5138 16584
rect 5261 16575 5319 16581
rect 5261 16572 5273 16575
rect 5132 16544 5273 16572
rect 5132 16532 5138 16544
rect 5261 16541 5273 16544
rect 5307 16541 5319 16575
rect 5261 16535 5319 16541
rect 5626 16532 5632 16584
rect 5684 16532 5690 16584
rect 6365 16575 6423 16581
rect 6365 16541 6377 16575
rect 6411 16572 6423 16575
rect 6932 16572 6960 16748
rect 7466 16736 7472 16748
rect 7524 16736 7530 16788
rect 8294 16736 8300 16788
rect 8352 16776 8358 16788
rect 9309 16779 9367 16785
rect 9309 16776 9321 16779
rect 8352 16748 9321 16776
rect 8352 16736 8358 16748
rect 9309 16745 9321 16748
rect 9355 16745 9367 16779
rect 9309 16739 9367 16745
rect 10502 16736 10508 16788
rect 10560 16776 10566 16788
rect 10597 16779 10655 16785
rect 10597 16776 10609 16779
rect 10560 16748 10609 16776
rect 10560 16736 10566 16748
rect 10597 16745 10609 16748
rect 10643 16745 10655 16779
rect 10597 16739 10655 16745
rect 7190 16668 7196 16720
rect 7248 16708 7254 16720
rect 9950 16708 9956 16720
rect 7248 16680 8156 16708
rect 7248 16668 7254 16680
rect 7929 16643 7987 16649
rect 7929 16640 7941 16643
rect 7024 16612 7941 16640
rect 7024 16581 7052 16612
rect 7929 16609 7941 16612
rect 7975 16609 7987 16643
rect 7929 16603 7987 16609
rect 8128 16640 8156 16680
rect 9140 16680 9956 16708
rect 9140 16649 9168 16680
rect 9950 16668 9956 16680
rect 10008 16668 10014 16720
rect 9125 16643 9183 16649
rect 9125 16640 9137 16643
rect 8128 16612 9137 16640
rect 8128 16584 8156 16612
rect 9125 16609 9137 16612
rect 9171 16609 9183 16643
rect 9125 16603 9183 16609
rect 9674 16600 9680 16652
rect 9732 16640 9738 16652
rect 9732 16612 10916 16640
rect 9732 16600 9738 16612
rect 6411 16544 6960 16572
rect 7009 16575 7067 16581
rect 6411 16541 6423 16544
rect 6365 16535 6423 16541
rect 7009 16541 7021 16575
rect 7055 16541 7067 16575
rect 7009 16535 7067 16541
rect 7282 16532 7288 16584
rect 7340 16581 7346 16584
rect 7340 16575 7369 16581
rect 7357 16541 7369 16575
rect 7340 16535 7369 16541
rect 7340 16532 7346 16535
rect 7466 16532 7472 16584
rect 7524 16532 7530 16584
rect 8110 16532 8116 16584
rect 8168 16532 8174 16584
rect 9401 16575 9459 16581
rect 9401 16541 9413 16575
rect 9447 16572 9459 16575
rect 9490 16572 9496 16584
rect 9447 16544 9496 16572
rect 9447 16541 9459 16544
rect 9401 16535 9459 16541
rect 9490 16532 9496 16544
rect 9548 16532 9554 16584
rect 10594 16532 10600 16584
rect 10652 16532 10658 16584
rect 10888 16581 10916 16612
rect 10873 16575 10931 16581
rect 10873 16541 10885 16575
rect 10919 16572 10931 16575
rect 10962 16572 10968 16584
rect 10919 16544 10968 16572
rect 10919 16541 10931 16544
rect 10873 16535 10931 16541
rect 10962 16532 10968 16544
rect 11020 16532 11026 16584
rect 5166 16504 5172 16516
rect 4816 16476 5172 16504
rect 5166 16464 5172 16476
rect 5224 16464 5230 16516
rect 7101 16507 7159 16513
rect 7101 16473 7113 16507
rect 7147 16473 7159 16507
rect 7101 16467 7159 16473
rect 2590 16396 2596 16448
rect 2648 16396 2654 16448
rect 2961 16439 3019 16445
rect 2961 16405 2973 16439
rect 3007 16436 3019 16439
rect 3326 16436 3332 16448
rect 3007 16408 3332 16436
rect 3007 16405 3019 16408
rect 2961 16399 3019 16405
rect 3326 16396 3332 16408
rect 3384 16396 3390 16448
rect 7116 16436 7144 16467
rect 7190 16464 7196 16516
rect 7248 16464 7254 16516
rect 8297 16507 8355 16513
rect 8297 16473 8309 16507
rect 8343 16504 8355 16507
rect 8386 16504 8392 16516
rect 8343 16476 8392 16504
rect 8343 16473 8355 16476
rect 8297 16467 8355 16473
rect 8386 16464 8392 16476
rect 8444 16504 8450 16516
rect 10410 16504 10416 16516
rect 8444 16476 10416 16504
rect 8444 16464 8450 16476
rect 10410 16464 10416 16476
rect 10468 16504 10474 16516
rect 10689 16507 10747 16513
rect 10689 16504 10701 16507
rect 10468 16476 10701 16504
rect 10468 16464 10474 16476
rect 10689 16473 10701 16476
rect 10735 16473 10747 16507
rect 10689 16467 10747 16473
rect 9125 16439 9183 16445
rect 9125 16436 9137 16439
rect 7116 16408 9137 16436
rect 9125 16405 9137 16408
rect 9171 16405 9183 16439
rect 9125 16399 9183 16405
rect 1104 16346 22976 16368
rect 1104 16294 6378 16346
rect 6430 16294 6442 16346
rect 6494 16294 6506 16346
rect 6558 16294 6570 16346
rect 6622 16294 6634 16346
rect 6686 16294 11806 16346
rect 11858 16294 11870 16346
rect 11922 16294 11934 16346
rect 11986 16294 11998 16346
rect 12050 16294 12062 16346
rect 12114 16294 17234 16346
rect 17286 16294 17298 16346
rect 17350 16294 17362 16346
rect 17414 16294 17426 16346
rect 17478 16294 17490 16346
rect 17542 16294 22662 16346
rect 22714 16294 22726 16346
rect 22778 16294 22790 16346
rect 22842 16294 22854 16346
rect 22906 16294 22918 16346
rect 22970 16294 22976 16346
rect 1104 16272 22976 16294
rect 2593 16235 2651 16241
rect 2593 16201 2605 16235
rect 2639 16232 2651 16235
rect 2682 16232 2688 16244
rect 2639 16204 2688 16232
rect 2639 16201 2651 16204
rect 2593 16195 2651 16201
rect 2682 16192 2688 16204
rect 2740 16192 2746 16244
rect 4798 16192 4804 16244
rect 4856 16232 4862 16244
rect 4893 16235 4951 16241
rect 4893 16232 4905 16235
rect 4856 16204 4905 16232
rect 4856 16192 4862 16204
rect 4893 16201 4905 16204
rect 4939 16201 4951 16235
rect 4893 16195 4951 16201
rect 6914 16192 6920 16244
rect 6972 16232 6978 16244
rect 7190 16232 7196 16244
rect 6972 16204 7196 16232
rect 6972 16192 6978 16204
rect 7190 16192 7196 16204
rect 7248 16192 7254 16244
rect 7466 16192 7472 16244
rect 7524 16232 7530 16244
rect 14366 16232 14372 16244
rect 7524 16204 14372 16232
rect 7524 16192 7530 16204
rect 14366 16192 14372 16204
rect 14424 16192 14430 16244
rect 10045 16167 10103 16173
rect 10045 16133 10057 16167
rect 10091 16164 10103 16167
rect 10134 16164 10140 16176
rect 10091 16136 10140 16164
rect 10091 16133 10103 16136
rect 10045 16127 10103 16133
rect 10134 16124 10140 16136
rect 10192 16124 10198 16176
rect 10597 16167 10655 16173
rect 10597 16133 10609 16167
rect 10643 16164 10655 16167
rect 10686 16164 10692 16176
rect 10643 16136 10692 16164
rect 10643 16133 10655 16136
rect 10597 16127 10655 16133
rect 10686 16124 10692 16136
rect 10744 16164 10750 16176
rect 11793 16167 11851 16173
rect 11793 16164 11805 16167
rect 10744 16136 11805 16164
rect 10744 16124 10750 16136
rect 11793 16133 11805 16136
rect 11839 16133 11851 16167
rect 11793 16127 11851 16133
rect 2501 16099 2559 16105
rect 2501 16065 2513 16099
rect 2547 16096 2559 16099
rect 3050 16096 3056 16108
rect 2547 16068 3056 16096
rect 2547 16065 2559 16068
rect 2501 16059 2559 16065
rect 3050 16056 3056 16068
rect 3108 16056 3114 16108
rect 4801 16099 4859 16105
rect 4801 16065 4813 16099
rect 4847 16096 4859 16099
rect 5258 16096 5264 16108
rect 4847 16068 5264 16096
rect 4847 16065 4859 16068
rect 4801 16059 4859 16065
rect 5258 16056 5264 16068
rect 5316 16056 5322 16108
rect 8297 16099 8355 16105
rect 8297 16065 8309 16099
rect 8343 16096 8355 16099
rect 9490 16096 9496 16108
rect 8343 16068 9496 16096
rect 8343 16065 8355 16068
rect 8297 16059 8355 16065
rect 9490 16056 9496 16068
rect 9548 16056 9554 16108
rect 9674 16056 9680 16108
rect 9732 16096 9738 16108
rect 9732 16068 10180 16096
rect 9732 16056 9738 16068
rect 2682 15988 2688 16040
rect 2740 15988 2746 16040
rect 5077 16031 5135 16037
rect 5077 15997 5089 16031
rect 5123 16028 5135 16031
rect 5166 16028 5172 16040
rect 5123 16000 5172 16028
rect 5123 15997 5135 16000
rect 5077 15991 5135 15997
rect 5166 15988 5172 16000
rect 5224 15988 5230 16040
rect 8110 15988 8116 16040
rect 8168 15988 8174 16040
rect 8386 15988 8392 16040
rect 8444 15988 8450 16040
rect 10152 16037 10180 16068
rect 11054 16056 11060 16108
rect 11112 16096 11118 16108
rect 11701 16099 11759 16105
rect 11701 16096 11713 16099
rect 11112 16068 11713 16096
rect 11112 16056 11118 16068
rect 11701 16065 11713 16068
rect 11747 16065 11759 16099
rect 11701 16059 11759 16065
rect 11885 16099 11943 16105
rect 11885 16065 11897 16099
rect 11931 16065 11943 16099
rect 11885 16059 11943 16065
rect 8481 16031 8539 16037
rect 8481 15997 8493 16031
rect 8527 15997 8539 16031
rect 8481 15991 8539 15997
rect 8573 16031 8631 16037
rect 8573 15997 8585 16031
rect 8619 16028 8631 16031
rect 9861 16031 9919 16037
rect 9861 16028 9873 16031
rect 8619 16000 9873 16028
rect 8619 15997 8631 16000
rect 8573 15991 8631 15997
rect 9861 15997 9873 16000
rect 9907 15997 9919 16031
rect 9861 15991 9919 15997
rect 10137 16031 10195 16037
rect 10137 15997 10149 16031
rect 10183 15997 10195 16031
rect 10137 15991 10195 15997
rect 8128 15960 8156 15988
rect 8496 15960 8524 15991
rect 10318 15988 10324 16040
rect 10376 16028 10382 16040
rect 11900 16028 11928 16059
rect 10376 16000 11928 16028
rect 10376 15988 10382 16000
rect 10597 15963 10655 15969
rect 10597 15960 10609 15963
rect 8128 15932 10609 15960
rect 10597 15929 10609 15932
rect 10643 15929 10655 15963
rect 10597 15923 10655 15929
rect 2038 15852 2044 15904
rect 2096 15892 2102 15904
rect 2133 15895 2191 15901
rect 2133 15892 2145 15895
rect 2096 15864 2145 15892
rect 2096 15852 2102 15864
rect 2133 15861 2145 15864
rect 2179 15861 2191 15895
rect 2133 15855 2191 15861
rect 4433 15895 4491 15901
rect 4433 15861 4445 15895
rect 4479 15892 4491 15895
rect 4522 15892 4528 15904
rect 4479 15864 4528 15892
rect 4479 15861 4491 15864
rect 4433 15855 4491 15861
rect 4522 15852 4528 15864
rect 4580 15852 4586 15904
rect 7190 15852 7196 15904
rect 7248 15892 7254 15904
rect 8113 15895 8171 15901
rect 8113 15892 8125 15895
rect 7248 15864 8125 15892
rect 7248 15852 7254 15864
rect 8113 15861 8125 15864
rect 8159 15861 8171 15895
rect 8113 15855 8171 15861
rect 1104 15802 22816 15824
rect 1104 15750 3664 15802
rect 3716 15750 3728 15802
rect 3780 15750 3792 15802
rect 3844 15750 3856 15802
rect 3908 15750 3920 15802
rect 3972 15750 9092 15802
rect 9144 15750 9156 15802
rect 9208 15750 9220 15802
rect 9272 15750 9284 15802
rect 9336 15750 9348 15802
rect 9400 15750 14520 15802
rect 14572 15750 14584 15802
rect 14636 15750 14648 15802
rect 14700 15750 14712 15802
rect 14764 15750 14776 15802
rect 14828 15750 19948 15802
rect 20000 15750 20012 15802
rect 20064 15750 20076 15802
rect 20128 15750 20140 15802
rect 20192 15750 20204 15802
rect 20256 15750 22816 15802
rect 1104 15728 22816 15750
rect 10410 15648 10416 15700
rect 10468 15648 10474 15700
rect 10962 15580 10968 15632
rect 11020 15580 11026 15632
rect 4706 15512 4712 15564
rect 4764 15552 4770 15564
rect 4801 15555 4859 15561
rect 4801 15552 4813 15555
rect 4764 15524 4813 15552
rect 4764 15512 4770 15524
rect 4801 15521 4813 15524
rect 4847 15521 4859 15555
rect 4801 15515 4859 15521
rect 4985 15555 5043 15561
rect 4985 15521 4997 15555
rect 5031 15552 5043 15555
rect 5166 15552 5172 15564
rect 5031 15524 5172 15552
rect 5031 15521 5043 15524
rect 4985 15515 5043 15521
rect 5166 15512 5172 15524
rect 5224 15512 5230 15564
rect 6914 15444 6920 15496
rect 6972 15484 6978 15496
rect 7009 15487 7067 15493
rect 7009 15484 7021 15487
rect 6972 15456 7021 15484
rect 6972 15444 6978 15456
rect 7009 15453 7021 15456
rect 7055 15453 7067 15487
rect 7009 15447 7067 15453
rect 7190 15444 7196 15496
rect 7248 15444 7254 15496
rect 9309 15487 9367 15493
rect 9309 15453 9321 15487
rect 9355 15453 9367 15487
rect 9309 15447 9367 15453
rect 9324 15416 9352 15447
rect 10318 15444 10324 15496
rect 10376 15444 10382 15496
rect 10505 15487 10563 15493
rect 10505 15453 10517 15487
rect 10551 15484 10563 15487
rect 11054 15484 11060 15496
rect 10551 15456 11060 15484
rect 10551 15453 10563 15456
rect 10505 15447 10563 15453
rect 11054 15444 11060 15456
rect 11112 15484 11118 15496
rect 11333 15487 11391 15493
rect 11333 15484 11345 15487
rect 11112 15456 11345 15484
rect 11112 15444 11118 15456
rect 11333 15453 11345 15456
rect 11379 15453 11391 15487
rect 11333 15447 11391 15453
rect 10870 15416 10876 15428
rect 9324 15388 10876 15416
rect 10870 15376 10876 15388
rect 10928 15416 10934 15428
rect 11149 15419 11207 15425
rect 11149 15416 11161 15419
rect 10928 15388 11161 15416
rect 10928 15376 10934 15388
rect 11149 15385 11161 15388
rect 11195 15385 11207 15419
rect 11149 15379 11207 15385
rect 4341 15351 4399 15357
rect 4341 15317 4353 15351
rect 4387 15348 4399 15351
rect 4430 15348 4436 15360
rect 4387 15320 4436 15348
rect 4387 15317 4399 15320
rect 4341 15311 4399 15317
rect 4430 15308 4436 15320
rect 4488 15308 4494 15360
rect 4709 15351 4767 15357
rect 4709 15317 4721 15351
rect 4755 15348 4767 15351
rect 5074 15348 5080 15360
rect 4755 15320 5080 15348
rect 4755 15317 4767 15320
rect 4709 15311 4767 15317
rect 5074 15308 5080 15320
rect 5132 15308 5138 15360
rect 5534 15308 5540 15360
rect 5592 15348 5598 15360
rect 7009 15351 7067 15357
rect 7009 15348 7021 15351
rect 5592 15320 7021 15348
rect 5592 15308 5598 15320
rect 7009 15317 7021 15320
rect 7055 15317 7067 15351
rect 7009 15311 7067 15317
rect 9214 15308 9220 15360
rect 9272 15308 9278 15360
rect 1104 15258 22976 15280
rect 1104 15206 6378 15258
rect 6430 15206 6442 15258
rect 6494 15206 6506 15258
rect 6558 15206 6570 15258
rect 6622 15206 6634 15258
rect 6686 15206 11806 15258
rect 11858 15206 11870 15258
rect 11922 15206 11934 15258
rect 11986 15206 11998 15258
rect 12050 15206 12062 15258
rect 12114 15206 17234 15258
rect 17286 15206 17298 15258
rect 17350 15206 17362 15258
rect 17414 15206 17426 15258
rect 17478 15206 17490 15258
rect 17542 15206 22662 15258
rect 22714 15206 22726 15258
rect 22778 15206 22790 15258
rect 22842 15206 22854 15258
rect 22906 15206 22918 15258
rect 22970 15206 22976 15258
rect 1104 15184 22976 15206
rect 8021 15147 8079 15153
rect 8021 15113 8033 15147
rect 8067 15144 8079 15147
rect 8110 15144 8116 15156
rect 8067 15116 8116 15144
rect 8067 15113 8079 15116
rect 8021 15107 8079 15113
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 8202 15104 8208 15156
rect 8260 15144 8266 15156
rect 8665 15147 8723 15153
rect 8665 15144 8677 15147
rect 8260 15116 8677 15144
rect 8260 15104 8266 15116
rect 8665 15113 8677 15116
rect 8711 15113 8723 15147
rect 8665 15107 8723 15113
rect 2041 15079 2099 15085
rect 2041 15045 2053 15079
rect 2087 15076 2099 15079
rect 2406 15076 2412 15088
rect 2087 15048 2412 15076
rect 2087 15045 2099 15048
rect 2041 15039 2099 15045
rect 2406 15036 2412 15048
rect 2464 15036 2470 15088
rect 3234 15076 3240 15088
rect 2746 15048 3240 15076
rect 1854 14968 1860 15020
rect 1912 14968 1918 15020
rect 2130 14968 2136 15020
rect 2188 15008 2194 15020
rect 2746 15008 2774 15048
rect 3234 15036 3240 15048
rect 3292 15036 3298 15088
rect 4709 15079 4767 15085
rect 4709 15045 4721 15079
rect 4755 15076 4767 15079
rect 5534 15076 5540 15088
rect 4755 15048 5540 15076
rect 4755 15045 4767 15048
rect 4709 15039 4767 15045
rect 5534 15036 5540 15048
rect 5592 15036 5598 15088
rect 7009 15079 7067 15085
rect 7009 15045 7021 15079
rect 7055 15076 7067 15079
rect 9953 15079 10011 15085
rect 9953 15076 9965 15079
rect 7055 15048 9965 15076
rect 7055 15045 7067 15048
rect 7009 15039 7067 15045
rect 9953 15045 9965 15048
rect 9999 15045 10011 15079
rect 10965 15079 11023 15085
rect 10965 15076 10977 15079
rect 9953 15039 10011 15045
rect 10152 15048 10977 15076
rect 10152 15020 10180 15048
rect 10965 15045 10977 15048
rect 11011 15045 11023 15079
rect 10965 15039 11023 15045
rect 2188 14980 2774 15008
rect 2961 15011 3019 15017
rect 2188 14968 2194 14980
rect 2961 14977 2973 15011
rect 3007 15008 3019 15011
rect 3050 15008 3056 15020
rect 3007 14980 3056 15008
rect 3007 14977 3019 14980
rect 2961 14971 3019 14977
rect 3050 14968 3056 14980
rect 3108 14968 3114 15020
rect 3145 15011 3203 15017
rect 3145 14977 3157 15011
rect 3191 15008 3203 15011
rect 3326 15008 3332 15020
rect 3191 14980 3332 15008
rect 3191 14977 3203 14980
rect 3145 14971 3203 14977
rect 3326 14968 3332 14980
rect 3384 14968 3390 15020
rect 4062 14968 4068 15020
rect 4120 15008 4126 15020
rect 4525 15011 4583 15017
rect 4525 15008 4537 15011
rect 4120 14980 4537 15008
rect 4120 14968 4126 14980
rect 4525 14977 4537 14980
rect 4571 14977 4583 15011
rect 4525 14971 4583 14977
rect 4798 14968 4804 15020
rect 4856 14968 4862 15020
rect 4890 14968 4896 15020
rect 4948 14968 4954 15020
rect 5258 14968 5264 15020
rect 5316 15008 5322 15020
rect 6917 15011 6975 15017
rect 6917 15008 6929 15011
rect 5316 14980 6929 15008
rect 5316 14968 5322 14980
rect 6917 14977 6929 14980
rect 6963 14977 6975 15011
rect 6917 14971 6975 14977
rect 8113 15011 8171 15017
rect 8113 14977 8125 15011
rect 8159 15008 8171 15011
rect 8294 15008 8300 15020
rect 8159 14980 8300 15008
rect 8159 14977 8171 14980
rect 8113 14971 8171 14977
rect 8294 14968 8300 14980
rect 8352 14968 8358 15020
rect 8938 14968 8944 15020
rect 8996 15008 9002 15020
rect 9214 15008 9220 15020
rect 8996 14980 9220 15008
rect 8996 14968 9002 14980
rect 9214 14968 9220 14980
rect 9272 14968 9278 15020
rect 10134 14968 10140 15020
rect 10192 14968 10198 15020
rect 10413 15011 10471 15017
rect 10413 15008 10425 15011
rect 10244 14980 10425 15008
rect 7006 14900 7012 14952
rect 7064 14940 7070 14952
rect 7101 14943 7159 14949
rect 7101 14940 7113 14943
rect 7064 14912 7113 14940
rect 7064 14900 7070 14912
rect 7101 14909 7113 14912
rect 7147 14909 7159 14943
rect 7101 14903 7159 14909
rect 8846 14900 8852 14952
rect 8904 14900 8910 14952
rect 9309 14943 9367 14949
rect 9309 14909 9321 14943
rect 9355 14909 9367 14943
rect 9309 14903 9367 14909
rect 8110 14832 8116 14884
rect 8168 14872 8174 14884
rect 9324 14872 9352 14903
rect 9490 14900 9496 14952
rect 9548 14940 9554 14952
rect 10045 14943 10103 14949
rect 10045 14940 10057 14943
rect 9548 14912 10057 14940
rect 9548 14900 9554 14912
rect 10045 14909 10057 14912
rect 10091 14909 10103 14943
rect 10045 14903 10103 14909
rect 10244 14872 10272 14980
rect 10413 14977 10425 14980
rect 10459 14977 10471 15011
rect 10413 14971 10471 14977
rect 10870 14968 10876 15020
rect 10928 14968 10934 15020
rect 11054 14968 11060 15020
rect 11112 14968 11118 15020
rect 10321 14943 10379 14949
rect 10321 14909 10333 14943
rect 10367 14940 10379 14943
rect 10962 14940 10968 14952
rect 10367 14912 10968 14940
rect 10367 14909 10379 14912
rect 10321 14903 10379 14909
rect 10962 14900 10968 14912
rect 11020 14900 11026 14952
rect 8168 14844 10272 14872
rect 8168 14832 8174 14844
rect 1762 14764 1768 14816
rect 1820 14804 1826 14816
rect 1857 14807 1915 14813
rect 1857 14804 1869 14807
rect 1820 14776 1869 14804
rect 1820 14764 1826 14776
rect 1857 14773 1869 14776
rect 1903 14773 1915 14807
rect 1857 14767 1915 14773
rect 3053 14807 3111 14813
rect 3053 14773 3065 14807
rect 3099 14804 3111 14807
rect 3418 14804 3424 14816
rect 3099 14776 3424 14804
rect 3099 14773 3111 14776
rect 3053 14767 3111 14773
rect 3418 14764 3424 14776
rect 3476 14764 3482 14816
rect 5077 14807 5135 14813
rect 5077 14773 5089 14807
rect 5123 14804 5135 14807
rect 5534 14804 5540 14816
rect 5123 14776 5540 14804
rect 5123 14773 5135 14776
rect 5077 14767 5135 14773
rect 5534 14764 5540 14776
rect 5592 14764 5598 14816
rect 6549 14807 6607 14813
rect 6549 14773 6561 14807
rect 6595 14804 6607 14807
rect 6638 14804 6644 14816
rect 6595 14776 6644 14804
rect 6595 14773 6607 14776
rect 6549 14767 6607 14773
rect 6638 14764 6644 14776
rect 6696 14764 6702 14816
rect 1104 14714 22816 14736
rect 1104 14662 3664 14714
rect 3716 14662 3728 14714
rect 3780 14662 3792 14714
rect 3844 14662 3856 14714
rect 3908 14662 3920 14714
rect 3972 14662 9092 14714
rect 9144 14662 9156 14714
rect 9208 14662 9220 14714
rect 9272 14662 9284 14714
rect 9336 14662 9348 14714
rect 9400 14662 14520 14714
rect 14572 14662 14584 14714
rect 14636 14662 14648 14714
rect 14700 14662 14712 14714
rect 14764 14662 14776 14714
rect 14828 14662 19948 14714
rect 20000 14662 20012 14714
rect 20064 14662 20076 14714
rect 20128 14662 20140 14714
rect 20192 14662 20204 14714
rect 20256 14662 22816 14714
rect 1104 14640 22816 14662
rect 1578 14560 1584 14612
rect 1636 14600 1642 14612
rect 1765 14603 1823 14609
rect 1765 14600 1777 14603
rect 1636 14572 1777 14600
rect 1636 14560 1642 14572
rect 1765 14569 1777 14572
rect 1811 14569 1823 14603
rect 1765 14563 1823 14569
rect 3973 14603 4031 14609
rect 3973 14569 3985 14603
rect 4019 14600 4031 14603
rect 4062 14600 4068 14612
rect 4019 14572 4068 14600
rect 4019 14569 4031 14572
rect 3973 14563 4031 14569
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 5077 14603 5135 14609
rect 5077 14569 5089 14603
rect 5123 14569 5135 14603
rect 5077 14563 5135 14569
rect 3329 14535 3387 14541
rect 3329 14501 3341 14535
rect 3375 14532 3387 14535
rect 3510 14532 3516 14544
rect 3375 14504 3516 14532
rect 3375 14501 3387 14504
rect 3329 14495 3387 14501
rect 3510 14492 3516 14504
rect 3568 14532 3574 14544
rect 5092 14532 5120 14563
rect 5166 14560 5172 14612
rect 5224 14600 5230 14612
rect 5224 14572 6592 14600
rect 5224 14560 5230 14572
rect 3568 14504 5120 14532
rect 3568 14492 3574 14504
rect 4338 14424 4344 14476
rect 4396 14424 4402 14476
rect 6564 14473 6592 14572
rect 9490 14560 9496 14612
rect 9548 14560 9554 14612
rect 8846 14492 8852 14544
rect 8904 14532 8910 14544
rect 8904 14504 9628 14532
rect 8904 14492 8910 14504
rect 6549 14467 6607 14473
rect 5000 14436 6500 14464
rect 1949 14399 2007 14405
rect 1949 14365 1961 14399
rect 1995 14365 2007 14399
rect 1949 14359 2007 14365
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14396 2191 14399
rect 2406 14396 2412 14408
rect 2179 14368 2412 14396
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 1964 14328 1992 14359
rect 2406 14356 2412 14368
rect 2464 14356 2470 14408
rect 2682 14356 2688 14408
rect 2740 14396 2746 14408
rect 5000 14405 5028 14436
rect 4157 14399 4215 14405
rect 4157 14396 4169 14399
rect 2740 14368 4169 14396
rect 2740 14356 2746 14368
rect 4157 14365 4169 14368
rect 4203 14365 4215 14399
rect 4157 14359 4215 14365
rect 4433 14399 4491 14405
rect 4433 14365 4445 14399
rect 4479 14365 4491 14399
rect 4433 14359 4491 14365
rect 4985 14399 5043 14405
rect 4985 14365 4997 14399
rect 5031 14365 5043 14399
rect 4985 14359 5043 14365
rect 5169 14399 5227 14405
rect 5169 14365 5181 14399
rect 5215 14390 5227 14399
rect 5258 14390 5264 14408
rect 5215 14365 5264 14390
rect 5169 14362 5264 14365
rect 5169 14359 5227 14362
rect 2314 14328 2320 14340
rect 1964 14300 2320 14328
rect 2314 14288 2320 14300
rect 2372 14288 2378 14340
rect 2961 14331 3019 14337
rect 2961 14297 2973 14331
rect 3007 14328 3019 14331
rect 3050 14328 3056 14340
rect 3007 14300 3056 14328
rect 3007 14297 3019 14300
rect 2961 14291 3019 14297
rect 3050 14288 3056 14300
rect 3108 14288 3114 14340
rect 3145 14331 3203 14337
rect 3145 14297 3157 14331
rect 3191 14328 3203 14331
rect 3326 14328 3332 14340
rect 3191 14300 3332 14328
rect 3191 14297 3203 14300
rect 3145 14291 3203 14297
rect 3326 14288 3332 14300
rect 3384 14288 3390 14340
rect 4172 14260 4200 14359
rect 4448 14328 4476 14359
rect 5258 14356 5264 14362
rect 5316 14356 5322 14408
rect 5350 14356 5356 14408
rect 5408 14396 5414 14408
rect 5537 14399 5595 14405
rect 5537 14396 5549 14399
rect 5408 14368 5549 14396
rect 5408 14356 5414 14368
rect 5537 14365 5549 14368
rect 5583 14365 5595 14399
rect 5537 14359 5595 14365
rect 5810 14328 5816 14340
rect 4448 14300 5816 14328
rect 5810 14288 5816 14300
rect 5868 14288 5874 14340
rect 6472 14328 6500 14436
rect 6549 14433 6561 14467
rect 6595 14433 6607 14467
rect 6549 14427 6607 14433
rect 6564 14396 6592 14427
rect 6638 14424 6644 14476
rect 6696 14424 6702 14476
rect 8294 14424 8300 14476
rect 8352 14464 8358 14476
rect 9600 14473 9628 14504
rect 9401 14467 9459 14473
rect 9401 14464 9413 14467
rect 8352 14436 9413 14464
rect 8352 14424 8358 14436
rect 9401 14433 9413 14436
rect 9447 14433 9459 14467
rect 9401 14427 9459 14433
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14464 9643 14467
rect 9674 14464 9680 14476
rect 9631 14436 9680 14464
rect 9631 14433 9643 14436
rect 9585 14427 9643 14433
rect 9674 14424 9680 14436
rect 9732 14464 9738 14476
rect 10318 14464 10324 14476
rect 9732 14436 10324 14464
rect 9732 14424 9738 14436
rect 10318 14424 10324 14436
rect 10376 14424 10382 14476
rect 6564 14368 8156 14396
rect 6733 14331 6791 14337
rect 6733 14328 6745 14331
rect 6472 14300 6745 14328
rect 6733 14297 6745 14300
rect 6779 14328 6791 14331
rect 7374 14328 7380 14340
rect 6779 14300 7380 14328
rect 6779 14297 6791 14300
rect 6733 14291 6791 14297
rect 7374 14288 7380 14300
rect 7432 14328 7438 14340
rect 8018 14328 8024 14340
rect 7432 14300 8024 14328
rect 7432 14288 7438 14300
rect 8018 14288 8024 14300
rect 8076 14288 8082 14340
rect 8128 14328 8156 14368
rect 8938 14356 8944 14408
rect 8996 14396 9002 14408
rect 9309 14399 9367 14405
rect 9309 14396 9321 14399
rect 8996 14368 9321 14396
rect 8996 14356 9002 14368
rect 9309 14365 9321 14368
rect 9355 14365 9367 14399
rect 9309 14359 9367 14365
rect 9490 14356 9496 14408
rect 9548 14396 9554 14408
rect 11333 14399 11391 14405
rect 11333 14396 11345 14399
rect 9548 14368 11345 14396
rect 9548 14356 9554 14368
rect 11333 14365 11345 14368
rect 11379 14396 11391 14399
rect 11514 14396 11520 14408
rect 11379 14368 11520 14396
rect 11379 14365 11391 14368
rect 11333 14359 11391 14365
rect 11514 14356 11520 14368
rect 11572 14356 11578 14408
rect 10502 14328 10508 14340
rect 8128 14300 10508 14328
rect 10502 14288 10508 14300
rect 10560 14288 10566 14340
rect 10778 14288 10784 14340
rect 10836 14288 10842 14340
rect 5166 14260 5172 14272
rect 4172 14232 5172 14260
rect 5166 14220 5172 14232
rect 5224 14220 5230 14272
rect 5353 14263 5411 14269
rect 5353 14229 5365 14263
rect 5399 14260 5411 14263
rect 5626 14260 5632 14272
rect 5399 14232 5632 14260
rect 5399 14229 5411 14232
rect 5353 14223 5411 14229
rect 5626 14220 5632 14232
rect 5684 14220 5690 14272
rect 7101 14263 7159 14269
rect 7101 14229 7113 14263
rect 7147 14260 7159 14263
rect 7282 14260 7288 14272
rect 7147 14232 7288 14260
rect 7147 14229 7159 14232
rect 7101 14223 7159 14229
rect 7282 14220 7288 14232
rect 7340 14220 7346 14272
rect 1104 14170 22976 14192
rect 1104 14118 6378 14170
rect 6430 14118 6442 14170
rect 6494 14118 6506 14170
rect 6558 14118 6570 14170
rect 6622 14118 6634 14170
rect 6686 14118 11806 14170
rect 11858 14118 11870 14170
rect 11922 14118 11934 14170
rect 11986 14118 11998 14170
rect 12050 14118 12062 14170
rect 12114 14118 17234 14170
rect 17286 14118 17298 14170
rect 17350 14118 17362 14170
rect 17414 14118 17426 14170
rect 17478 14118 17490 14170
rect 17542 14118 22662 14170
rect 22714 14118 22726 14170
rect 22778 14118 22790 14170
rect 22842 14118 22854 14170
rect 22906 14118 22918 14170
rect 22970 14118 22976 14170
rect 1104 14096 22976 14118
rect 1854 14016 1860 14068
rect 1912 14056 1918 14068
rect 2317 14059 2375 14065
rect 2317 14056 2329 14059
rect 1912 14028 2329 14056
rect 1912 14016 1918 14028
rect 2317 14025 2329 14028
rect 2363 14025 2375 14059
rect 2317 14019 2375 14025
rect 3598 14059 3656 14065
rect 3598 14025 3610 14059
rect 3644 14056 3656 14059
rect 5261 14059 5319 14065
rect 3644 14028 5212 14056
rect 3644 14025 3656 14028
rect 3598 14019 3656 14025
rect 2406 13988 2412 14000
rect 2056 13960 2412 13988
rect 2056 13929 2084 13960
rect 2406 13948 2412 13960
rect 2464 13948 2470 14000
rect 3697 13991 3755 13997
rect 3697 13988 3709 13991
rect 2746 13960 3709 13988
rect 2041 13923 2099 13929
rect 2041 13889 2053 13923
rect 2087 13889 2099 13923
rect 2041 13883 2099 13889
rect 2130 13880 2136 13932
rect 2188 13920 2194 13932
rect 2746 13920 2774 13960
rect 3697 13957 3709 13960
rect 3743 13957 3755 13991
rect 3697 13951 3755 13957
rect 4338 13948 4344 14000
rect 4396 13988 4402 14000
rect 4982 13988 4988 14000
rect 4396 13960 4988 13988
rect 4396 13948 4402 13960
rect 2188 13892 2774 13920
rect 2188 13880 2194 13892
rect 3418 13880 3424 13932
rect 3476 13880 3482 13932
rect 3510 13880 3516 13932
rect 3568 13880 3574 13932
rect 2317 13855 2375 13861
rect 2317 13821 2329 13855
rect 2363 13852 2375 13855
rect 2682 13852 2688 13864
rect 2363 13824 2688 13852
rect 2363 13821 2375 13824
rect 2317 13815 2375 13821
rect 2682 13812 2688 13824
rect 2740 13812 2746 13864
rect 4540 13852 4568 13960
rect 4982 13948 4988 13960
rect 5040 13948 5046 14000
rect 5184 13988 5212 14028
rect 5261 14025 5273 14059
rect 5307 14056 5319 14059
rect 7193 14059 7251 14065
rect 7193 14056 7205 14059
rect 5307 14028 7205 14056
rect 5307 14025 5319 14028
rect 5261 14019 5319 14025
rect 7193 14025 7205 14028
rect 7239 14025 7251 14059
rect 7193 14019 7251 14025
rect 5184 13960 6684 13988
rect 4617 13923 4675 13929
rect 4617 13889 4629 13923
rect 4663 13920 4675 13923
rect 5442 13920 5448 13932
rect 4663 13892 5448 13920
rect 4663 13889 4675 13892
rect 4617 13883 4675 13889
rect 5442 13880 5448 13892
rect 5500 13880 5506 13932
rect 6656 13929 6684 13960
rect 6822 13948 6828 14000
rect 6880 13948 6886 14000
rect 6917 13991 6975 13997
rect 6917 13957 6929 13991
rect 6963 13988 6975 13991
rect 8202 13988 8208 14000
rect 6963 13960 8208 13988
rect 6963 13957 6975 13960
rect 6917 13951 6975 13957
rect 8202 13948 8208 13960
rect 8260 13948 8266 14000
rect 9217 13991 9275 13997
rect 9217 13988 9229 13991
rect 8312 13960 9229 13988
rect 6549 13923 6607 13929
rect 6549 13920 6561 13923
rect 5552 13892 6561 13920
rect 4801 13855 4859 13861
rect 4801 13852 4813 13855
rect 4540 13824 4813 13852
rect 4801 13821 4813 13824
rect 4847 13821 4859 13855
rect 4801 13815 4859 13821
rect 4893 13855 4951 13861
rect 4893 13821 4905 13855
rect 4939 13821 4951 13855
rect 4893 13815 4951 13821
rect 4908 13784 4936 13815
rect 4982 13812 4988 13864
rect 5040 13852 5046 13864
rect 5350 13852 5356 13864
rect 5040 13824 5356 13852
rect 5040 13812 5046 13824
rect 5350 13812 5356 13824
rect 5408 13812 5414 13864
rect 5552 13784 5580 13892
rect 6549 13889 6561 13892
rect 6595 13889 6607 13923
rect 6549 13883 6607 13889
rect 6641 13923 6699 13929
rect 6641 13889 6653 13923
rect 6687 13889 6699 13923
rect 6641 13883 6699 13889
rect 7009 13923 7067 13929
rect 7009 13889 7021 13923
rect 7055 13920 7067 13923
rect 7098 13920 7104 13932
rect 7055 13892 7104 13920
rect 7055 13889 7067 13892
rect 7009 13883 7067 13889
rect 7098 13880 7104 13892
rect 7156 13880 7162 13932
rect 8312 13929 8340 13960
rect 9217 13957 9229 13960
rect 9263 13957 9275 13991
rect 9585 13991 9643 13997
rect 9585 13988 9597 13991
rect 9217 13951 9275 13957
rect 9324 13960 9597 13988
rect 8297 13923 8355 13929
rect 8297 13889 8309 13923
rect 8343 13889 8355 13923
rect 8297 13883 8355 13889
rect 8573 13923 8631 13929
rect 8573 13889 8585 13923
rect 8619 13889 8631 13923
rect 8573 13883 8631 13889
rect 8110 13812 8116 13864
rect 8168 13812 8174 13864
rect 8588 13852 8616 13883
rect 8754 13880 8760 13932
rect 8812 13920 8818 13932
rect 9324 13920 9352 13960
rect 9585 13957 9597 13960
rect 9631 13957 9643 13991
rect 9585 13951 9643 13957
rect 8812 13892 9352 13920
rect 9401 13923 9459 13929
rect 8812 13880 8818 13892
rect 9401 13889 9413 13923
rect 9447 13920 9459 13923
rect 9490 13920 9496 13932
rect 9447 13892 9496 13920
rect 9447 13889 9459 13892
rect 9401 13883 9459 13889
rect 9490 13880 9496 13892
rect 9548 13880 9554 13932
rect 9677 13923 9735 13929
rect 9677 13889 9689 13923
rect 9723 13889 9735 13923
rect 9677 13883 9735 13889
rect 8938 13852 8944 13864
rect 8588 13824 8944 13852
rect 8938 13812 8944 13824
rect 8996 13852 9002 13864
rect 9692 13852 9720 13883
rect 10778 13880 10784 13932
rect 10836 13880 10842 13932
rect 13078 13880 13084 13932
rect 13136 13880 13142 13932
rect 13262 13880 13268 13932
rect 13320 13880 13326 13932
rect 13446 13880 13452 13932
rect 13504 13920 13510 13932
rect 15289 13923 15347 13929
rect 15289 13920 15301 13923
rect 13504 13892 15301 13920
rect 13504 13880 13510 13892
rect 15289 13889 15301 13892
rect 15335 13889 15347 13923
rect 15289 13883 15347 13889
rect 8996 13824 9720 13852
rect 10796 13852 10824 13880
rect 13538 13852 13544 13864
rect 10796 13824 13544 13852
rect 8996 13812 9002 13824
rect 13538 13812 13544 13824
rect 13596 13812 13602 13864
rect 13630 13812 13636 13864
rect 13688 13812 13694 13864
rect 15194 13812 15200 13864
rect 15252 13812 15258 13864
rect 4816 13756 5580 13784
rect 15657 13787 15715 13793
rect 4816 13728 4844 13756
rect 15657 13753 15669 13787
rect 15703 13784 15715 13787
rect 16758 13784 16764 13796
rect 15703 13756 16764 13784
rect 15703 13753 15715 13756
rect 15657 13747 15715 13753
rect 16758 13744 16764 13756
rect 16816 13744 16822 13796
rect 4798 13676 4804 13728
rect 4856 13676 4862 13728
rect 10502 13676 10508 13728
rect 10560 13716 10566 13728
rect 10597 13719 10655 13725
rect 10597 13716 10609 13719
rect 10560 13688 10609 13716
rect 10560 13676 10566 13688
rect 10597 13685 10609 13688
rect 10643 13685 10655 13719
rect 10597 13679 10655 13685
rect 1104 13626 22816 13648
rect 1104 13574 3664 13626
rect 3716 13574 3728 13626
rect 3780 13574 3792 13626
rect 3844 13574 3856 13626
rect 3908 13574 3920 13626
rect 3972 13574 9092 13626
rect 9144 13574 9156 13626
rect 9208 13574 9220 13626
rect 9272 13574 9284 13626
rect 9336 13574 9348 13626
rect 9400 13574 14520 13626
rect 14572 13574 14584 13626
rect 14636 13574 14648 13626
rect 14700 13574 14712 13626
rect 14764 13574 14776 13626
rect 14828 13574 19948 13626
rect 20000 13574 20012 13626
rect 20064 13574 20076 13626
rect 20128 13574 20140 13626
rect 20192 13574 20204 13626
rect 20256 13574 22816 13626
rect 1104 13552 22816 13574
rect 13262 13472 13268 13524
rect 13320 13472 13326 13524
rect 14366 13472 14372 13524
rect 14424 13472 14430 13524
rect 17681 13515 17739 13521
rect 17681 13481 17693 13515
rect 17727 13512 17739 13515
rect 19521 13515 19579 13521
rect 19521 13512 19533 13515
rect 17727 13484 19533 13512
rect 17727 13481 17739 13484
rect 17681 13475 17739 13481
rect 19521 13481 19533 13484
rect 19567 13512 19579 13515
rect 19794 13512 19800 13524
rect 19567 13484 19800 13512
rect 19567 13481 19579 13484
rect 19521 13475 19579 13481
rect 19794 13472 19800 13484
rect 19852 13472 19858 13524
rect 15838 13404 15844 13456
rect 15896 13444 15902 13456
rect 17586 13444 17592 13456
rect 15896 13416 17592 13444
rect 15896 13404 15902 13416
rect 17586 13404 17592 13416
rect 17644 13444 17650 13456
rect 17644 13416 17724 13444
rect 17644 13404 17650 13416
rect 2501 13379 2559 13385
rect 2501 13345 2513 13379
rect 2547 13376 2559 13379
rect 2682 13376 2688 13388
rect 2547 13348 2688 13376
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 2682 13336 2688 13348
rect 2740 13376 2746 13388
rect 9490 13376 9496 13388
rect 2740 13348 9496 13376
rect 2740 13336 2746 13348
rect 1854 13268 1860 13320
rect 1912 13308 1918 13320
rect 2225 13311 2283 13317
rect 2225 13308 2237 13311
rect 1912 13280 2237 13308
rect 1912 13268 1918 13280
rect 2225 13277 2237 13280
rect 2271 13277 2283 13311
rect 2225 13271 2283 13277
rect 3142 13268 3148 13320
rect 3200 13268 3206 13320
rect 3237 13311 3295 13317
rect 3237 13277 3249 13311
rect 3283 13308 3295 13311
rect 3602 13308 3608 13320
rect 3283 13280 3608 13308
rect 3283 13277 3295 13280
rect 3237 13271 3295 13277
rect 3602 13268 3608 13280
rect 3660 13268 3666 13320
rect 8938 13268 8944 13320
rect 8996 13308 9002 13320
rect 9324 13317 9352 13348
rect 9490 13336 9496 13348
rect 9548 13336 9554 13388
rect 12069 13379 12127 13385
rect 12069 13376 12081 13379
rect 10704 13348 12081 13376
rect 10704 13320 10732 13348
rect 12069 13345 12081 13348
rect 12115 13345 12127 13379
rect 12069 13339 12127 13345
rect 12805 13379 12863 13385
rect 12805 13345 12817 13379
rect 12851 13376 12863 13379
rect 13814 13376 13820 13388
rect 12851 13348 13820 13376
rect 12851 13345 12863 13348
rect 12805 13339 12863 13345
rect 13814 13336 13820 13348
rect 13872 13336 13878 13388
rect 13906 13336 13912 13388
rect 13964 13376 13970 13388
rect 15565 13379 15623 13385
rect 15565 13376 15577 13379
rect 13964 13348 15577 13376
rect 13964 13336 13970 13348
rect 15565 13345 15577 13348
rect 15611 13376 15623 13379
rect 17034 13376 17040 13388
rect 15611 13348 17040 13376
rect 15611 13345 15623 13348
rect 15565 13339 15623 13345
rect 17034 13336 17040 13348
rect 17092 13336 17098 13388
rect 9125 13311 9183 13317
rect 9125 13308 9137 13311
rect 8996 13280 9137 13308
rect 8996 13268 9002 13280
rect 9125 13277 9137 13280
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13277 9367 13311
rect 9309 13271 9367 13277
rect 10502 13268 10508 13320
rect 10560 13268 10566 13320
rect 10686 13268 10692 13320
rect 10744 13268 10750 13320
rect 10781 13311 10839 13317
rect 10781 13277 10793 13311
rect 10827 13277 10839 13311
rect 10781 13271 10839 13277
rect 10873 13311 10931 13317
rect 10873 13277 10885 13311
rect 10919 13308 10931 13311
rect 11606 13308 11612 13320
rect 10919 13280 11612 13308
rect 10919 13277 10931 13280
rect 10873 13271 10931 13277
rect 3421 13243 3479 13249
rect 3421 13240 3433 13243
rect 2240 13212 3433 13240
rect 2240 13184 2268 13212
rect 3421 13209 3433 13212
rect 3467 13240 3479 13243
rect 4798 13240 4804 13252
rect 3467 13212 4804 13240
rect 3467 13209 3479 13212
rect 3421 13203 3479 13209
rect 4798 13200 4804 13212
rect 4856 13200 4862 13252
rect 10796 13240 10824 13271
rect 11606 13268 11612 13280
rect 11664 13268 11670 13320
rect 11793 13311 11851 13317
rect 11793 13277 11805 13311
rect 11839 13277 11851 13311
rect 11793 13271 11851 13277
rect 12161 13311 12219 13317
rect 12161 13277 12173 13311
rect 12207 13308 12219 13311
rect 12434 13308 12440 13320
rect 12207 13280 12440 13308
rect 12207 13277 12219 13280
rect 12161 13271 12219 13277
rect 10962 13240 10968 13252
rect 10796 13212 10968 13240
rect 10962 13200 10968 13212
rect 11020 13240 11026 13252
rect 11808 13240 11836 13271
rect 12434 13268 12440 13280
rect 12492 13268 12498 13320
rect 13446 13268 13452 13320
rect 13504 13268 13510 13320
rect 13541 13311 13599 13317
rect 13541 13277 13553 13311
rect 13587 13308 13599 13311
rect 13722 13308 13728 13320
rect 13587 13280 13728 13308
rect 13587 13277 13599 13280
rect 13541 13271 13599 13277
rect 13722 13268 13728 13280
rect 13780 13268 13786 13320
rect 13998 13268 14004 13320
rect 14056 13308 14062 13320
rect 14369 13311 14427 13317
rect 14369 13308 14381 13311
rect 14056 13280 14381 13308
rect 14056 13268 14062 13280
rect 14369 13277 14381 13280
rect 14415 13277 14427 13311
rect 14369 13271 14427 13277
rect 15473 13311 15531 13317
rect 15473 13277 15485 13311
rect 15519 13277 15531 13311
rect 15473 13271 15531 13277
rect 11020 13212 11836 13240
rect 11020 13200 11026 13212
rect 13262 13200 13268 13252
rect 13320 13200 13326 13252
rect 13740 13240 13768 13268
rect 15194 13240 15200 13252
rect 13740 13212 15200 13240
rect 15194 13200 15200 13212
rect 15252 13240 15258 13252
rect 15488 13240 15516 13271
rect 16022 13268 16028 13320
rect 16080 13268 16086 13320
rect 16482 13268 16488 13320
rect 16540 13268 16546 13320
rect 16578 13311 16636 13317
rect 16578 13277 16590 13311
rect 16624 13277 16636 13311
rect 16578 13271 16636 13277
rect 17405 13311 17463 13317
rect 17405 13277 17417 13311
rect 17451 13277 17463 13311
rect 17696 13308 17724 13416
rect 17770 13404 17776 13456
rect 17828 13444 17834 13456
rect 17865 13447 17923 13453
rect 17865 13444 17877 13447
rect 17828 13416 17877 13444
rect 17828 13404 17834 13416
rect 17865 13413 17877 13416
rect 17911 13413 17923 13447
rect 17865 13407 17923 13413
rect 18230 13404 18236 13456
rect 18288 13444 18294 13456
rect 18601 13447 18659 13453
rect 18601 13444 18613 13447
rect 18288 13416 18613 13444
rect 18288 13404 18294 13416
rect 18601 13413 18613 13416
rect 18647 13413 18659 13447
rect 18601 13407 18659 13413
rect 17773 13311 17831 13317
rect 17773 13308 17785 13311
rect 17696 13280 17785 13308
rect 17405 13271 17463 13277
rect 17773 13277 17785 13280
rect 17819 13308 17831 13311
rect 18785 13311 18843 13317
rect 18785 13308 18797 13311
rect 17819 13280 18797 13308
rect 17819 13277 17831 13280
rect 17773 13271 17831 13277
rect 18785 13277 18797 13280
rect 18831 13277 18843 13311
rect 18785 13271 18843 13277
rect 18877 13311 18935 13317
rect 18877 13277 18889 13311
rect 18923 13308 18935 13311
rect 19426 13308 19432 13320
rect 18923 13280 19432 13308
rect 18923 13277 18935 13280
rect 18877 13271 18935 13277
rect 16040 13240 16068 13268
rect 16592 13240 16620 13271
rect 15252 13212 15976 13240
rect 16040 13212 16620 13240
rect 17420 13240 17448 13271
rect 17678 13240 17684 13252
rect 17420 13212 17684 13240
rect 15252 13200 15258 13212
rect 2222 13132 2228 13184
rect 2280 13132 2286 13184
rect 2958 13132 2964 13184
rect 3016 13172 3022 13184
rect 3145 13175 3203 13181
rect 3145 13172 3157 13175
rect 3016 13144 3157 13172
rect 3016 13132 3022 13144
rect 3145 13141 3157 13144
rect 3191 13141 3203 13175
rect 3145 13135 3203 13141
rect 8386 13132 8392 13184
rect 8444 13172 8450 13184
rect 9217 13175 9275 13181
rect 9217 13172 9229 13175
rect 8444 13144 9229 13172
rect 8444 13132 8450 13144
rect 9217 13141 9229 13144
rect 9263 13141 9275 13175
rect 9217 13135 9275 13141
rect 9766 13132 9772 13184
rect 9824 13172 9830 13184
rect 11149 13175 11207 13181
rect 11149 13172 11161 13175
rect 9824 13144 11161 13172
rect 9824 13132 9830 13144
rect 11149 13141 11161 13144
rect 11195 13141 11207 13175
rect 11149 13135 11207 13141
rect 15838 13132 15844 13184
rect 15896 13132 15902 13184
rect 15948 13172 15976 13212
rect 17678 13200 17684 13212
rect 17736 13200 17742 13252
rect 18064 13212 18460 13240
rect 16482 13172 16488 13184
rect 15948 13144 16488 13172
rect 16482 13132 16488 13144
rect 16540 13132 16546 13184
rect 16850 13132 16856 13184
rect 16908 13132 16914 13184
rect 17497 13175 17555 13181
rect 17497 13141 17509 13175
rect 17543 13172 17555 13175
rect 18064 13172 18092 13212
rect 17543 13144 18092 13172
rect 18141 13175 18199 13181
rect 17543 13141 17555 13144
rect 17497 13135 17555 13141
rect 18141 13141 18153 13175
rect 18187 13172 18199 13175
rect 18322 13172 18328 13184
rect 18187 13144 18328 13172
rect 18187 13141 18199 13144
rect 18141 13135 18199 13141
rect 18322 13132 18328 13144
rect 18380 13132 18386 13184
rect 18432 13172 18460 13212
rect 18506 13200 18512 13252
rect 18564 13240 18570 13252
rect 18601 13243 18659 13249
rect 18601 13240 18613 13243
rect 18564 13212 18613 13240
rect 18564 13200 18570 13212
rect 18601 13209 18613 13212
rect 18647 13209 18659 13243
rect 18800 13240 18828 13271
rect 19426 13268 19432 13280
rect 19484 13268 19490 13320
rect 19518 13268 19524 13320
rect 19576 13268 19582 13320
rect 19334 13240 19340 13252
rect 18800 13212 19340 13240
rect 18601 13203 18659 13209
rect 19334 13200 19340 13212
rect 19392 13200 19398 13252
rect 20622 13172 20628 13184
rect 18432 13144 20628 13172
rect 20622 13132 20628 13144
rect 20680 13132 20686 13184
rect 1104 13082 22976 13104
rect 1104 13030 6378 13082
rect 6430 13030 6442 13082
rect 6494 13030 6506 13082
rect 6558 13030 6570 13082
rect 6622 13030 6634 13082
rect 6686 13030 11806 13082
rect 11858 13030 11870 13082
rect 11922 13030 11934 13082
rect 11986 13030 11998 13082
rect 12050 13030 12062 13082
rect 12114 13030 17234 13082
rect 17286 13030 17298 13082
rect 17350 13030 17362 13082
rect 17414 13030 17426 13082
rect 17478 13030 17490 13082
rect 17542 13030 22662 13082
rect 22714 13030 22726 13082
rect 22778 13030 22790 13082
rect 22842 13030 22854 13082
rect 22906 13030 22918 13082
rect 22970 13030 22976 13082
rect 1104 13008 22976 13030
rect 3602 12928 3608 12980
rect 3660 12968 3666 12980
rect 4154 12968 4160 12980
rect 3660 12940 4160 12968
rect 3660 12928 3666 12940
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 4632 12940 5856 12968
rect 2866 12860 2872 12912
rect 2924 12900 2930 12912
rect 3237 12903 3295 12909
rect 3237 12900 3249 12903
rect 2924 12872 3249 12900
rect 2924 12860 2930 12872
rect 3237 12869 3249 12872
rect 3283 12869 3295 12903
rect 3237 12863 3295 12869
rect 3418 12860 3424 12912
rect 3476 12909 3482 12912
rect 3476 12903 3495 12909
rect 3483 12869 3495 12903
rect 3476 12863 3495 12869
rect 3476 12860 3482 12863
rect 2682 12792 2688 12844
rect 2740 12792 2746 12844
rect 4632 12841 4660 12940
rect 5718 12860 5724 12912
rect 5776 12860 5782 12912
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 4706 12832 4712 12844
rect 4663 12804 4712 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 4706 12792 4712 12804
rect 4764 12792 4770 12844
rect 4798 12792 4804 12844
rect 4856 12832 4862 12844
rect 5828 12841 5856 12940
rect 8938 12928 8944 12980
rect 8996 12968 9002 12980
rect 9125 12971 9183 12977
rect 9125 12968 9137 12971
rect 8996 12940 9137 12968
rect 8996 12928 9002 12940
rect 9125 12937 9137 12940
rect 9171 12937 9183 12971
rect 10318 12968 10324 12980
rect 9125 12931 9183 12937
rect 9416 12940 10324 12968
rect 7926 12860 7932 12912
rect 7984 12900 7990 12912
rect 9277 12903 9335 12909
rect 9277 12900 9289 12903
rect 7984 12872 9289 12900
rect 7984 12860 7990 12872
rect 9277 12869 9289 12872
rect 9323 12900 9335 12903
rect 9416 12900 9444 12940
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 11606 12928 11612 12980
rect 11664 12968 11670 12980
rect 11793 12971 11851 12977
rect 11793 12968 11805 12971
rect 11664 12940 11805 12968
rect 11664 12928 11670 12940
rect 11793 12937 11805 12940
rect 11839 12937 11851 12971
rect 11793 12931 11851 12937
rect 12434 12928 12440 12980
rect 12492 12928 12498 12980
rect 13541 12971 13599 12977
rect 13541 12937 13553 12971
rect 13587 12968 13599 12971
rect 15378 12968 15384 12980
rect 13587 12940 15384 12968
rect 13587 12937 13599 12940
rect 13541 12931 13599 12937
rect 15378 12928 15384 12940
rect 15436 12928 15442 12980
rect 15657 12971 15715 12977
rect 15657 12937 15669 12971
rect 15703 12968 15715 12971
rect 16022 12968 16028 12980
rect 15703 12940 16028 12968
rect 15703 12937 15715 12940
rect 15657 12931 15715 12937
rect 16022 12928 16028 12940
rect 16080 12928 16086 12980
rect 19426 12928 19432 12980
rect 19484 12968 19490 12980
rect 20073 12971 20131 12977
rect 20073 12968 20085 12971
rect 19484 12940 20085 12968
rect 19484 12928 19490 12940
rect 20073 12937 20085 12940
rect 20119 12937 20131 12971
rect 20073 12931 20131 12937
rect 20257 12971 20315 12977
rect 20257 12937 20269 12971
rect 20303 12968 20315 12971
rect 20530 12968 20536 12980
rect 20303 12940 20536 12968
rect 20303 12937 20315 12940
rect 20257 12931 20315 12937
rect 9323 12872 9444 12900
rect 9493 12903 9551 12909
rect 9323 12869 9335 12872
rect 9277 12863 9335 12869
rect 9493 12869 9505 12903
rect 9539 12900 9551 12903
rect 9539 12872 9628 12900
rect 9539 12869 9551 12872
rect 9493 12863 9551 12869
rect 5537 12835 5595 12841
rect 5537 12832 5549 12835
rect 4856 12804 5549 12832
rect 4856 12792 4862 12804
rect 5537 12801 5549 12804
rect 5583 12801 5595 12835
rect 5537 12795 5595 12801
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12801 5871 12835
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 5813 12795 5871 12801
rect 5920 12804 6561 12832
rect 2222 12724 2228 12776
rect 2280 12764 2286 12776
rect 2409 12767 2467 12773
rect 2409 12764 2421 12767
rect 2280 12736 2421 12764
rect 2280 12724 2286 12736
rect 2409 12733 2421 12736
rect 2455 12733 2467 12767
rect 2409 12727 2467 12733
rect 5552 12696 5580 12795
rect 5920 12696 5948 12804
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 6825 12835 6883 12841
rect 6825 12801 6837 12835
rect 6871 12832 6883 12835
rect 7006 12832 7012 12844
rect 6871 12804 7012 12832
rect 6871 12801 6883 12804
rect 6825 12795 6883 12801
rect 7006 12792 7012 12804
rect 7064 12792 7070 12844
rect 7098 12792 7104 12844
rect 7156 12832 7162 12844
rect 7469 12835 7527 12841
rect 7469 12832 7481 12835
rect 7156 12804 7481 12832
rect 7156 12792 7162 12804
rect 7469 12801 7481 12804
rect 7515 12801 7527 12835
rect 7469 12795 7527 12801
rect 8386 12792 8392 12844
rect 8444 12792 8450 12844
rect 9600 12776 9628 12872
rect 13464 12872 15240 12900
rect 10318 12792 10324 12844
rect 10376 12792 10382 12844
rect 10410 12792 10416 12844
rect 10468 12832 10474 12844
rect 10505 12835 10563 12841
rect 10505 12832 10517 12835
rect 10468 12804 10517 12832
rect 10468 12792 10474 12804
rect 10505 12801 10517 12804
rect 10551 12801 10563 12835
rect 10505 12795 10563 12801
rect 10870 12792 10876 12844
rect 10928 12792 10934 12844
rect 10962 12792 10968 12844
rect 11020 12792 11026 12844
rect 11146 12792 11152 12844
rect 11204 12792 11210 12844
rect 11606 12792 11612 12844
rect 11664 12832 11670 12844
rect 11701 12835 11759 12841
rect 11701 12832 11713 12835
rect 11664 12804 11713 12832
rect 11664 12792 11670 12804
rect 11701 12801 11713 12804
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 12342 12792 12348 12844
rect 12400 12792 12406 12844
rect 12618 12792 12624 12844
rect 12676 12832 12682 12844
rect 13464 12841 13492 12872
rect 13449 12835 13507 12841
rect 13449 12832 13461 12835
rect 12676 12804 13461 12832
rect 12676 12792 12682 12804
rect 13449 12801 13461 12804
rect 13495 12801 13507 12835
rect 13449 12795 13507 12801
rect 13633 12835 13691 12841
rect 13633 12801 13645 12835
rect 13679 12832 13691 12835
rect 15102 12832 15108 12844
rect 13679 12804 15108 12832
rect 13679 12801 13691 12804
rect 13633 12795 13691 12801
rect 15102 12792 15108 12804
rect 15160 12792 15166 12844
rect 15212 12832 15240 12872
rect 16758 12860 16764 12912
rect 16816 12900 16822 12912
rect 16853 12903 16911 12909
rect 16853 12900 16865 12903
rect 16816 12872 16865 12900
rect 16816 12860 16822 12872
rect 16853 12869 16865 12872
rect 16899 12900 16911 12903
rect 16942 12900 16948 12912
rect 16899 12872 16948 12900
rect 16899 12869 16911 12872
rect 16853 12863 16911 12869
rect 16942 12860 16948 12872
rect 17000 12860 17006 12912
rect 19518 12900 19524 12912
rect 18156 12872 19524 12900
rect 15212 12804 15332 12832
rect 7285 12767 7343 12773
rect 7285 12764 7297 12767
rect 5552 12668 5948 12696
rect 6104 12736 7297 12764
rect 3234 12588 3240 12640
rect 3292 12628 3298 12640
rect 3421 12631 3479 12637
rect 3421 12628 3433 12631
rect 3292 12600 3433 12628
rect 3292 12588 3298 12600
rect 3421 12597 3433 12600
rect 3467 12597 3479 12631
rect 3421 12591 3479 12597
rect 4614 12588 4620 12640
rect 4672 12588 4678 12640
rect 5537 12631 5595 12637
rect 5537 12597 5549 12631
rect 5583 12628 5595 12631
rect 5626 12628 5632 12640
rect 5583 12600 5632 12628
rect 5583 12597 5595 12600
rect 5537 12591 5595 12597
rect 5626 12588 5632 12600
rect 5684 12588 5690 12640
rect 5718 12588 5724 12640
rect 5776 12628 5782 12640
rect 6104 12628 6132 12736
rect 7285 12733 7297 12736
rect 7331 12733 7343 12767
rect 7285 12727 7343 12733
rect 8662 12724 8668 12776
rect 8720 12764 8726 12776
rect 9582 12764 9588 12776
rect 8720 12736 9588 12764
rect 8720 12724 8726 12736
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 15304 12773 15332 12804
rect 15470 12792 15476 12844
rect 15528 12792 15534 12844
rect 17034 12792 17040 12844
rect 17092 12792 17098 12844
rect 17862 12792 17868 12844
rect 17920 12832 17926 12844
rect 18156 12841 18184 12872
rect 19518 12860 19524 12872
rect 19576 12860 19582 12912
rect 20088 12900 20116 12931
rect 20530 12928 20536 12940
rect 20588 12928 20594 12980
rect 20346 12900 20352 12912
rect 20088 12872 20352 12900
rect 20346 12860 20352 12872
rect 20404 12860 20410 12912
rect 18141 12835 18199 12841
rect 18141 12832 18153 12835
rect 17920 12804 18153 12832
rect 17920 12792 17926 12804
rect 18141 12801 18153 12804
rect 18187 12801 18199 12835
rect 18141 12795 18199 12801
rect 18230 12792 18236 12844
rect 18288 12792 18294 12844
rect 18322 12792 18328 12844
rect 18380 12792 18386 12844
rect 18509 12835 18567 12841
rect 18509 12801 18521 12835
rect 18555 12801 18567 12835
rect 18509 12795 18567 12801
rect 13265 12767 13323 12773
rect 13265 12733 13277 12767
rect 13311 12764 13323 12767
rect 15197 12767 15255 12773
rect 15197 12764 15209 12767
rect 13311 12736 15209 12764
rect 13311 12733 13323 12736
rect 13265 12727 13323 12733
rect 6733 12699 6791 12705
rect 6733 12665 6745 12699
rect 6779 12696 6791 12699
rect 7742 12696 7748 12708
rect 6779 12668 7748 12696
rect 6779 12665 6791 12668
rect 6733 12659 6791 12665
rect 7742 12656 7748 12668
rect 7800 12696 7806 12708
rect 8573 12699 8631 12705
rect 8573 12696 8585 12699
rect 7800 12668 8585 12696
rect 7800 12656 7806 12668
rect 8573 12665 8585 12668
rect 8619 12665 8631 12699
rect 8573 12659 8631 12665
rect 5776 12600 6132 12628
rect 6825 12631 6883 12637
rect 5776 12588 5782 12600
rect 6825 12597 6837 12631
rect 6871 12628 6883 12631
rect 7190 12628 7196 12640
rect 6871 12600 7196 12628
rect 6871 12597 6883 12600
rect 6825 12591 6883 12597
rect 7190 12588 7196 12600
rect 7248 12588 7254 12640
rect 7653 12631 7711 12637
rect 7653 12597 7665 12631
rect 7699 12628 7711 12631
rect 7926 12628 7932 12640
rect 7699 12600 7932 12628
rect 7699 12597 7711 12600
rect 7653 12591 7711 12597
rect 7926 12588 7932 12600
rect 7984 12588 7990 12640
rect 8202 12588 8208 12640
rect 8260 12588 8266 12640
rect 8938 12588 8944 12640
rect 8996 12628 9002 12640
rect 9309 12631 9367 12637
rect 9309 12628 9321 12631
rect 8996 12600 9321 12628
rect 8996 12588 9002 12600
rect 9309 12597 9321 12600
rect 9355 12597 9367 12631
rect 9309 12591 9367 12597
rect 13722 12588 13728 12640
rect 13780 12628 13786 12640
rect 13817 12631 13875 12637
rect 13817 12628 13829 12631
rect 13780 12600 13829 12628
rect 13780 12588 13786 12600
rect 13817 12597 13829 12600
rect 13863 12597 13875 12631
rect 15120 12628 15148 12736
rect 15197 12733 15209 12736
rect 15243 12733 15255 12767
rect 15197 12727 15255 12733
rect 15289 12767 15347 12773
rect 15289 12733 15301 12767
rect 15335 12733 15347 12767
rect 15289 12727 15347 12733
rect 15378 12724 15384 12776
rect 15436 12764 15442 12776
rect 15838 12764 15844 12776
rect 15436 12736 15844 12764
rect 15436 12724 15442 12736
rect 15838 12724 15844 12736
rect 15896 12724 15902 12776
rect 18524 12764 18552 12795
rect 19334 12792 19340 12844
rect 19392 12792 19398 12844
rect 19426 12792 19432 12844
rect 19484 12792 19490 12844
rect 20198 12835 20256 12841
rect 20198 12832 20210 12835
rect 19536 12804 20210 12832
rect 18598 12764 18604 12776
rect 17236 12736 18604 12764
rect 17236 12640 17264 12736
rect 18598 12724 18604 12736
rect 18656 12724 18662 12776
rect 17678 12656 17684 12708
rect 17736 12696 17742 12708
rect 19536 12696 19564 12804
rect 20198 12801 20210 12804
rect 20244 12801 20256 12835
rect 20198 12795 20256 12801
rect 20622 12792 20628 12844
rect 20680 12792 20686 12844
rect 22186 12792 22192 12844
rect 22244 12792 22250 12844
rect 19613 12767 19671 12773
rect 19613 12733 19625 12767
rect 19659 12764 19671 12767
rect 20438 12764 20444 12776
rect 19659 12736 20444 12764
rect 19659 12733 19671 12736
rect 19613 12727 19671 12733
rect 20438 12724 20444 12736
rect 20496 12724 20502 12776
rect 20717 12767 20775 12773
rect 20717 12733 20729 12767
rect 20763 12764 20775 12767
rect 21726 12764 21732 12776
rect 20763 12736 21732 12764
rect 20763 12733 20775 12736
rect 20717 12727 20775 12733
rect 21726 12724 21732 12736
rect 21784 12764 21790 12776
rect 22097 12767 22155 12773
rect 22097 12764 22109 12767
rect 21784 12736 22109 12764
rect 21784 12724 21790 12736
rect 22097 12733 22109 12736
rect 22143 12733 22155 12767
rect 22097 12727 22155 12733
rect 17736 12668 19564 12696
rect 17736 12656 17742 12668
rect 16022 12628 16028 12640
rect 15120 12600 16028 12628
rect 13817 12591 13875 12597
rect 16022 12588 16028 12600
rect 16080 12588 16086 12640
rect 17129 12631 17187 12637
rect 17129 12597 17141 12631
rect 17175 12628 17187 12631
rect 17218 12628 17224 12640
rect 17175 12600 17224 12628
rect 17175 12597 17187 12600
rect 17129 12591 17187 12597
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 17865 12631 17923 12637
rect 17865 12597 17877 12631
rect 17911 12628 17923 12631
rect 18138 12628 18144 12640
rect 17911 12600 18144 12628
rect 17911 12597 17923 12600
rect 17865 12591 17923 12597
rect 18138 12588 18144 12600
rect 18196 12588 18202 12640
rect 19518 12588 19524 12640
rect 19576 12588 19582 12640
rect 1104 12538 22816 12560
rect 1104 12486 3664 12538
rect 3716 12486 3728 12538
rect 3780 12486 3792 12538
rect 3844 12486 3856 12538
rect 3908 12486 3920 12538
rect 3972 12486 9092 12538
rect 9144 12486 9156 12538
rect 9208 12486 9220 12538
rect 9272 12486 9284 12538
rect 9336 12486 9348 12538
rect 9400 12486 14520 12538
rect 14572 12486 14584 12538
rect 14636 12486 14648 12538
rect 14700 12486 14712 12538
rect 14764 12486 14776 12538
rect 14828 12486 19948 12538
rect 20000 12486 20012 12538
rect 20064 12486 20076 12538
rect 20128 12486 20140 12538
rect 20192 12486 20204 12538
rect 20256 12486 22816 12538
rect 1104 12464 22816 12486
rect 3142 12384 3148 12436
rect 3200 12384 3206 12436
rect 7006 12384 7012 12436
rect 7064 12384 7070 12436
rect 7742 12384 7748 12436
rect 7800 12384 7806 12436
rect 10686 12384 10692 12436
rect 10744 12424 10750 12436
rect 10965 12427 11023 12433
rect 10965 12424 10977 12427
rect 10744 12396 10977 12424
rect 10744 12384 10750 12396
rect 10965 12393 10977 12396
rect 11011 12393 11023 12427
rect 10965 12387 11023 12393
rect 13078 12384 13084 12436
rect 13136 12384 13142 12436
rect 13170 12384 13176 12436
rect 13228 12424 13234 12436
rect 13538 12424 13544 12436
rect 13228 12396 13544 12424
rect 13228 12384 13234 12396
rect 13538 12384 13544 12396
rect 13596 12384 13602 12436
rect 13630 12384 13636 12436
rect 13688 12424 13694 12436
rect 17862 12424 17868 12436
rect 13688 12396 17868 12424
rect 13688 12384 13694 12396
rect 17862 12384 17868 12396
rect 17920 12384 17926 12436
rect 18598 12384 18604 12436
rect 18656 12424 18662 12436
rect 21082 12424 21088 12436
rect 18656 12396 21088 12424
rect 18656 12384 18662 12396
rect 21082 12384 21088 12396
rect 21140 12384 21146 12436
rect 2866 12316 2872 12368
rect 2924 12356 2930 12368
rect 5813 12359 5871 12365
rect 5813 12356 5825 12359
rect 2924 12328 4016 12356
rect 2924 12316 2930 12328
rect 2317 12291 2375 12297
rect 2317 12257 2329 12291
rect 2363 12288 2375 12291
rect 2774 12288 2780 12300
rect 2363 12260 2780 12288
rect 2363 12257 2375 12260
rect 2317 12251 2375 12257
rect 2774 12248 2780 12260
rect 2832 12288 2838 12300
rect 3988 12297 4016 12328
rect 4724 12328 5825 12356
rect 4724 12300 4752 12328
rect 5813 12325 5825 12328
rect 5859 12356 5871 12359
rect 5859 12328 6040 12356
rect 5859 12325 5871 12328
rect 5813 12319 5871 12325
rect 3973 12291 4031 12297
rect 2832 12260 2912 12288
rect 2832 12248 2838 12260
rect 2130 12180 2136 12232
rect 2188 12180 2194 12232
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12220 2467 12223
rect 2498 12220 2504 12232
rect 2455 12192 2504 12220
rect 2455 12189 2467 12192
rect 2409 12183 2467 12189
rect 2498 12180 2504 12192
rect 2556 12180 2562 12232
rect 2884 12229 2912 12260
rect 3973 12257 3985 12291
rect 4019 12257 4031 12291
rect 3973 12251 4031 12257
rect 4706 12248 4712 12300
rect 4764 12248 4770 12300
rect 5718 12248 5724 12300
rect 5776 12288 5782 12300
rect 5905 12291 5963 12297
rect 5905 12288 5917 12291
rect 5776 12260 5917 12288
rect 5776 12248 5782 12260
rect 5905 12257 5917 12260
rect 5951 12257 5963 12291
rect 5905 12251 5963 12257
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12220 2927 12223
rect 3418 12220 3424 12232
rect 2915 12192 3424 12220
rect 2915 12189 2927 12192
rect 2869 12183 2927 12189
rect 3418 12180 3424 12192
rect 3476 12220 3482 12232
rect 3476 12192 4384 12220
rect 3476 12180 3482 12192
rect 2516 12152 2544 12180
rect 2961 12155 3019 12161
rect 2961 12152 2973 12155
rect 2516 12124 2973 12152
rect 2884 12096 2912 12124
rect 2961 12121 2973 12124
rect 3007 12121 3019 12155
rect 2961 12115 3019 12121
rect 3142 12112 3148 12164
rect 3200 12112 3206 12164
rect 4356 12161 4384 12192
rect 5626 12180 5632 12232
rect 5684 12180 5690 12232
rect 4341 12155 4399 12161
rect 4341 12121 4353 12155
rect 4387 12121 4399 12155
rect 4341 12115 4399 12121
rect 1946 12044 1952 12096
rect 2004 12044 2010 12096
rect 2866 12044 2872 12096
rect 2924 12044 2930 12096
rect 3160 12084 3188 12112
rect 4157 12087 4215 12093
rect 4157 12084 4169 12087
rect 3160 12056 4169 12084
rect 4157 12053 4169 12056
rect 4203 12053 4215 12087
rect 4157 12047 4215 12053
rect 4246 12044 4252 12096
rect 4304 12044 4310 12096
rect 5350 12044 5356 12096
rect 5408 12084 5414 12096
rect 5445 12087 5503 12093
rect 5445 12084 5457 12087
rect 5408 12056 5457 12084
rect 5408 12044 5414 12056
rect 5445 12053 5457 12056
rect 5491 12053 5503 12087
rect 5920 12084 5948 12251
rect 6012 12220 6040 12328
rect 9858 12316 9864 12368
rect 9916 12356 9922 12368
rect 11425 12359 11483 12365
rect 11425 12356 11437 12359
rect 9916 12328 11437 12356
rect 9916 12316 9922 12328
rect 11425 12325 11437 12328
rect 11471 12325 11483 12359
rect 11425 12319 11483 12325
rect 11514 12316 11520 12368
rect 11572 12356 11578 12368
rect 11572 12328 13860 12356
rect 11572 12316 11578 12328
rect 8113 12291 8171 12297
rect 8113 12288 8125 12291
rect 6886 12260 8125 12288
rect 6733 12223 6791 12229
rect 6733 12220 6745 12223
rect 6012 12192 6745 12220
rect 6733 12189 6745 12192
rect 6779 12220 6791 12223
rect 6886 12220 6914 12260
rect 8113 12257 8125 12260
rect 8159 12288 8171 12291
rect 8938 12288 8944 12300
rect 8159 12260 8944 12288
rect 8159 12257 8171 12260
rect 8113 12251 8171 12257
rect 8938 12248 8944 12260
rect 8996 12248 9002 12300
rect 10318 12248 10324 12300
rect 10376 12248 10382 12300
rect 11146 12288 11152 12300
rect 10704 12260 11152 12288
rect 6779 12192 6914 12220
rect 6779 12189 6791 12192
rect 6733 12183 6791 12189
rect 7926 12180 7932 12232
rect 7984 12180 7990 12232
rect 7009 12155 7067 12161
rect 7009 12121 7021 12155
rect 7055 12152 7067 12155
rect 7098 12152 7104 12164
rect 7055 12124 7104 12152
rect 7055 12121 7067 12124
rect 7009 12115 7067 12121
rect 7098 12112 7104 12124
rect 7156 12112 7162 12164
rect 8956 12152 8984 12248
rect 9582 12180 9588 12232
rect 9640 12220 9646 12232
rect 10704 12229 10732 12260
rect 11146 12248 11152 12260
rect 11204 12248 11210 12300
rect 12084 12297 12112 12328
rect 12069 12291 12127 12297
rect 12069 12257 12081 12291
rect 12115 12257 12127 12291
rect 12069 12251 12127 12257
rect 13265 12291 13323 12297
rect 13265 12257 13277 12291
rect 13311 12288 13323 12291
rect 13722 12288 13728 12300
rect 13311 12260 13728 12288
rect 13311 12257 13323 12260
rect 13265 12251 13323 12257
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 10689 12223 10747 12229
rect 10689 12220 10701 12223
rect 9640 12192 10701 12220
rect 9640 12180 9646 12192
rect 10689 12189 10701 12192
rect 10735 12189 10747 12223
rect 10689 12183 10747 12189
rect 10781 12223 10839 12229
rect 10781 12189 10793 12223
rect 10827 12220 10839 12223
rect 10870 12220 10876 12232
rect 10827 12192 10876 12220
rect 10827 12189 10839 12192
rect 10781 12183 10839 12189
rect 10870 12180 10876 12192
rect 10928 12220 10934 12232
rect 11793 12223 11851 12229
rect 11793 12220 11805 12223
rect 10928 12192 11805 12220
rect 10928 12180 10934 12192
rect 11793 12189 11805 12192
rect 11839 12189 11851 12223
rect 11793 12183 11851 12189
rect 13354 12180 13360 12232
rect 13412 12180 13418 12232
rect 13446 12180 13452 12232
rect 13504 12180 13510 12232
rect 13541 12223 13599 12229
rect 13541 12189 13553 12223
rect 13587 12220 13599 12223
rect 13832 12220 13860 12328
rect 15304 12328 15608 12356
rect 15304 12297 15332 12328
rect 15289 12291 15347 12297
rect 15289 12257 15301 12291
rect 15335 12257 15347 12291
rect 15580 12288 15608 12328
rect 16758 12316 16764 12368
rect 16816 12356 16822 12368
rect 17129 12359 17187 12365
rect 17129 12356 17141 12359
rect 16816 12328 17141 12356
rect 16816 12316 16822 12328
rect 17129 12325 17141 12328
rect 17175 12356 17187 12359
rect 19702 12356 19708 12368
rect 17175 12328 19708 12356
rect 17175 12325 17187 12328
rect 17129 12319 17187 12325
rect 19702 12316 19708 12328
rect 19760 12316 19766 12368
rect 19794 12316 19800 12368
rect 19852 12356 19858 12368
rect 20714 12356 20720 12368
rect 19852 12328 20720 12356
rect 19852 12316 19858 12328
rect 20714 12316 20720 12328
rect 20772 12316 20778 12368
rect 16850 12288 16856 12300
rect 15580 12260 16856 12288
rect 15289 12251 15347 12257
rect 16850 12248 16856 12260
rect 16908 12248 16914 12300
rect 20162 12288 20168 12300
rect 17880 12260 20168 12288
rect 13906 12220 13912 12232
rect 13587 12192 13912 12220
rect 13587 12189 13599 12192
rect 13541 12183 13599 12189
rect 13906 12180 13912 12192
rect 13964 12180 13970 12232
rect 14918 12180 14924 12232
rect 14976 12220 14982 12232
rect 15013 12223 15071 12229
rect 15013 12220 15025 12223
rect 14976 12192 15025 12220
rect 14976 12180 14982 12192
rect 15013 12189 15025 12192
rect 15059 12189 15071 12223
rect 15013 12183 15071 12189
rect 15197 12223 15255 12229
rect 15197 12189 15209 12223
rect 15243 12189 15255 12223
rect 15197 12183 15255 12189
rect 10410 12152 10416 12164
rect 8956 12124 10416 12152
rect 10410 12112 10416 12124
rect 10468 12112 10474 12164
rect 13372 12152 13400 12180
rect 15212 12152 15240 12183
rect 15378 12180 15384 12232
rect 15436 12180 15442 12232
rect 15565 12223 15623 12229
rect 15565 12189 15577 12223
rect 15611 12220 15623 12223
rect 16393 12223 16451 12229
rect 16393 12220 16405 12223
rect 15611 12192 16405 12220
rect 15611 12189 15623 12192
rect 15565 12183 15623 12189
rect 16393 12189 16405 12192
rect 16439 12220 16451 12223
rect 16482 12220 16488 12232
rect 16439 12192 16488 12220
rect 16439 12189 16451 12192
rect 16393 12183 16451 12189
rect 16482 12180 16488 12192
rect 16540 12180 16546 12232
rect 16574 12180 16580 12232
rect 16632 12180 16638 12232
rect 16666 12180 16672 12232
rect 16724 12220 16730 12232
rect 17218 12220 17224 12232
rect 16724 12192 17224 12220
rect 16724 12180 16730 12192
rect 17218 12180 17224 12192
rect 17276 12180 17282 12232
rect 17310 12180 17316 12232
rect 17368 12220 17374 12232
rect 17678 12220 17684 12232
rect 17368 12192 17684 12220
rect 17368 12180 17374 12192
rect 17678 12180 17684 12192
rect 17736 12180 17742 12232
rect 17880 12229 17908 12260
rect 20162 12248 20168 12260
rect 20220 12248 20226 12300
rect 20438 12248 20444 12300
rect 20496 12288 20502 12300
rect 20990 12288 20996 12300
rect 20496 12260 20996 12288
rect 20496 12248 20502 12260
rect 20990 12248 20996 12260
rect 21048 12248 21054 12300
rect 17865 12223 17923 12229
rect 17865 12189 17877 12223
rect 17911 12189 17923 12223
rect 17865 12183 17923 12189
rect 19334 12180 19340 12232
rect 19392 12220 19398 12232
rect 20257 12223 20315 12229
rect 20257 12220 20269 12223
rect 19392 12192 20269 12220
rect 19392 12180 19398 12192
rect 20257 12189 20269 12192
rect 20303 12189 20315 12223
rect 20257 12183 20315 12189
rect 20346 12180 20352 12232
rect 20404 12180 20410 12232
rect 20533 12223 20591 12229
rect 20533 12189 20545 12223
rect 20579 12220 20591 12223
rect 20714 12220 20720 12232
rect 20579 12192 20720 12220
rect 20579 12189 20591 12192
rect 20533 12183 20591 12189
rect 20714 12180 20720 12192
rect 20772 12180 20778 12232
rect 20806 12180 20812 12232
rect 20864 12220 20870 12232
rect 21545 12223 21603 12229
rect 21545 12220 21557 12223
rect 20864 12192 21557 12220
rect 20864 12180 20870 12192
rect 21545 12189 21557 12192
rect 21591 12189 21603 12223
rect 21545 12183 21603 12189
rect 21726 12180 21732 12232
rect 21784 12180 21790 12232
rect 21637 12155 21695 12161
rect 13372 12124 13584 12152
rect 15212 12124 20208 12152
rect 13556 12096 13584 12124
rect 6270 12084 6276 12096
rect 5920 12056 6276 12084
rect 5445 12047 5503 12053
rect 6270 12044 6276 12056
rect 6328 12084 6334 12096
rect 6825 12087 6883 12093
rect 6825 12084 6837 12087
rect 6328 12056 6837 12084
rect 6328 12044 6334 12056
rect 6825 12053 6837 12056
rect 6871 12053 6883 12087
rect 6825 12047 6883 12053
rect 8478 12044 8484 12096
rect 8536 12084 8542 12096
rect 8754 12084 8760 12096
rect 8536 12056 8760 12084
rect 8536 12044 8542 12056
rect 8754 12044 8760 12056
rect 8812 12084 8818 12096
rect 10505 12087 10563 12093
rect 10505 12084 10517 12087
rect 8812 12056 10517 12084
rect 8812 12044 8818 12056
rect 10505 12053 10517 12056
rect 10551 12084 10563 12087
rect 11606 12084 11612 12096
rect 10551 12056 11612 12084
rect 10551 12053 10563 12056
rect 10505 12047 10563 12053
rect 11606 12044 11612 12056
rect 11664 12044 11670 12096
rect 11698 12044 11704 12096
rect 11756 12084 11762 12096
rect 11885 12087 11943 12093
rect 11885 12084 11897 12087
rect 11756 12056 11897 12084
rect 11756 12044 11762 12056
rect 11885 12053 11897 12056
rect 11931 12084 11943 12087
rect 12342 12084 12348 12096
rect 11931 12056 12348 12084
rect 11931 12053 11943 12056
rect 11885 12047 11943 12053
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 13538 12044 13544 12096
rect 13596 12044 13602 12096
rect 15746 12044 15752 12096
rect 15804 12044 15810 12096
rect 16485 12087 16543 12093
rect 16485 12053 16497 12087
rect 16531 12084 16543 12087
rect 17678 12084 17684 12096
rect 16531 12056 17684 12084
rect 16531 12053 16543 12056
rect 16485 12047 16543 12053
rect 17678 12044 17684 12056
rect 17736 12044 17742 12096
rect 17773 12087 17831 12093
rect 17773 12053 17785 12087
rect 17819 12084 17831 12087
rect 18690 12084 18696 12096
rect 17819 12056 18696 12084
rect 17819 12053 17831 12056
rect 17773 12047 17831 12053
rect 18690 12044 18696 12056
rect 18748 12044 18754 12096
rect 20070 12044 20076 12096
rect 20128 12044 20134 12096
rect 20180 12084 20208 12124
rect 21637 12121 21649 12155
rect 21683 12121 21695 12155
rect 21637 12115 21695 12121
rect 21266 12084 21272 12096
rect 20180 12056 21272 12084
rect 21266 12044 21272 12056
rect 21324 12084 21330 12096
rect 21652 12084 21680 12115
rect 21324 12056 21680 12084
rect 21324 12044 21330 12056
rect 1104 11994 22976 12016
rect 1104 11942 6378 11994
rect 6430 11942 6442 11994
rect 6494 11942 6506 11994
rect 6558 11942 6570 11994
rect 6622 11942 6634 11994
rect 6686 11942 11806 11994
rect 11858 11942 11870 11994
rect 11922 11942 11934 11994
rect 11986 11942 11998 11994
rect 12050 11942 12062 11994
rect 12114 11942 17234 11994
rect 17286 11942 17298 11994
rect 17350 11942 17362 11994
rect 17414 11942 17426 11994
rect 17478 11942 17490 11994
rect 17542 11942 22662 11994
rect 22714 11942 22726 11994
rect 22778 11942 22790 11994
rect 22842 11942 22854 11994
rect 22906 11942 22918 11994
rect 22970 11942 22976 11994
rect 1104 11920 22976 11942
rect 15378 11840 15384 11892
rect 15436 11880 15442 11892
rect 16574 11880 16580 11892
rect 15436 11852 16580 11880
rect 15436 11840 15442 11852
rect 16574 11840 16580 11852
rect 16632 11840 16638 11892
rect 17494 11840 17500 11892
rect 17552 11880 17558 11892
rect 17770 11880 17776 11892
rect 17552 11852 17776 11880
rect 17552 11840 17558 11852
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 20806 11880 20812 11892
rect 17972 11852 20812 11880
rect 2317 11815 2375 11821
rect 2317 11781 2329 11815
rect 2363 11812 2375 11815
rect 2498 11812 2504 11824
rect 2363 11784 2504 11812
rect 2363 11781 2375 11784
rect 2317 11775 2375 11781
rect 2498 11772 2504 11784
rect 2556 11772 2562 11824
rect 2133 11747 2191 11753
rect 2133 11713 2145 11747
rect 2179 11744 2191 11747
rect 2222 11744 2228 11756
rect 2179 11716 2228 11744
rect 2179 11713 2191 11716
rect 2133 11707 2191 11713
rect 2222 11704 2228 11716
rect 2280 11704 2286 11756
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11744 2467 11747
rect 2774 11744 2780 11756
rect 2455 11716 2780 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 2774 11704 2780 11716
rect 2832 11704 2838 11756
rect 4154 11704 4160 11756
rect 4212 11744 4218 11756
rect 4433 11747 4491 11753
rect 4433 11744 4445 11747
rect 4212 11716 4445 11744
rect 4212 11704 4218 11716
rect 4433 11713 4445 11716
rect 4479 11713 4491 11747
rect 4433 11707 4491 11713
rect 4614 11704 4620 11756
rect 4672 11704 4678 11756
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11744 15623 11747
rect 16758 11744 16764 11756
rect 15611 11716 16764 11744
rect 15611 11713 15623 11716
rect 15565 11707 15623 11713
rect 16758 11704 16764 11716
rect 16816 11704 16822 11756
rect 16850 11704 16856 11756
rect 16908 11744 16914 11756
rect 17129 11747 17187 11753
rect 17129 11744 17141 11747
rect 16908 11716 17141 11744
rect 16908 11704 16914 11716
rect 17129 11713 17141 11716
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 17222 11747 17280 11753
rect 17222 11713 17234 11747
rect 17268 11713 17280 11747
rect 17222 11707 17280 11713
rect 4338 11636 4344 11688
rect 4396 11636 4402 11688
rect 15381 11679 15439 11685
rect 15381 11645 15393 11679
rect 15427 11645 15439 11679
rect 15381 11639 15439 11645
rect 2130 11568 2136 11620
rect 2188 11568 2194 11620
rect 4798 11500 4804 11552
rect 4856 11500 4862 11552
rect 14918 11500 14924 11552
rect 14976 11540 14982 11552
rect 15396 11540 15424 11639
rect 16482 11636 16488 11688
rect 16540 11676 16546 11688
rect 17236 11676 17264 11707
rect 17402 11704 17408 11756
rect 17460 11704 17466 11756
rect 17678 11753 17684 11756
rect 17497 11747 17555 11753
rect 17497 11713 17509 11747
rect 17543 11713 17555 11747
rect 17497 11707 17555 11713
rect 17635 11747 17684 11753
rect 17635 11713 17647 11747
rect 17681 11713 17684 11747
rect 17635 11707 17684 11713
rect 16540 11648 17264 11676
rect 17512 11676 17540 11707
rect 17678 11704 17684 11707
rect 17736 11704 17742 11756
rect 17972 11676 18000 11852
rect 20806 11840 20812 11852
rect 20864 11840 20870 11892
rect 19518 11772 19524 11824
rect 19576 11812 19582 11824
rect 19981 11815 20039 11821
rect 19981 11812 19993 11815
rect 19576 11784 19993 11812
rect 19576 11772 19582 11784
rect 19981 11781 19993 11784
rect 20027 11781 20039 11815
rect 19981 11775 20039 11781
rect 20070 11772 20076 11824
rect 20128 11772 20134 11824
rect 19705 11747 19763 11753
rect 19705 11744 19717 11747
rect 19536 11716 19717 11744
rect 19536 11688 19564 11716
rect 19705 11713 19717 11716
rect 19751 11713 19763 11747
rect 19705 11707 19763 11713
rect 20990 11704 20996 11756
rect 21048 11744 21054 11756
rect 21177 11747 21235 11753
rect 21177 11744 21189 11747
rect 21048 11716 21189 11744
rect 21048 11704 21054 11716
rect 21177 11713 21189 11716
rect 21223 11713 21235 11747
rect 21177 11707 21235 11713
rect 21361 11747 21419 11753
rect 21361 11713 21373 11747
rect 21407 11713 21419 11747
rect 21361 11707 21419 11713
rect 17512 11648 18000 11676
rect 16540 11636 16546 11648
rect 15930 11568 15936 11620
rect 15988 11608 15994 11620
rect 17512 11608 17540 11648
rect 19518 11636 19524 11688
rect 19576 11636 19582 11688
rect 19613 11679 19671 11685
rect 19613 11645 19625 11679
rect 19659 11645 19671 11679
rect 19613 11639 19671 11645
rect 18230 11608 18236 11620
rect 15988 11580 17540 11608
rect 17696 11580 18236 11608
rect 15988 11568 15994 11580
rect 17696 11540 17724 11580
rect 18230 11568 18236 11580
rect 18288 11568 18294 11620
rect 19334 11568 19340 11620
rect 19392 11608 19398 11620
rect 19628 11608 19656 11639
rect 20714 11636 20720 11688
rect 20772 11676 20778 11688
rect 21376 11676 21404 11707
rect 20772 11648 21404 11676
rect 20772 11636 20778 11648
rect 19392 11580 19656 11608
rect 19392 11568 19398 11580
rect 14976 11512 17724 11540
rect 17773 11543 17831 11549
rect 14976 11500 14982 11512
rect 17773 11509 17785 11543
rect 17819 11540 17831 11543
rect 17862 11540 17868 11552
rect 17819 11512 17868 11540
rect 17819 11509 17831 11512
rect 17773 11503 17831 11509
rect 17862 11500 17868 11512
rect 17920 11500 17926 11552
rect 19429 11543 19487 11549
rect 19429 11509 19441 11543
rect 19475 11540 19487 11543
rect 19610 11540 19616 11552
rect 19475 11512 19616 11540
rect 19475 11509 19487 11512
rect 19429 11503 19487 11509
rect 19610 11500 19616 11512
rect 19668 11500 19674 11552
rect 21174 11500 21180 11552
rect 21232 11500 21238 11552
rect 1104 11450 22816 11472
rect 1104 11398 3664 11450
rect 3716 11398 3728 11450
rect 3780 11398 3792 11450
rect 3844 11398 3856 11450
rect 3908 11398 3920 11450
rect 3972 11398 9092 11450
rect 9144 11398 9156 11450
rect 9208 11398 9220 11450
rect 9272 11398 9284 11450
rect 9336 11398 9348 11450
rect 9400 11398 14520 11450
rect 14572 11398 14584 11450
rect 14636 11398 14648 11450
rect 14700 11398 14712 11450
rect 14764 11398 14776 11450
rect 14828 11398 19948 11450
rect 20000 11398 20012 11450
rect 20064 11398 20076 11450
rect 20128 11398 20140 11450
rect 20192 11398 20204 11450
rect 20256 11398 22816 11450
rect 1104 11376 22816 11398
rect 6270 11296 6276 11348
rect 6328 11336 6334 11348
rect 6457 11339 6515 11345
rect 6457 11336 6469 11339
rect 6328 11308 6469 11336
rect 6328 11296 6334 11308
rect 6457 11305 6469 11308
rect 6503 11305 6515 11339
rect 6457 11299 6515 11305
rect 7098 11296 7104 11348
rect 7156 11336 7162 11348
rect 8297 11339 8355 11345
rect 8297 11336 8309 11339
rect 7156 11308 8309 11336
rect 7156 11296 7162 11308
rect 8297 11305 8309 11308
rect 8343 11305 8355 11339
rect 8297 11299 8355 11305
rect 14550 11296 14556 11348
rect 14608 11336 14614 11348
rect 15378 11336 15384 11348
rect 14608 11308 15384 11336
rect 14608 11296 14614 11308
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 17402 11296 17408 11348
rect 17460 11336 17466 11348
rect 18785 11339 18843 11345
rect 18785 11336 18797 11339
rect 17460 11308 18797 11336
rect 17460 11296 17466 11308
rect 18785 11305 18797 11308
rect 18831 11305 18843 11339
rect 18785 11299 18843 11305
rect 21266 11296 21272 11348
rect 21324 11296 21330 11348
rect 1854 11228 1860 11280
rect 1912 11228 1918 11280
rect 14182 11268 14188 11280
rect 13464 11240 14188 11268
rect 934 11092 940 11144
rect 992 11132 998 11144
rect 1673 11135 1731 11141
rect 1673 11132 1685 11135
rect 992 11104 1685 11132
rect 992 11092 998 11104
rect 1673 11101 1685 11104
rect 1719 11101 1731 11135
rect 1673 11095 1731 11101
rect 4154 11092 4160 11144
rect 4212 11132 4218 11144
rect 5350 11141 5356 11144
rect 5077 11135 5135 11141
rect 5077 11132 5089 11135
rect 4212 11104 5089 11132
rect 4212 11092 4218 11104
rect 5077 11101 5089 11104
rect 5123 11101 5135 11135
rect 5344 11132 5356 11141
rect 5311 11104 5356 11132
rect 5077 11095 5135 11101
rect 5344 11095 5356 11104
rect 5350 11092 5356 11095
rect 5408 11092 5414 11144
rect 6914 11092 6920 11144
rect 6972 11092 6978 11144
rect 7190 11141 7196 11144
rect 7184 11095 7196 11141
rect 7190 11092 7196 11095
rect 7248 11092 7254 11144
rect 13464 11141 13492 11240
rect 14182 11228 14188 11240
rect 14240 11228 14246 11280
rect 14737 11271 14795 11277
rect 14737 11237 14749 11271
rect 14783 11268 14795 11271
rect 14783 11240 14872 11268
rect 14783 11237 14795 11240
rect 14737 11231 14795 11237
rect 14274 11200 14280 11212
rect 13648 11172 14280 11200
rect 13648 11141 13676 11172
rect 14274 11160 14280 11172
rect 14332 11160 14338 11212
rect 14844 11200 14872 11240
rect 16390 11228 16396 11280
rect 16448 11268 16454 11280
rect 21174 11268 21180 11280
rect 16448 11240 21180 11268
rect 16448 11228 16454 11240
rect 21174 11228 21180 11240
rect 21232 11228 21238 11280
rect 15654 11200 15660 11212
rect 14844 11172 15660 11200
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 15856 11172 16896 11200
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11101 13415 11135
rect 13357 11095 13415 11101
rect 13449 11135 13507 11141
rect 13449 11101 13461 11135
rect 13495 11101 13507 11135
rect 13449 11095 13507 11101
rect 13633 11135 13691 11141
rect 13633 11101 13645 11135
rect 13679 11101 13691 11135
rect 13633 11095 13691 11101
rect 13372 11064 13400 11095
rect 13722 11092 13728 11144
rect 13780 11092 13786 11144
rect 14458 11092 14464 11144
rect 14516 11092 14522 11144
rect 14550 11092 14556 11144
rect 14608 11092 14614 11144
rect 14829 11135 14887 11141
rect 14829 11101 14841 11135
rect 14875 11132 14887 11135
rect 14918 11132 14924 11144
rect 14875 11104 14924 11132
rect 14875 11101 14887 11104
rect 14829 11095 14887 11101
rect 13998 11064 14004 11076
rect 13372 11036 14004 11064
rect 13998 11024 14004 11036
rect 14056 11024 14062 11076
rect 14182 11024 14188 11076
rect 14240 11064 14246 11076
rect 14844 11064 14872 11095
rect 14918 11092 14924 11104
rect 14976 11092 14982 11144
rect 15470 11092 15476 11144
rect 15528 11092 15534 11144
rect 15565 11135 15623 11141
rect 15565 11101 15577 11135
rect 15611 11101 15623 11135
rect 15565 11095 15623 11101
rect 14240 11036 14872 11064
rect 14240 11024 14246 11036
rect 15286 11024 15292 11076
rect 15344 11024 15350 11076
rect 15580 11064 15608 11095
rect 15746 11092 15752 11144
rect 15804 11092 15810 11144
rect 15856 11141 15884 11172
rect 15841 11135 15899 11141
rect 15841 11101 15853 11135
rect 15887 11101 15899 11135
rect 16666 11132 16672 11144
rect 15841 11095 15899 11101
rect 16408 11104 16672 11132
rect 16408 11064 16436 11104
rect 16666 11092 16672 11104
rect 16724 11092 16730 11144
rect 16758 11092 16764 11144
rect 16816 11092 16822 11144
rect 16868 11132 16896 11172
rect 17678 11160 17684 11212
rect 17736 11160 17742 11212
rect 17862 11160 17868 11212
rect 17920 11160 17926 11212
rect 18138 11160 18144 11212
rect 18196 11160 18202 11212
rect 19794 11200 19800 11212
rect 19444 11172 19800 11200
rect 17770 11132 17776 11144
rect 16868 11104 17776 11132
rect 17770 11092 17776 11104
rect 17828 11092 17834 11144
rect 17954 11092 17960 11144
rect 18012 11092 18018 11144
rect 18049 11135 18107 11141
rect 18049 11101 18061 11135
rect 18095 11132 18107 11135
rect 18230 11132 18236 11144
rect 18095 11104 18236 11132
rect 18095 11101 18107 11104
rect 18049 11095 18107 11101
rect 18230 11092 18236 11104
rect 18288 11092 18294 11144
rect 18690 11092 18696 11144
rect 18748 11092 18754 11144
rect 18874 11092 18880 11144
rect 18932 11092 18938 11144
rect 15580 11036 16436 11064
rect 16482 11024 16488 11076
rect 16540 11024 16546 11076
rect 16850 11024 16856 11076
rect 16908 11064 16914 11076
rect 17862 11064 17868 11076
rect 16908 11036 17868 11064
rect 16908 11024 16914 11036
rect 17862 11024 17868 11036
rect 17920 11024 17926 11076
rect 19444 11064 19472 11172
rect 19794 11160 19800 11172
rect 19852 11200 19858 11212
rect 21361 11203 21419 11209
rect 21361 11200 21373 11203
rect 19852 11172 21373 11200
rect 19852 11160 19858 11172
rect 21192 11144 21220 11172
rect 21361 11169 21373 11172
rect 21407 11169 21419 11203
rect 21361 11163 21419 11169
rect 19610 11092 19616 11144
rect 19668 11092 19674 11144
rect 19702 11092 19708 11144
rect 19760 11132 19766 11144
rect 19981 11135 20039 11141
rect 19760 11104 19932 11132
rect 19760 11092 19766 11104
rect 19168 11036 19472 11064
rect 13170 10956 13176 11008
rect 13228 10956 13234 11008
rect 13906 10956 13912 11008
rect 13964 10996 13970 11008
rect 14277 10999 14335 11005
rect 14277 10996 14289 10999
rect 13964 10968 14289 10996
rect 13964 10956 13970 10968
rect 14277 10965 14289 10968
rect 14323 10965 14335 10999
rect 14277 10959 14335 10965
rect 16666 10956 16672 11008
rect 16724 10996 16730 11008
rect 17494 10996 17500 11008
rect 16724 10968 17500 10996
rect 16724 10956 16730 10968
rect 17494 10956 17500 10968
rect 17552 10996 17558 11008
rect 17770 10996 17776 11008
rect 17552 10968 17776 10996
rect 17552 10956 17558 10968
rect 17770 10956 17776 10968
rect 17828 10956 17834 11008
rect 17880 10996 17908 11024
rect 19168 10996 19196 11036
rect 19794 11024 19800 11076
rect 19852 11024 19858 11076
rect 19904 11064 19932 11104
rect 19981 11101 19993 11135
rect 20027 11132 20039 11135
rect 20809 11135 20867 11141
rect 20809 11132 20821 11135
rect 20027 11104 20821 11132
rect 20027 11101 20039 11104
rect 19981 11095 20039 11101
rect 20809 11101 20821 11104
rect 20855 11101 20867 11135
rect 20809 11095 20867 11101
rect 21082 11092 21088 11144
rect 21140 11092 21146 11144
rect 21174 11092 21180 11144
rect 21232 11092 21238 11144
rect 21545 11135 21603 11141
rect 21545 11101 21557 11135
rect 21591 11132 21603 11135
rect 22002 11132 22008 11144
rect 21591 11104 22008 11132
rect 21591 11101 21603 11104
rect 21545 11095 21603 11101
rect 22002 11092 22008 11104
rect 22060 11092 22066 11144
rect 20438 11064 20444 11076
rect 19904 11036 20444 11064
rect 20438 11024 20444 11036
rect 20496 11024 20502 11076
rect 17880 10968 19196 10996
rect 19242 10956 19248 11008
rect 19300 10996 19306 11008
rect 19429 10999 19487 11005
rect 19429 10996 19441 10999
rect 19300 10968 19441 10996
rect 19300 10956 19306 10968
rect 19429 10965 19441 10968
rect 19475 10965 19487 10999
rect 19429 10959 19487 10965
rect 1104 10906 22976 10928
rect 1104 10854 6378 10906
rect 6430 10854 6442 10906
rect 6494 10854 6506 10906
rect 6558 10854 6570 10906
rect 6622 10854 6634 10906
rect 6686 10854 11806 10906
rect 11858 10854 11870 10906
rect 11922 10854 11934 10906
rect 11986 10854 11998 10906
rect 12050 10854 12062 10906
rect 12114 10854 17234 10906
rect 17286 10854 17298 10906
rect 17350 10854 17362 10906
rect 17414 10854 17426 10906
rect 17478 10854 17490 10906
rect 17542 10854 22662 10906
rect 22714 10854 22726 10906
rect 22778 10854 22790 10906
rect 22842 10854 22854 10906
rect 22906 10854 22918 10906
rect 22970 10854 22976 10906
rect 1104 10832 22976 10854
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 3053 10795 3111 10801
rect 3053 10792 3065 10795
rect 2832 10764 3065 10792
rect 2832 10752 2838 10764
rect 3053 10761 3065 10764
rect 3099 10761 3111 10795
rect 3053 10755 3111 10761
rect 4525 10795 4583 10801
rect 4525 10761 4537 10795
rect 4571 10792 4583 10795
rect 4890 10792 4896 10804
rect 4571 10764 4896 10792
rect 4571 10761 4583 10764
rect 4525 10755 4583 10761
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 8573 10795 8631 10801
rect 8573 10761 8585 10795
rect 8619 10792 8631 10795
rect 8662 10792 8668 10804
rect 8619 10764 8668 10792
rect 8619 10761 8631 10764
rect 8573 10755 8631 10761
rect 8662 10752 8668 10764
rect 8720 10752 8726 10804
rect 10870 10752 10876 10804
rect 10928 10752 10934 10804
rect 13722 10792 13728 10804
rect 12268 10764 13728 10792
rect 1946 10733 1952 10736
rect 1940 10724 1952 10733
rect 1907 10696 1952 10724
rect 1940 10687 1952 10696
rect 1946 10684 1952 10687
rect 2004 10684 2010 10736
rect 5534 10684 5540 10736
rect 5592 10724 5598 10736
rect 5638 10727 5696 10733
rect 5638 10724 5650 10727
rect 5592 10696 5650 10724
rect 5592 10684 5598 10696
rect 5638 10693 5650 10696
rect 5684 10693 5696 10727
rect 5638 10687 5696 10693
rect 7460 10727 7518 10733
rect 7460 10693 7472 10727
rect 7506 10724 7518 10727
rect 8202 10724 8208 10736
rect 7506 10696 8208 10724
rect 7506 10693 7518 10696
rect 7460 10687 7518 10693
rect 8202 10684 8208 10696
rect 8260 10684 8266 10736
rect 9766 10733 9772 10736
rect 9760 10724 9772 10733
rect 9727 10696 9772 10724
rect 9760 10687 9772 10696
rect 9766 10684 9772 10687
rect 9824 10684 9830 10736
rect 6914 10656 6920 10668
rect 6886 10616 6920 10656
rect 6972 10656 6978 10668
rect 7193 10659 7251 10665
rect 7193 10656 7205 10659
rect 6972 10628 7205 10656
rect 6972 10616 6978 10628
rect 7193 10625 7205 10628
rect 7239 10625 7251 10659
rect 7193 10619 7251 10625
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 1670 10548 1676 10600
rect 1728 10548 1734 10600
rect 5905 10591 5963 10597
rect 5905 10557 5917 10591
rect 5951 10588 5963 10591
rect 6730 10588 6736 10600
rect 5951 10560 6736 10588
rect 5951 10557 5963 10560
rect 5905 10551 5963 10557
rect 6730 10548 6736 10560
rect 6788 10588 6794 10600
rect 6886 10588 6914 10616
rect 6788 10560 6914 10588
rect 6788 10548 6794 10560
rect 9490 10548 9496 10600
rect 9548 10548 9554 10600
rect 11992 10588 12020 10619
rect 12158 10616 12164 10668
rect 12216 10616 12222 10668
rect 12268 10665 12296 10764
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 13817 10795 13875 10801
rect 13817 10761 13829 10795
rect 13863 10792 13875 10795
rect 14458 10792 14464 10804
rect 13863 10764 14464 10792
rect 13863 10761 13875 10764
rect 13817 10755 13875 10761
rect 14458 10752 14464 10764
rect 14516 10752 14522 10804
rect 15470 10752 15476 10804
rect 15528 10792 15534 10804
rect 15565 10795 15623 10801
rect 15565 10792 15577 10795
rect 15528 10764 15577 10792
rect 15528 10752 15534 10764
rect 15565 10761 15577 10764
rect 15611 10761 15623 10795
rect 15565 10755 15623 10761
rect 16022 10752 16028 10804
rect 16080 10792 16086 10804
rect 18785 10795 18843 10801
rect 16080 10764 17264 10792
rect 16080 10752 16086 10764
rect 13170 10684 13176 10736
rect 13228 10724 13234 10736
rect 13265 10727 13323 10733
rect 13265 10724 13277 10727
rect 13228 10696 13277 10724
rect 13228 10684 13234 10696
rect 13265 10693 13277 10696
rect 13311 10693 13323 10727
rect 13265 10687 13323 10693
rect 15197 10727 15255 10733
rect 15197 10693 15209 10727
rect 15243 10724 15255 10727
rect 16666 10724 16672 10736
rect 15243 10696 16672 10724
rect 15243 10693 15255 10696
rect 15197 10687 15255 10693
rect 16666 10684 16672 10696
rect 16724 10684 16730 10736
rect 12253 10659 12311 10665
rect 12253 10625 12265 10659
rect 12299 10625 12311 10659
rect 12253 10619 12311 10625
rect 12989 10659 13047 10665
rect 12989 10625 13001 10659
rect 13035 10656 13047 10659
rect 13906 10656 13912 10668
rect 13035 10628 13912 10656
rect 13035 10625 13047 10628
rect 12989 10619 13047 10625
rect 13906 10616 13912 10628
rect 13964 10616 13970 10668
rect 14093 10659 14151 10665
rect 14093 10625 14105 10659
rect 14139 10656 14151 10659
rect 15930 10656 15936 10668
rect 14139 10628 15936 10656
rect 14139 10625 14151 10628
rect 14093 10619 14151 10625
rect 15930 10616 15936 10628
rect 15988 10616 15994 10668
rect 16206 10616 16212 10668
rect 16264 10616 16270 10668
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10656 16911 10659
rect 16942 10656 16948 10668
rect 16899 10628 16948 10656
rect 16899 10625 16911 10628
rect 16853 10619 16911 10625
rect 16942 10616 16948 10628
rect 17000 10616 17006 10668
rect 17236 10665 17264 10764
rect 18785 10761 18797 10795
rect 18831 10792 18843 10795
rect 19334 10792 19340 10804
rect 18831 10764 19340 10792
rect 18831 10761 18843 10764
rect 18785 10755 18843 10761
rect 19334 10752 19340 10764
rect 19392 10752 19398 10804
rect 19426 10752 19432 10804
rect 19484 10792 19490 10804
rect 19610 10792 19616 10804
rect 19484 10764 19616 10792
rect 19484 10752 19490 10764
rect 19610 10752 19616 10764
rect 19668 10752 19674 10804
rect 20990 10752 20996 10804
rect 21048 10752 21054 10804
rect 17954 10684 17960 10736
rect 18012 10724 18018 10736
rect 19245 10727 19303 10733
rect 19245 10724 19257 10727
rect 18012 10696 19257 10724
rect 18012 10684 18018 10696
rect 19245 10693 19257 10696
rect 19291 10693 19303 10727
rect 19245 10687 19303 10693
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 17129 10659 17187 10665
rect 17129 10625 17141 10659
rect 17175 10625 17187 10659
rect 17129 10619 17187 10625
rect 17221 10659 17279 10665
rect 17221 10625 17233 10659
rect 17267 10625 17279 10659
rect 17221 10619 17279 10625
rect 12342 10588 12348 10600
rect 11992 10560 12348 10588
rect 12342 10548 12348 10560
rect 12400 10548 12406 10600
rect 12894 10548 12900 10600
rect 12952 10548 12958 10600
rect 13357 10591 13415 10597
rect 13357 10557 13369 10591
rect 13403 10557 13415 10591
rect 13357 10551 13415 10557
rect 13817 10591 13875 10597
rect 13817 10557 13829 10591
rect 13863 10557 13875 10591
rect 13817 10551 13875 10557
rect 11977 10523 12035 10529
rect 11977 10489 11989 10523
rect 12023 10520 12035 10523
rect 13078 10520 13084 10532
rect 12023 10492 13084 10520
rect 12023 10489 12035 10492
rect 11977 10483 12035 10489
rect 13078 10480 13084 10492
rect 13136 10520 13142 10532
rect 13372 10520 13400 10551
rect 13136 10492 13400 10520
rect 13832 10520 13860 10551
rect 13998 10548 14004 10600
rect 14056 10588 14062 10600
rect 15010 10588 15016 10600
rect 14056 10560 15016 10588
rect 14056 10548 14062 10560
rect 15010 10548 15016 10560
rect 15068 10548 15074 10600
rect 15102 10548 15108 10600
rect 15160 10548 15166 10600
rect 16298 10548 16304 10600
rect 16356 10588 16362 10600
rect 17052 10588 17080 10619
rect 16356 10560 17080 10588
rect 16356 10548 16362 10560
rect 14182 10520 14188 10532
rect 13832 10492 14188 10520
rect 13136 10480 13142 10492
rect 14182 10480 14188 10492
rect 14240 10480 14246 10532
rect 16942 10480 16948 10532
rect 17000 10520 17006 10532
rect 17144 10520 17172 10619
rect 17402 10616 17408 10668
rect 17460 10656 17466 10668
rect 18509 10659 18567 10665
rect 18509 10656 18521 10659
rect 17460 10628 18521 10656
rect 17460 10616 17466 10628
rect 18509 10625 18521 10628
rect 18555 10625 18567 10659
rect 18509 10619 18567 10625
rect 19426 10616 19432 10668
rect 19484 10616 19490 10668
rect 19521 10659 19579 10665
rect 19521 10625 19533 10659
rect 19567 10625 19579 10659
rect 19521 10619 19579 10625
rect 17862 10548 17868 10600
rect 17920 10588 17926 10600
rect 18325 10591 18383 10597
rect 18325 10588 18337 10591
rect 17920 10560 18337 10588
rect 17920 10548 17926 10560
rect 18325 10557 18337 10560
rect 18371 10557 18383 10591
rect 18325 10551 18383 10557
rect 18414 10548 18420 10600
rect 18472 10548 18478 10600
rect 18601 10591 18659 10597
rect 18601 10557 18613 10591
rect 18647 10588 18659 10591
rect 18874 10588 18880 10600
rect 18647 10560 18880 10588
rect 18647 10557 18659 10560
rect 18601 10551 18659 10557
rect 18616 10520 18644 10551
rect 18874 10548 18880 10560
rect 18932 10588 18938 10600
rect 19536 10588 19564 10619
rect 19702 10616 19708 10668
rect 19760 10616 19766 10668
rect 19797 10659 19855 10665
rect 19797 10625 19809 10659
rect 19843 10625 19855 10659
rect 19797 10619 19855 10625
rect 18932 10560 19564 10588
rect 18932 10548 18938 10560
rect 19610 10548 19616 10600
rect 19668 10588 19674 10600
rect 19812 10588 19840 10619
rect 20622 10616 20628 10668
rect 20680 10656 20686 10668
rect 22005 10659 22063 10665
rect 22005 10656 22017 10659
rect 20680 10628 22017 10656
rect 20680 10616 20686 10628
rect 22005 10625 22017 10628
rect 22051 10625 22063 10659
rect 22005 10619 22063 10625
rect 22186 10616 22192 10668
rect 22244 10616 22250 10668
rect 19668 10560 19840 10588
rect 19668 10548 19674 10560
rect 21266 10548 21272 10600
rect 21324 10588 21330 10600
rect 21453 10591 21511 10597
rect 21453 10588 21465 10591
rect 21324 10560 21465 10588
rect 21324 10548 21330 10560
rect 21453 10557 21465 10560
rect 21499 10557 21511 10591
rect 21453 10551 21511 10557
rect 21542 10548 21548 10600
rect 21600 10588 21606 10600
rect 22204 10588 22232 10616
rect 21600 10560 22232 10588
rect 21600 10548 21606 10560
rect 17000 10492 18644 10520
rect 21085 10523 21143 10529
rect 17000 10480 17006 10492
rect 21085 10489 21097 10523
rect 21131 10489 21143 10523
rect 21085 10483 21143 10489
rect 11238 10412 11244 10464
rect 11296 10452 11302 10464
rect 12713 10455 12771 10461
rect 12713 10452 12725 10455
rect 11296 10424 12725 10452
rect 11296 10412 11302 10424
rect 12713 10421 12725 10424
rect 12759 10421 12771 10455
rect 12713 10415 12771 10421
rect 13262 10412 13268 10464
rect 13320 10452 13326 10464
rect 16117 10455 16175 10461
rect 16117 10452 16129 10455
rect 13320 10424 16129 10452
rect 13320 10412 13326 10424
rect 16117 10421 16129 10424
rect 16163 10452 16175 10455
rect 16758 10452 16764 10464
rect 16163 10424 16764 10452
rect 16163 10421 16175 10424
rect 16117 10415 16175 10421
rect 16758 10412 16764 10424
rect 16816 10452 16822 10464
rect 17402 10452 17408 10464
rect 16816 10424 17408 10452
rect 16816 10412 16822 10424
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 17494 10412 17500 10464
rect 17552 10412 17558 10464
rect 17862 10412 17868 10464
rect 17920 10452 17926 10464
rect 21100 10452 21128 10483
rect 17920 10424 21128 10452
rect 17920 10412 17926 10424
rect 22002 10412 22008 10464
rect 22060 10412 22066 10464
rect 1104 10362 22816 10384
rect 1104 10310 3664 10362
rect 3716 10310 3728 10362
rect 3780 10310 3792 10362
rect 3844 10310 3856 10362
rect 3908 10310 3920 10362
rect 3972 10310 9092 10362
rect 9144 10310 9156 10362
rect 9208 10310 9220 10362
rect 9272 10310 9284 10362
rect 9336 10310 9348 10362
rect 9400 10310 14520 10362
rect 14572 10310 14584 10362
rect 14636 10310 14648 10362
rect 14700 10310 14712 10362
rect 14764 10310 14776 10362
rect 14828 10310 19948 10362
rect 20000 10310 20012 10362
rect 20064 10310 20076 10362
rect 20128 10310 20140 10362
rect 20192 10310 20204 10362
rect 20256 10310 22816 10362
rect 1104 10288 22816 10310
rect 2406 10208 2412 10260
rect 2464 10248 2470 10260
rect 3053 10251 3111 10257
rect 3053 10248 3065 10251
rect 2464 10220 3065 10248
rect 2464 10208 2470 10220
rect 3053 10217 3065 10220
rect 3099 10217 3111 10251
rect 3053 10211 3111 10217
rect 5074 10208 5080 10260
rect 5132 10248 5138 10260
rect 5537 10251 5595 10257
rect 5537 10248 5549 10251
rect 5132 10220 5549 10248
rect 5132 10208 5138 10220
rect 5537 10217 5549 10220
rect 5583 10217 5595 10251
rect 5537 10211 5595 10217
rect 8478 10208 8484 10260
rect 8536 10208 8542 10260
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 10873 10251 10931 10257
rect 10873 10248 10885 10251
rect 9732 10220 10885 10248
rect 9732 10208 9738 10220
rect 10873 10217 10885 10220
rect 10919 10217 10931 10251
rect 10873 10211 10931 10217
rect 12894 10208 12900 10260
rect 12952 10248 12958 10260
rect 13449 10251 13507 10257
rect 13449 10248 13461 10251
rect 12952 10220 13461 10248
rect 12952 10208 12958 10220
rect 13449 10217 13461 10220
rect 13495 10248 13507 10251
rect 13630 10248 13636 10260
rect 13495 10220 13636 10248
rect 13495 10217 13507 10220
rect 13449 10211 13507 10217
rect 13630 10208 13636 10220
rect 13688 10208 13694 10260
rect 15654 10208 15660 10260
rect 15712 10208 15718 10260
rect 16206 10208 16212 10260
rect 16264 10248 16270 10260
rect 16945 10251 17003 10257
rect 16945 10248 16957 10251
rect 16264 10220 16957 10248
rect 16264 10208 16270 10220
rect 16945 10217 16957 10220
rect 16991 10217 17003 10251
rect 16945 10211 17003 10217
rect 19610 10208 19616 10260
rect 19668 10208 19674 10260
rect 19794 10208 19800 10260
rect 19852 10248 19858 10260
rect 19981 10251 20039 10257
rect 19981 10248 19993 10251
rect 19852 10220 19993 10248
rect 19852 10208 19858 10220
rect 19981 10217 19993 10220
rect 20027 10217 20039 10251
rect 19981 10211 20039 10217
rect 20530 10208 20536 10260
rect 20588 10248 20594 10260
rect 20625 10251 20683 10257
rect 20625 10248 20637 10251
rect 20588 10220 20637 10248
rect 20588 10208 20594 10220
rect 20625 10217 20637 10220
rect 20671 10217 20683 10251
rect 20625 10211 20683 10217
rect 17494 10180 17500 10192
rect 13556 10152 17500 10180
rect 4154 10072 4160 10124
rect 4212 10072 4218 10124
rect 6730 10072 6736 10124
rect 6788 10112 6794 10124
rect 13556 10121 13584 10152
rect 17494 10140 17500 10152
rect 17552 10140 17558 10192
rect 20441 10183 20499 10189
rect 20441 10149 20453 10183
rect 20487 10149 20499 10183
rect 20441 10143 20499 10149
rect 7101 10115 7159 10121
rect 7101 10112 7113 10115
rect 6788 10084 7113 10112
rect 6788 10072 6794 10084
rect 7101 10081 7113 10084
rect 7147 10081 7159 10115
rect 7101 10075 7159 10081
rect 13541 10115 13599 10121
rect 13541 10081 13553 10115
rect 13587 10081 13599 10115
rect 13541 10075 13599 10081
rect 16301 10115 16359 10121
rect 16301 10081 16313 10115
rect 16347 10112 16359 10115
rect 16942 10112 16948 10124
rect 16347 10084 16948 10112
rect 16347 10081 16359 10084
rect 16301 10075 16359 10081
rect 1670 10004 1676 10056
rect 1728 10004 1734 10056
rect 1762 10004 1768 10056
rect 1820 10044 1826 10056
rect 4430 10053 4436 10056
rect 1929 10047 1987 10053
rect 1929 10044 1941 10047
rect 1820 10016 1941 10044
rect 1820 10004 1826 10016
rect 1929 10013 1941 10016
rect 1975 10013 1987 10047
rect 4424 10044 4436 10053
rect 4391 10016 4436 10044
rect 1929 10007 1987 10013
rect 4424 10007 4436 10016
rect 4430 10004 4436 10007
rect 4488 10004 4494 10056
rect 7116 10044 7144 10075
rect 16942 10072 16948 10084
rect 17000 10072 17006 10124
rect 19702 10072 19708 10124
rect 19760 10112 19766 10124
rect 20456 10112 20484 10143
rect 19760 10084 20484 10112
rect 19760 10072 19766 10084
rect 9490 10044 9496 10056
rect 7116 10016 9496 10044
rect 9490 10004 9496 10016
rect 9548 10004 9554 10056
rect 9760 10047 9818 10053
rect 9760 10013 9772 10047
rect 9806 10044 9818 10047
rect 10962 10044 10968 10056
rect 9806 10016 10968 10044
rect 9806 10013 9818 10016
rect 9760 10007 9818 10013
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 13078 10044 13084 10056
rect 13039 10016 13084 10044
rect 13078 10004 13084 10016
rect 13136 10004 13142 10056
rect 16666 10044 16672 10056
rect 15028 10016 16672 10044
rect 7368 9979 7426 9985
rect 7368 9945 7380 9979
rect 7414 9976 7426 9979
rect 8110 9976 8116 9988
rect 7414 9948 8116 9976
rect 7414 9945 7426 9948
rect 7368 9939 7426 9945
rect 8110 9936 8116 9948
rect 8168 9936 8174 9988
rect 12342 9936 12348 9988
rect 12400 9976 12406 9988
rect 15028 9976 15056 10016
rect 16666 10004 16672 10016
rect 16724 10004 16730 10056
rect 16758 10004 16764 10056
rect 16816 10044 16822 10056
rect 17037 10047 17095 10053
rect 17037 10044 17049 10047
rect 16816 10016 17049 10044
rect 16816 10004 16822 10016
rect 17037 10013 17049 10016
rect 17083 10044 17095 10047
rect 17586 10044 17592 10056
rect 17083 10016 17592 10044
rect 17083 10013 17095 10016
rect 17037 10007 17095 10013
rect 17586 10004 17592 10016
rect 17644 10004 17650 10056
rect 19429 10047 19487 10053
rect 19429 10013 19441 10047
rect 19475 10044 19487 10047
rect 19794 10044 19800 10056
rect 19475 10016 19800 10044
rect 19475 10013 19487 10016
rect 19429 10007 19487 10013
rect 19794 10004 19800 10016
rect 19852 10044 19858 10056
rect 20346 10044 20352 10056
rect 19852 10016 20352 10044
rect 19852 10004 19858 10016
rect 20346 10004 20352 10016
rect 20404 10004 20410 10056
rect 12400 9948 15056 9976
rect 12400 9936 12406 9948
rect 15102 9936 15108 9988
rect 15160 9976 15166 9988
rect 20809 9979 20867 9985
rect 20809 9976 20821 9979
rect 15160 9948 20821 9976
rect 15160 9936 15166 9948
rect 20809 9945 20821 9948
rect 20855 9976 20867 9979
rect 21266 9976 21272 9988
rect 20855 9948 21272 9976
rect 20855 9945 20867 9948
rect 20809 9939 20867 9945
rect 21266 9936 21272 9948
rect 21324 9936 21330 9988
rect 12710 9868 12716 9920
rect 12768 9908 12774 9920
rect 12897 9911 12955 9917
rect 12897 9908 12909 9911
rect 12768 9880 12909 9908
rect 12768 9868 12774 9880
rect 12897 9877 12909 9880
rect 12943 9877 12955 9911
rect 12897 9871 12955 9877
rect 13078 9868 13084 9920
rect 13136 9868 13142 9920
rect 16022 9868 16028 9920
rect 16080 9868 16086 9920
rect 16117 9911 16175 9917
rect 16117 9877 16129 9911
rect 16163 9908 16175 9911
rect 16206 9908 16212 9920
rect 16163 9880 16212 9908
rect 16163 9877 16175 9880
rect 16117 9871 16175 9877
rect 16206 9868 16212 9880
rect 16264 9868 16270 9920
rect 20254 9868 20260 9920
rect 20312 9908 20318 9920
rect 20599 9911 20657 9917
rect 20599 9908 20611 9911
rect 20312 9880 20611 9908
rect 20312 9868 20318 9880
rect 20599 9877 20611 9880
rect 20645 9908 20657 9911
rect 20714 9908 20720 9920
rect 20645 9880 20720 9908
rect 20645 9877 20657 9880
rect 20599 9871 20657 9877
rect 20714 9868 20720 9880
rect 20772 9868 20778 9920
rect 1104 9818 22976 9840
rect 1104 9766 6378 9818
rect 6430 9766 6442 9818
rect 6494 9766 6506 9818
rect 6558 9766 6570 9818
rect 6622 9766 6634 9818
rect 6686 9766 11806 9818
rect 11858 9766 11870 9818
rect 11922 9766 11934 9818
rect 11986 9766 11998 9818
rect 12050 9766 12062 9818
rect 12114 9766 17234 9818
rect 17286 9766 17298 9818
rect 17350 9766 17362 9818
rect 17414 9766 17426 9818
rect 17478 9766 17490 9818
rect 17542 9766 22662 9818
rect 22714 9766 22726 9818
rect 22778 9766 22790 9818
rect 22842 9766 22854 9818
rect 22906 9766 22918 9818
rect 22970 9766 22976 9818
rect 1104 9744 22976 9766
rect 9766 9664 9772 9716
rect 9824 9704 9830 9716
rect 12158 9704 12164 9716
rect 9824 9676 12164 9704
rect 9824 9664 9830 9676
rect 12158 9664 12164 9676
rect 12216 9704 12222 9716
rect 14182 9704 14188 9716
rect 12216 9676 14188 9704
rect 12216 9664 12222 9676
rect 14182 9664 14188 9676
rect 14240 9664 14246 9716
rect 15010 9664 15016 9716
rect 15068 9704 15074 9716
rect 15841 9707 15899 9713
rect 15841 9704 15853 9707
rect 15068 9676 15853 9704
rect 15068 9664 15074 9676
rect 15841 9673 15853 9676
rect 15887 9673 15899 9707
rect 15841 9667 15899 9673
rect 16482 9664 16488 9716
rect 16540 9664 16546 9716
rect 16942 9664 16948 9716
rect 17000 9664 17006 9716
rect 17126 9664 17132 9716
rect 17184 9704 17190 9716
rect 17678 9704 17684 9716
rect 17184 9676 17684 9704
rect 17184 9664 17190 9676
rect 17678 9664 17684 9676
rect 17736 9704 17742 9716
rect 17862 9704 17868 9716
rect 17736 9676 17868 9704
rect 17736 9664 17742 9676
rect 17862 9664 17868 9676
rect 17920 9664 17926 9716
rect 19242 9664 19248 9716
rect 19300 9704 19306 9716
rect 20622 9704 20628 9716
rect 19300 9676 20628 9704
rect 19300 9664 19306 9676
rect 20622 9664 20628 9676
rect 20680 9664 20686 9716
rect 1670 9596 1676 9648
rect 1728 9636 1734 9648
rect 2866 9636 2872 9648
rect 1728 9608 2872 9636
rect 1728 9596 1734 9608
rect 1780 9577 1808 9608
rect 2866 9596 2872 9608
rect 2924 9636 2930 9648
rect 9858 9645 9864 9648
rect 9852 9636 9864 9645
rect 2924 9608 4200 9636
rect 9819 9608 9864 9636
rect 2924 9596 2930 9608
rect 4172 9580 4200 9608
rect 9852 9599 9864 9608
rect 9858 9596 9864 9599
rect 9916 9596 9922 9648
rect 16500 9636 16528 9664
rect 15764 9608 17172 9636
rect 2038 9577 2044 9580
rect 1765 9571 1823 9577
rect 1765 9537 1777 9571
rect 1811 9537 1823 9571
rect 2032 9568 2044 9577
rect 1999 9540 2044 9568
rect 1765 9531 1823 9537
rect 2032 9531 2044 9540
rect 2038 9528 2044 9531
rect 2096 9528 2102 9580
rect 4154 9528 4160 9580
rect 4212 9568 4218 9580
rect 4522 9577 4528 9580
rect 4249 9571 4307 9577
rect 4249 9568 4261 9571
rect 4212 9540 4261 9568
rect 4212 9528 4218 9540
rect 4249 9537 4261 9540
rect 4295 9537 4307 9571
rect 4516 9568 4528 9577
rect 4483 9540 4528 9568
rect 4249 9531 4307 9537
rect 4516 9531 4528 9540
rect 4522 9528 4528 9531
rect 4580 9528 4586 9580
rect 9490 9528 9496 9580
rect 9548 9568 9554 9580
rect 15764 9577 15792 9608
rect 9585 9571 9643 9577
rect 9585 9568 9597 9571
rect 9548 9540 9597 9568
rect 9548 9528 9554 9540
rect 9585 9537 9597 9540
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 15749 9571 15807 9577
rect 15749 9537 15761 9571
rect 15795 9537 15807 9571
rect 15749 9531 15807 9537
rect 15933 9571 15991 9577
rect 15933 9537 15945 9571
rect 15979 9568 15991 9571
rect 16482 9568 16488 9580
rect 15979 9540 16488 9568
rect 15979 9537 15991 9540
rect 15933 9531 15991 9537
rect 16482 9528 16488 9540
rect 16540 9528 16546 9580
rect 16850 9528 16856 9580
rect 16908 9528 16914 9580
rect 17144 9577 17172 9608
rect 17586 9596 17592 9648
rect 17644 9636 17650 9648
rect 18049 9639 18107 9645
rect 17644 9608 17908 9636
rect 17644 9596 17650 9608
rect 17880 9580 17908 9608
rect 18049 9605 18061 9639
rect 18095 9636 18107 9639
rect 18095 9608 20944 9636
rect 18095 9605 18107 9608
rect 18049 9599 18107 9605
rect 17129 9571 17187 9577
rect 17129 9537 17141 9571
rect 17175 9537 17187 9571
rect 17129 9531 17187 9537
rect 17144 9500 17172 9531
rect 17218 9528 17224 9580
rect 17276 9568 17282 9580
rect 17770 9568 17776 9580
rect 17276 9540 17776 9568
rect 17276 9528 17282 9540
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 17862 9528 17868 9580
rect 17920 9568 17926 9580
rect 18509 9571 18567 9577
rect 18509 9568 18521 9571
rect 17920 9540 18521 9568
rect 17920 9528 17926 9540
rect 18509 9537 18521 9540
rect 18555 9537 18567 9571
rect 18509 9531 18567 9537
rect 18693 9571 18751 9577
rect 18693 9537 18705 9571
rect 18739 9537 18751 9571
rect 18693 9531 18751 9537
rect 17144 9472 18000 9500
rect 3050 9392 3056 9444
rect 3108 9432 3114 9444
rect 3145 9435 3203 9441
rect 3145 9432 3157 9435
rect 3108 9404 3157 9432
rect 3108 9392 3114 9404
rect 3145 9401 3157 9404
rect 3191 9401 3203 9435
rect 3145 9395 3203 9401
rect 5258 9392 5264 9444
rect 5316 9432 5322 9444
rect 5629 9435 5687 9441
rect 5629 9432 5641 9435
rect 5316 9404 5641 9432
rect 5316 9392 5322 9404
rect 5629 9401 5641 9404
rect 5675 9401 5687 9435
rect 5629 9395 5687 9401
rect 10965 9435 11023 9441
rect 10965 9401 10977 9435
rect 11011 9432 11023 9435
rect 11698 9432 11704 9444
rect 11011 9404 11704 9432
rect 11011 9401 11023 9404
rect 10965 9395 11023 9401
rect 11698 9392 11704 9404
rect 11756 9392 11762 9444
rect 17678 9392 17684 9444
rect 17736 9432 17742 9444
rect 17865 9435 17923 9441
rect 17865 9432 17877 9435
rect 17736 9404 17877 9432
rect 17736 9392 17742 9404
rect 17865 9401 17877 9404
rect 17911 9401 17923 9435
rect 17865 9395 17923 9401
rect 17129 9367 17187 9373
rect 17129 9333 17141 9367
rect 17175 9364 17187 9367
rect 17770 9364 17776 9376
rect 17175 9336 17776 9364
rect 17175 9333 17187 9336
rect 17129 9327 17187 9333
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 17972 9364 18000 9472
rect 18046 9460 18052 9512
rect 18104 9500 18110 9512
rect 18414 9500 18420 9512
rect 18104 9472 18420 9500
rect 18104 9460 18110 9472
rect 18414 9460 18420 9472
rect 18472 9500 18478 9512
rect 18708 9500 18736 9531
rect 18782 9528 18788 9580
rect 18840 9528 18846 9580
rect 20714 9528 20720 9580
rect 20772 9568 20778 9580
rect 20916 9577 20944 9608
rect 20990 9596 20996 9648
rect 21048 9636 21054 9648
rect 21177 9639 21235 9645
rect 21177 9636 21189 9639
rect 21048 9608 21189 9636
rect 21048 9596 21054 9608
rect 21177 9605 21189 9608
rect 21223 9636 21235 9639
rect 21542 9636 21548 9648
rect 21223 9608 21548 9636
rect 21223 9605 21235 9608
rect 21177 9599 21235 9605
rect 21542 9596 21548 9608
rect 21600 9596 21606 9648
rect 20809 9571 20867 9577
rect 20809 9568 20821 9571
rect 20772 9540 20821 9568
rect 20772 9528 20778 9540
rect 20809 9537 20821 9540
rect 20855 9537 20867 9571
rect 20809 9531 20867 9537
rect 20902 9571 20960 9577
rect 20902 9537 20914 9571
rect 20948 9537 20960 9571
rect 20902 9531 20960 9537
rect 21085 9571 21143 9577
rect 21085 9537 21097 9571
rect 21131 9537 21143 9571
rect 21085 9531 21143 9537
rect 18472 9472 18736 9500
rect 18472 9460 18478 9472
rect 18506 9392 18512 9444
rect 18564 9392 18570 9444
rect 20254 9392 20260 9444
rect 20312 9432 20318 9444
rect 20622 9432 20628 9444
rect 20312 9404 20628 9432
rect 20312 9392 20318 9404
rect 20622 9392 20628 9404
rect 20680 9432 20686 9444
rect 21100 9432 21128 9531
rect 21266 9528 21272 9580
rect 21324 9577 21330 9580
rect 21324 9568 21332 9577
rect 22005 9571 22063 9577
rect 22005 9568 22017 9571
rect 21324 9540 22017 9568
rect 21324 9531 21332 9540
rect 22005 9537 22017 9540
rect 22051 9537 22063 9571
rect 22005 9531 22063 9537
rect 21324 9528 21330 9531
rect 22094 9528 22100 9580
rect 22152 9568 22158 9580
rect 22189 9571 22247 9577
rect 22189 9568 22201 9571
rect 22152 9540 22201 9568
rect 22152 9528 22158 9540
rect 22189 9537 22201 9540
rect 22235 9537 22247 9571
rect 22189 9531 22247 9537
rect 20680 9404 21128 9432
rect 20680 9392 20686 9404
rect 20272 9364 20300 9392
rect 17972 9336 20300 9364
rect 20714 9324 20720 9376
rect 20772 9364 20778 9376
rect 21082 9364 21088 9376
rect 20772 9336 21088 9364
rect 20772 9324 20778 9336
rect 21082 9324 21088 9336
rect 21140 9324 21146 9376
rect 21266 9324 21272 9376
rect 21324 9364 21330 9376
rect 21453 9367 21511 9373
rect 21453 9364 21465 9367
rect 21324 9336 21465 9364
rect 21324 9324 21330 9336
rect 21453 9333 21465 9336
rect 21499 9333 21511 9367
rect 21453 9327 21511 9333
rect 22002 9324 22008 9376
rect 22060 9324 22066 9376
rect 1104 9274 22816 9296
rect 1104 9222 3664 9274
rect 3716 9222 3728 9274
rect 3780 9222 3792 9274
rect 3844 9222 3856 9274
rect 3908 9222 3920 9274
rect 3972 9222 9092 9274
rect 9144 9222 9156 9274
rect 9208 9222 9220 9274
rect 9272 9222 9284 9274
rect 9336 9222 9348 9274
rect 9400 9222 14520 9274
rect 14572 9222 14584 9274
rect 14636 9222 14648 9274
rect 14700 9222 14712 9274
rect 14764 9222 14776 9274
rect 14828 9222 19948 9274
rect 20000 9222 20012 9274
rect 20064 9222 20076 9274
rect 20128 9222 20140 9274
rect 20192 9222 20204 9274
rect 20256 9222 22816 9274
rect 1104 9200 22816 9222
rect 3326 9120 3332 9172
rect 3384 9160 3390 9172
rect 3421 9163 3479 9169
rect 3421 9160 3433 9163
rect 3384 9132 3433 9160
rect 3384 9120 3390 9132
rect 3421 9129 3433 9132
rect 3467 9129 3479 9163
rect 3421 9123 3479 9129
rect 10873 9163 10931 9169
rect 10873 9129 10885 9163
rect 10919 9160 10931 9163
rect 11054 9160 11060 9172
rect 10919 9132 11060 9160
rect 10919 9129 10931 9132
rect 10873 9123 10931 9129
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 13078 9120 13084 9172
rect 13136 9120 13142 9172
rect 14921 9163 14979 9169
rect 14921 9129 14933 9163
rect 14967 9160 14979 9163
rect 15102 9160 15108 9172
rect 14967 9132 15108 9160
rect 14967 9129 14979 9132
rect 14921 9123 14979 9129
rect 15102 9120 15108 9132
rect 15160 9120 15166 9172
rect 19334 9160 19340 9172
rect 15212 9132 19340 9160
rect 15212 9092 15240 9132
rect 19334 9120 19340 9132
rect 19392 9120 19398 9172
rect 12406 9064 15240 9092
rect 1670 8984 1676 9036
rect 1728 9024 1734 9036
rect 2041 9027 2099 9033
rect 2041 9024 2053 9027
rect 1728 8996 2053 9024
rect 1728 8984 1734 8996
rect 2041 8993 2053 8996
rect 2087 8993 2099 9027
rect 2041 8987 2099 8993
rect 9490 8984 9496 9036
rect 9548 8984 9554 9036
rect 2308 8959 2366 8965
rect 2308 8925 2320 8959
rect 2354 8956 2366 8959
rect 2590 8956 2596 8968
rect 2354 8928 2596 8956
rect 2354 8925 2366 8928
rect 2308 8919 2366 8925
rect 2590 8916 2596 8928
rect 2648 8916 2654 8968
rect 9760 8959 9818 8965
rect 9760 8925 9772 8959
rect 9806 8956 9818 8959
rect 12406 8956 12434 9064
rect 16574 9052 16580 9104
rect 16632 9092 16638 9104
rect 17313 9095 17371 9101
rect 17313 9092 17325 9095
rect 16632 9064 17325 9092
rect 16632 9052 16638 9064
rect 17313 9061 17325 9064
rect 17359 9061 17371 9095
rect 17313 9055 17371 9061
rect 20438 9052 20444 9104
rect 20496 9092 20502 9104
rect 20993 9095 21051 9101
rect 20993 9092 21005 9095
rect 20496 9064 21005 9092
rect 20496 9052 20502 9064
rect 20993 9061 21005 9064
rect 21039 9061 21051 9095
rect 20993 9055 21051 9061
rect 12802 8984 12808 9036
rect 12860 9024 12866 9036
rect 14553 9027 14611 9033
rect 14553 9024 14565 9027
rect 12860 8996 14565 9024
rect 12860 8984 12866 8996
rect 14553 8993 14565 8996
rect 14599 8993 14611 9027
rect 14553 8987 14611 8993
rect 15657 9027 15715 9033
rect 15657 8993 15669 9027
rect 15703 9024 15715 9027
rect 16758 9024 16764 9036
rect 15703 8996 16764 9024
rect 15703 8993 15715 8996
rect 15657 8987 15715 8993
rect 9806 8928 12434 8956
rect 12989 8959 13047 8965
rect 9806 8925 9818 8928
rect 9760 8919 9818 8925
rect 12989 8925 13001 8959
rect 13035 8925 13047 8959
rect 12989 8919 13047 8925
rect 13173 8959 13231 8965
rect 13173 8925 13185 8959
rect 13219 8956 13231 8959
rect 13354 8956 13360 8968
rect 13219 8928 13360 8956
rect 13219 8925 13231 8928
rect 13173 8919 13231 8925
rect 13004 8888 13032 8919
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 14737 8959 14795 8965
rect 14737 8925 14749 8959
rect 14783 8956 14795 8959
rect 14918 8956 14924 8968
rect 14783 8928 14924 8956
rect 14783 8925 14795 8928
rect 14737 8919 14795 8925
rect 14918 8916 14924 8928
rect 14976 8916 14982 8968
rect 16408 8965 16436 8996
rect 16758 8984 16764 8996
rect 16816 8984 16822 9036
rect 16942 8984 16948 9036
rect 17000 9024 17006 9036
rect 18049 9027 18107 9033
rect 18049 9024 18061 9027
rect 17000 8996 18061 9024
rect 17000 8984 17006 8996
rect 18049 8993 18061 8996
rect 18095 8993 18107 9027
rect 18049 8987 18107 8993
rect 18230 8984 18236 9036
rect 18288 9024 18294 9036
rect 22002 9024 22008 9036
rect 18288 8996 19380 9024
rect 18288 8984 18294 8996
rect 15749 8959 15807 8965
rect 15749 8925 15761 8959
rect 15795 8925 15807 8959
rect 15749 8919 15807 8925
rect 16393 8959 16451 8965
rect 16393 8925 16405 8959
rect 16439 8925 16451 8959
rect 16393 8919 16451 8925
rect 13262 8888 13268 8900
rect 13004 8860 13268 8888
rect 13262 8848 13268 8860
rect 13320 8848 13326 8900
rect 13538 8848 13544 8900
rect 13596 8888 13602 8900
rect 15473 8891 15531 8897
rect 15473 8888 15485 8891
rect 13596 8860 15485 8888
rect 13596 8848 13602 8860
rect 15473 8857 15485 8860
rect 15519 8857 15531 8891
rect 15764 8888 15792 8919
rect 16482 8916 16488 8968
rect 16540 8956 16546 8968
rect 16669 8959 16727 8965
rect 16669 8956 16681 8959
rect 16540 8928 16681 8956
rect 16540 8916 16546 8928
rect 16669 8925 16681 8928
rect 16715 8925 16727 8959
rect 16669 8919 16727 8925
rect 17405 8959 17463 8965
rect 17405 8925 17417 8959
rect 17451 8925 17463 8959
rect 17405 8919 17463 8925
rect 16942 8888 16948 8900
rect 15764 8860 16948 8888
rect 15473 8851 15531 8857
rect 16942 8848 16948 8860
rect 17000 8848 17006 8900
rect 17420 8888 17448 8919
rect 17586 8916 17592 8968
rect 17644 8916 17650 8968
rect 18417 8959 18475 8965
rect 18417 8925 18429 8959
rect 18463 8956 18475 8959
rect 19242 8956 19248 8968
rect 18463 8928 19248 8956
rect 18463 8925 18475 8928
rect 18417 8919 18475 8925
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 17678 8888 17684 8900
rect 17420 8860 17684 8888
rect 17678 8848 17684 8860
rect 17736 8888 17742 8900
rect 18601 8891 18659 8897
rect 18601 8888 18613 8891
rect 17736 8860 18613 8888
rect 17736 8848 17742 8860
rect 18601 8857 18613 8860
rect 18647 8888 18659 8891
rect 18782 8888 18788 8900
rect 18647 8860 18788 8888
rect 18647 8857 18659 8860
rect 18601 8851 18659 8857
rect 18782 8848 18788 8860
rect 18840 8848 18846 8900
rect 19352 8888 19380 8996
rect 20824 8996 22008 9024
rect 20824 8965 20852 8996
rect 22002 8984 22008 8996
rect 22060 8984 22066 9036
rect 20809 8959 20867 8965
rect 20809 8925 20821 8959
rect 20855 8925 20867 8959
rect 20809 8919 20867 8925
rect 20901 8959 20959 8965
rect 20901 8925 20913 8959
rect 20947 8925 20959 8959
rect 20901 8919 20959 8925
rect 21085 8959 21143 8965
rect 21085 8925 21097 8959
rect 21131 8956 21143 8959
rect 21174 8956 21180 8968
rect 21131 8928 21180 8956
rect 21131 8925 21143 8928
rect 21085 8919 21143 8925
rect 20916 8888 20944 8919
rect 21174 8916 21180 8928
rect 21232 8916 21238 8968
rect 21266 8916 21272 8968
rect 21324 8916 21330 8968
rect 19352 8860 20944 8888
rect 15010 8780 15016 8832
rect 15068 8820 15074 8832
rect 15749 8823 15807 8829
rect 15749 8820 15761 8823
rect 15068 8792 15761 8820
rect 15068 8780 15074 8792
rect 15749 8789 15761 8792
rect 15795 8789 15807 8823
rect 15749 8783 15807 8789
rect 16206 8780 16212 8832
rect 16264 8780 16270 8832
rect 16577 8823 16635 8829
rect 16577 8789 16589 8823
rect 16623 8820 16635 8823
rect 16850 8820 16856 8832
rect 16623 8792 16856 8820
rect 16623 8789 16635 8792
rect 16577 8783 16635 8789
rect 16850 8780 16856 8792
rect 16908 8820 16914 8832
rect 17218 8820 17224 8832
rect 16908 8792 17224 8820
rect 16908 8780 16914 8792
rect 17218 8780 17224 8792
rect 17276 8780 17282 8832
rect 17586 8780 17592 8832
rect 17644 8820 17650 8832
rect 19334 8820 19340 8832
rect 17644 8792 19340 8820
rect 17644 8780 17650 8792
rect 19334 8780 19340 8792
rect 19392 8780 19398 8832
rect 20622 8780 20628 8832
rect 20680 8780 20686 8832
rect 1104 8730 22976 8752
rect 1104 8678 6378 8730
rect 6430 8678 6442 8730
rect 6494 8678 6506 8730
rect 6558 8678 6570 8730
rect 6622 8678 6634 8730
rect 6686 8678 11806 8730
rect 11858 8678 11870 8730
rect 11922 8678 11934 8730
rect 11986 8678 11998 8730
rect 12050 8678 12062 8730
rect 12114 8678 17234 8730
rect 17286 8678 17298 8730
rect 17350 8678 17362 8730
rect 17414 8678 17426 8730
rect 17478 8678 17490 8730
rect 17542 8678 22662 8730
rect 22714 8678 22726 8730
rect 22778 8678 22790 8730
rect 22842 8678 22854 8730
rect 22906 8678 22918 8730
rect 22970 8678 22976 8730
rect 1104 8656 22976 8678
rect 4338 8576 4344 8628
rect 4396 8576 4402 8628
rect 8018 8576 8024 8628
rect 8076 8576 8082 8628
rect 10778 8576 10784 8628
rect 10836 8616 10842 8628
rect 10873 8619 10931 8625
rect 10873 8616 10885 8619
rect 10836 8588 10885 8616
rect 10836 8576 10842 8588
rect 10873 8585 10885 8588
rect 10919 8585 10931 8619
rect 10873 8579 10931 8585
rect 12802 8576 12808 8628
rect 12860 8576 12866 8628
rect 13354 8576 13360 8628
rect 13412 8576 13418 8628
rect 15286 8576 15292 8628
rect 15344 8576 15350 8628
rect 17586 8616 17592 8628
rect 15396 8588 17592 8616
rect 4798 8508 4804 8560
rect 4856 8548 4862 8560
rect 5454 8551 5512 8557
rect 5454 8548 5466 8551
rect 4856 8520 5466 8548
rect 4856 8508 4862 8520
rect 5454 8517 5466 8520
rect 5500 8517 5512 8551
rect 5454 8511 5512 8517
rect 6908 8551 6966 8557
rect 6908 8517 6920 8551
rect 6954 8548 6966 8551
rect 7282 8548 7288 8560
rect 6954 8520 7288 8548
rect 6954 8517 6966 8520
rect 6908 8511 6966 8517
rect 7282 8508 7288 8520
rect 7340 8508 7346 8560
rect 15304 8548 15332 8576
rect 15120 8520 15332 8548
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8480 5779 8483
rect 6641 8483 6699 8489
rect 6641 8480 6653 8483
rect 5767 8452 6653 8480
rect 5767 8449 5779 8452
rect 5721 8443 5779 8449
rect 6641 8449 6653 8452
rect 6687 8480 6699 8483
rect 6730 8480 6736 8492
rect 6687 8452 6736 8480
rect 6687 8449 6699 8452
rect 6641 8443 6699 8449
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 9490 8440 9496 8492
rect 9548 8440 9554 8492
rect 9769 8483 9827 8489
rect 9769 8449 9781 8483
rect 9815 8480 9827 8483
rect 11238 8480 11244 8492
rect 9815 8452 11244 8480
rect 9815 8449 9827 8452
rect 9769 8443 9827 8449
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 12250 8440 12256 8492
rect 12308 8480 12314 8492
rect 12713 8483 12771 8489
rect 12713 8480 12725 8483
rect 12308 8452 12725 8480
rect 12308 8440 12314 8452
rect 12713 8449 12725 8452
rect 12759 8449 12771 8483
rect 12713 8443 12771 8449
rect 13633 8483 13691 8489
rect 13633 8449 13645 8483
rect 13679 8480 13691 8483
rect 13722 8480 13728 8492
rect 13679 8452 13728 8480
rect 13679 8449 13691 8452
rect 13633 8443 13691 8449
rect 13722 8440 13728 8452
rect 13780 8480 13786 8492
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 13780 8452 14657 8480
rect 13780 8440 13786 8452
rect 14645 8449 14657 8452
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 14830 8483 14888 8489
rect 14830 8449 14842 8483
rect 14876 8449 14888 8483
rect 14830 8443 14888 8449
rect 14921 8483 14979 8489
rect 14921 8449 14933 8483
rect 14967 8480 14979 8483
rect 15120 8480 15148 8520
rect 15396 8492 15424 8588
rect 17586 8576 17592 8588
rect 17644 8576 17650 8628
rect 17865 8619 17923 8625
rect 17865 8585 17877 8619
rect 17911 8616 17923 8619
rect 18046 8616 18052 8628
rect 17911 8588 18052 8616
rect 17911 8585 17923 8588
rect 17865 8579 17923 8585
rect 18046 8576 18052 8588
rect 18104 8576 18110 8628
rect 19518 8576 19524 8628
rect 19576 8576 19582 8628
rect 20438 8576 20444 8628
rect 20496 8576 20502 8628
rect 15746 8508 15752 8560
rect 15804 8548 15810 8560
rect 15804 8520 15976 8548
rect 15804 8508 15810 8520
rect 14967 8452 15148 8480
rect 15197 8483 15255 8489
rect 14967 8449 14979 8452
rect 14921 8443 14979 8449
rect 15197 8449 15209 8483
rect 15243 8480 15255 8483
rect 15378 8480 15384 8492
rect 15243 8452 15384 8480
rect 15243 8449 15255 8452
rect 15197 8443 15255 8449
rect 13538 8372 13544 8424
rect 13596 8372 13602 8424
rect 13906 8372 13912 8424
rect 13964 8372 13970 8424
rect 14001 8415 14059 8421
rect 14001 8381 14013 8415
rect 14047 8412 14059 8415
rect 14182 8412 14188 8424
rect 14047 8384 14188 8412
rect 14047 8381 14059 8384
rect 14001 8375 14059 8381
rect 14182 8372 14188 8384
rect 14240 8372 14246 8424
rect 14844 8412 14872 8443
rect 15378 8440 15384 8452
rect 15436 8440 15442 8492
rect 15838 8440 15844 8492
rect 15896 8440 15902 8492
rect 15948 8489 15976 8520
rect 16482 8508 16488 8560
rect 16540 8548 16546 8560
rect 20609 8551 20667 8557
rect 16540 8520 20576 8548
rect 16540 8508 16546 8520
rect 15933 8483 15991 8489
rect 15933 8449 15945 8483
rect 15979 8449 15991 8483
rect 15933 8443 15991 8449
rect 16850 8440 16856 8492
rect 16908 8440 16914 8492
rect 17052 8489 17080 8520
rect 17037 8483 17095 8489
rect 17037 8449 17049 8483
rect 17083 8449 17095 8483
rect 17037 8443 17095 8449
rect 17494 8440 17500 8492
rect 17552 8440 17558 8492
rect 17678 8440 17684 8492
rect 17736 8480 17742 8492
rect 18877 8483 18935 8489
rect 18877 8480 18889 8483
rect 17736 8452 18889 8480
rect 17736 8440 17742 8452
rect 18877 8449 18889 8452
rect 18923 8449 18935 8483
rect 18877 8443 18935 8449
rect 19061 8483 19119 8489
rect 19061 8449 19073 8483
rect 19107 8449 19119 8483
rect 19061 8443 19119 8449
rect 15102 8412 15108 8424
rect 14844 8384 15108 8412
rect 15102 8372 15108 8384
rect 15160 8372 15166 8424
rect 15470 8372 15476 8424
rect 15528 8412 15534 8424
rect 16868 8412 16896 8440
rect 15528 8384 16896 8412
rect 15528 8372 15534 8384
rect 16942 8372 16948 8424
rect 17000 8372 17006 8424
rect 17402 8372 17408 8424
rect 17460 8412 17466 8424
rect 17589 8415 17647 8421
rect 17589 8412 17601 8415
rect 17460 8384 17601 8412
rect 17460 8372 17466 8384
rect 17589 8381 17601 8384
rect 17635 8381 17647 8415
rect 19076 8412 19104 8443
rect 19150 8440 19156 8492
rect 19208 8440 19214 8492
rect 19245 8483 19303 8489
rect 19245 8449 19257 8483
rect 19291 8480 19303 8483
rect 19334 8480 19340 8492
rect 19291 8452 19340 8480
rect 19291 8449 19303 8452
rect 19245 8443 19303 8449
rect 19334 8440 19340 8452
rect 19392 8440 19398 8492
rect 17589 8375 17647 8381
rect 17972 8384 19104 8412
rect 19168 8412 19196 8440
rect 20548 8424 20576 8520
rect 20609 8517 20621 8551
rect 20655 8548 20667 8551
rect 20714 8548 20720 8560
rect 20655 8520 20720 8548
rect 20655 8517 20667 8520
rect 20609 8511 20667 8517
rect 20714 8508 20720 8520
rect 20772 8508 20778 8560
rect 20806 8508 20812 8560
rect 20864 8508 20870 8560
rect 19702 8412 19708 8424
rect 19168 8384 19708 8412
rect 17972 8356 18000 8384
rect 19702 8372 19708 8384
rect 19760 8372 19766 8424
rect 20530 8372 20536 8424
rect 20588 8372 20594 8424
rect 17954 8304 17960 8356
rect 18012 8304 18018 8356
rect 14918 8236 14924 8288
rect 14976 8276 14982 8288
rect 15105 8279 15163 8285
rect 15105 8276 15117 8279
rect 14976 8248 15117 8276
rect 14976 8236 14982 8248
rect 15105 8245 15117 8248
rect 15151 8276 15163 8279
rect 15746 8276 15752 8288
rect 15151 8248 15752 8276
rect 15151 8245 15163 8248
rect 15105 8239 15163 8245
rect 15746 8236 15752 8248
rect 15804 8236 15810 8288
rect 15930 8236 15936 8288
rect 15988 8236 15994 8288
rect 17586 8236 17592 8288
rect 17644 8236 17650 8288
rect 20530 8236 20536 8288
rect 20588 8276 20594 8288
rect 20625 8279 20683 8285
rect 20625 8276 20637 8279
rect 20588 8248 20637 8276
rect 20588 8236 20594 8248
rect 20625 8245 20637 8248
rect 20671 8245 20683 8279
rect 20625 8239 20683 8245
rect 1104 8186 22816 8208
rect 1104 8134 3664 8186
rect 3716 8134 3728 8186
rect 3780 8134 3792 8186
rect 3844 8134 3856 8186
rect 3908 8134 3920 8186
rect 3972 8134 9092 8186
rect 9144 8134 9156 8186
rect 9208 8134 9220 8186
rect 9272 8134 9284 8186
rect 9336 8134 9348 8186
rect 9400 8134 14520 8186
rect 14572 8134 14584 8186
rect 14636 8134 14648 8186
rect 14700 8134 14712 8186
rect 14764 8134 14776 8186
rect 14828 8134 19948 8186
rect 20000 8134 20012 8186
rect 20064 8134 20076 8186
rect 20128 8134 20140 8186
rect 20192 8134 20204 8186
rect 20256 8134 22816 8186
rect 1104 8112 22816 8134
rect 10965 8075 11023 8081
rect 10965 8041 10977 8075
rect 11011 8072 11023 8075
rect 13446 8072 13452 8084
rect 11011 8044 13452 8072
rect 11011 8041 11023 8044
rect 10965 8035 11023 8041
rect 13446 8032 13452 8044
rect 13504 8032 13510 8084
rect 14921 8075 14979 8081
rect 14921 8041 14933 8075
rect 14967 8072 14979 8075
rect 15102 8072 15108 8084
rect 14967 8044 15108 8072
rect 14967 8041 14979 8044
rect 14921 8035 14979 8041
rect 15102 8032 15108 8044
rect 15160 8072 15166 8084
rect 15470 8072 15476 8084
rect 15160 8044 15476 8072
rect 15160 8032 15166 8044
rect 15470 8032 15476 8044
rect 15528 8032 15534 8084
rect 15746 8032 15752 8084
rect 15804 8072 15810 8084
rect 17310 8072 17316 8084
rect 15804 8044 17316 8072
rect 15804 8032 15810 8044
rect 17310 8032 17316 8044
rect 17368 8032 17374 8084
rect 17405 8075 17463 8081
rect 17405 8041 17417 8075
rect 17451 8072 17463 8075
rect 17586 8072 17592 8084
rect 17451 8044 17592 8072
rect 17451 8041 17463 8044
rect 17405 8035 17463 8041
rect 17586 8032 17592 8044
rect 17644 8032 17650 8084
rect 19426 8032 19432 8084
rect 19484 8072 19490 8084
rect 19797 8075 19855 8081
rect 19797 8072 19809 8075
rect 19484 8044 19809 8072
rect 19484 8032 19490 8044
rect 19797 8041 19809 8044
rect 19843 8041 19855 8075
rect 19797 8035 19855 8041
rect 12618 7964 12624 8016
rect 12676 8004 12682 8016
rect 13354 8004 13360 8016
rect 12676 7976 13360 8004
rect 12676 7964 12682 7976
rect 13354 7964 13360 7976
rect 13412 7964 13418 8016
rect 16206 7964 16212 8016
rect 16264 8004 16270 8016
rect 17037 8007 17095 8013
rect 17037 8004 17049 8007
rect 16264 7976 17049 8004
rect 16264 7964 16270 7976
rect 17037 7973 17049 7976
rect 17083 7973 17095 8007
rect 17328 8004 17356 8032
rect 20990 8004 20996 8016
rect 17328 7976 20996 8004
rect 17037 7967 17095 7973
rect 9490 7896 9496 7948
rect 9548 7936 9554 7948
rect 9585 7939 9643 7945
rect 9585 7936 9597 7939
rect 9548 7908 9597 7936
rect 9548 7896 9554 7908
rect 9585 7905 9597 7908
rect 9631 7905 9643 7939
rect 14918 7936 14924 7948
rect 9585 7899 9643 7905
rect 12912 7908 14924 7936
rect 2222 7828 2228 7880
rect 2280 7868 2286 7880
rect 2317 7871 2375 7877
rect 2317 7868 2329 7871
rect 2280 7840 2329 7868
rect 2280 7828 2286 7840
rect 2317 7837 2329 7840
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 2332 7800 2360 7831
rect 2498 7828 2504 7880
rect 2556 7828 2562 7880
rect 12158 7828 12164 7880
rect 12216 7868 12222 7880
rect 12912 7877 12940 7908
rect 14918 7896 14924 7908
rect 14976 7936 14982 7948
rect 14976 7908 15148 7936
rect 14976 7896 14982 7908
rect 12897 7871 12955 7877
rect 12897 7868 12909 7871
rect 12216 7840 12909 7868
rect 12216 7828 12222 7840
rect 12897 7837 12909 7840
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 13262 7828 13268 7880
rect 13320 7828 13326 7880
rect 13354 7828 13360 7880
rect 13412 7828 13418 7880
rect 15120 7877 15148 7908
rect 15286 7896 15292 7948
rect 15344 7936 15350 7948
rect 15838 7936 15844 7948
rect 15344 7908 15844 7936
rect 15344 7896 15350 7908
rect 15838 7896 15844 7908
rect 15896 7896 15902 7948
rect 16942 7896 16948 7948
rect 17000 7936 17006 7948
rect 17402 7936 17408 7948
rect 17000 7908 17408 7936
rect 17000 7896 17006 7908
rect 17402 7896 17408 7908
rect 17460 7896 17466 7948
rect 20625 7939 20683 7945
rect 20625 7936 20637 7939
rect 20088 7908 20637 7936
rect 20088 7877 20116 7908
rect 20625 7905 20637 7908
rect 20671 7905 20683 7939
rect 20625 7899 20683 7905
rect 15105 7871 15163 7877
rect 15105 7837 15117 7871
rect 15151 7837 15163 7871
rect 15105 7831 15163 7837
rect 20073 7871 20131 7877
rect 20073 7837 20085 7871
rect 20119 7837 20131 7871
rect 20073 7831 20131 7837
rect 20346 7828 20352 7880
rect 20404 7868 20410 7880
rect 20732 7877 20760 7976
rect 20990 7964 20996 7976
rect 21048 7964 21054 8016
rect 20533 7871 20591 7877
rect 20533 7868 20545 7871
rect 20404 7840 20545 7868
rect 20404 7828 20410 7840
rect 20533 7837 20545 7840
rect 20579 7837 20591 7871
rect 20533 7831 20591 7837
rect 20717 7871 20775 7877
rect 20717 7837 20729 7871
rect 20763 7837 20775 7871
rect 20717 7831 20775 7837
rect 2682 7800 2688 7812
rect 2332 7772 2688 7800
rect 2682 7760 2688 7772
rect 2740 7760 2746 7812
rect 5534 7760 5540 7812
rect 5592 7800 5598 7812
rect 5721 7803 5779 7809
rect 5721 7800 5733 7803
rect 5592 7772 5733 7800
rect 5592 7760 5598 7772
rect 5721 7769 5733 7772
rect 5767 7769 5779 7803
rect 7469 7803 7527 7809
rect 7469 7800 7481 7803
rect 5721 7763 5779 7769
rect 6886 7772 7481 7800
rect 2406 7692 2412 7744
rect 2464 7692 2470 7744
rect 4338 7692 4344 7744
rect 4396 7732 4402 7744
rect 6886 7732 6914 7772
rect 7469 7769 7481 7772
rect 7515 7800 7527 7803
rect 7834 7800 7840 7812
rect 7515 7772 7840 7800
rect 7515 7769 7527 7772
rect 7469 7763 7527 7769
rect 7834 7760 7840 7772
rect 7892 7760 7898 7812
rect 9852 7803 9910 7809
rect 9852 7769 9864 7803
rect 9898 7800 9910 7803
rect 12342 7800 12348 7812
rect 9898 7772 12348 7800
rect 9898 7769 9910 7772
rect 9852 7763 9910 7769
rect 12342 7760 12348 7772
rect 12400 7760 12406 7812
rect 12802 7760 12808 7812
rect 12860 7800 12866 7812
rect 13081 7803 13139 7809
rect 13081 7800 13093 7803
rect 12860 7772 13093 7800
rect 12860 7760 12866 7772
rect 13081 7769 13093 7772
rect 13127 7769 13139 7803
rect 13081 7763 13139 7769
rect 19797 7803 19855 7809
rect 19797 7769 19809 7803
rect 19843 7800 19855 7803
rect 20438 7800 20444 7812
rect 19843 7772 20444 7800
rect 19843 7769 19855 7772
rect 19797 7763 19855 7769
rect 20438 7760 20444 7772
rect 20496 7760 20502 7812
rect 4396 7704 6914 7732
rect 12621 7735 12679 7741
rect 4396 7692 4402 7704
rect 12621 7701 12633 7735
rect 12667 7732 12679 7735
rect 12894 7732 12900 7744
rect 12667 7704 12900 7732
rect 12667 7701 12679 7704
rect 12621 7695 12679 7701
rect 12894 7692 12900 7704
rect 12952 7692 12958 7744
rect 12989 7735 13047 7741
rect 12989 7701 13001 7735
rect 13035 7732 13047 7735
rect 13446 7732 13452 7744
rect 13035 7704 13452 7732
rect 13035 7701 13047 7704
rect 12989 7695 13047 7701
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 15102 7692 15108 7744
rect 15160 7732 15166 7744
rect 17405 7735 17463 7741
rect 17405 7732 17417 7735
rect 15160 7704 17417 7732
rect 15160 7692 15166 7704
rect 17405 7701 17417 7704
rect 17451 7701 17463 7735
rect 17405 7695 17463 7701
rect 17589 7735 17647 7741
rect 17589 7701 17601 7735
rect 17635 7732 17647 7735
rect 18138 7732 18144 7744
rect 17635 7704 18144 7732
rect 17635 7701 17647 7704
rect 17589 7695 17647 7701
rect 18138 7692 18144 7704
rect 18196 7692 18202 7744
rect 19702 7692 19708 7744
rect 19760 7732 19766 7744
rect 19981 7735 20039 7741
rect 19981 7732 19993 7735
rect 19760 7704 19993 7732
rect 19760 7692 19766 7704
rect 19981 7701 19993 7704
rect 20027 7701 20039 7735
rect 19981 7695 20039 7701
rect 1104 7642 22976 7664
rect 1104 7590 6378 7642
rect 6430 7590 6442 7642
rect 6494 7590 6506 7642
rect 6558 7590 6570 7642
rect 6622 7590 6634 7642
rect 6686 7590 11806 7642
rect 11858 7590 11870 7642
rect 11922 7590 11934 7642
rect 11986 7590 11998 7642
rect 12050 7590 12062 7642
rect 12114 7590 17234 7642
rect 17286 7590 17298 7642
rect 17350 7590 17362 7642
rect 17414 7590 17426 7642
rect 17478 7590 17490 7642
rect 17542 7590 22662 7642
rect 22714 7590 22726 7642
rect 22778 7590 22790 7642
rect 22842 7590 22854 7642
rect 22906 7590 22918 7642
rect 22970 7590 22976 7642
rect 1104 7568 22976 7590
rect 2866 7488 2872 7540
rect 2924 7488 2930 7540
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 13446 7528 13452 7540
rect 12492 7500 13452 7528
rect 12492 7488 12498 7500
rect 13446 7488 13452 7500
rect 13504 7488 13510 7540
rect 17586 7488 17592 7540
rect 17644 7528 17650 7540
rect 19242 7528 19248 7540
rect 17644 7500 19248 7528
rect 17644 7488 17650 7500
rect 19242 7488 19248 7500
rect 19300 7488 19306 7540
rect 19334 7488 19340 7540
rect 19392 7528 19398 7540
rect 19797 7531 19855 7537
rect 19797 7528 19809 7531
rect 19392 7500 19809 7528
rect 19392 7488 19398 7500
rect 19797 7497 19809 7500
rect 19843 7528 19855 7531
rect 20346 7528 20352 7540
rect 19843 7500 20352 7528
rect 19843 7497 19855 7500
rect 19797 7491 19855 7497
rect 20346 7488 20352 7500
rect 20404 7488 20410 7540
rect 4338 7420 4344 7472
rect 4396 7420 4402 7472
rect 8938 7420 8944 7472
rect 8996 7460 9002 7472
rect 9490 7460 9496 7472
rect 8996 7432 9496 7460
rect 8996 7420 9002 7432
rect 9490 7420 9496 7432
rect 9548 7420 9554 7472
rect 11698 7420 11704 7472
rect 11756 7460 11762 7472
rect 15378 7460 15384 7472
rect 11756 7432 15384 7460
rect 11756 7420 11762 7432
rect 15378 7420 15384 7432
rect 15436 7420 15442 7472
rect 17862 7420 17868 7472
rect 17920 7420 17926 7472
rect 20714 7460 20720 7472
rect 20364 7432 20720 7460
rect 7834 7352 7840 7404
rect 7892 7352 7898 7404
rect 12342 7352 12348 7404
rect 12400 7392 12406 7404
rect 12713 7395 12771 7401
rect 12713 7392 12725 7395
rect 12400 7364 12725 7392
rect 12400 7352 12406 7364
rect 12713 7361 12725 7364
rect 12759 7361 12771 7395
rect 12713 7355 12771 7361
rect 12894 7352 12900 7404
rect 12952 7352 12958 7404
rect 12986 7352 12992 7404
rect 13044 7352 13050 7404
rect 15105 7395 15163 7401
rect 15105 7361 15117 7395
rect 15151 7392 15163 7395
rect 15562 7392 15568 7404
rect 15151 7364 15568 7392
rect 15151 7361 15163 7364
rect 15105 7355 15163 7361
rect 15562 7352 15568 7364
rect 15620 7392 15626 7404
rect 17126 7392 17132 7404
rect 15620 7364 17132 7392
rect 15620 7352 15626 7364
rect 17126 7352 17132 7364
rect 17184 7352 17190 7404
rect 17681 7395 17739 7401
rect 17681 7361 17693 7395
rect 17727 7361 17739 7395
rect 17681 7355 17739 7361
rect 12805 7327 12863 7333
rect 12805 7293 12817 7327
rect 12851 7324 12863 7327
rect 15010 7324 15016 7336
rect 12851 7296 15016 7324
rect 12851 7293 12863 7296
rect 12805 7287 12863 7293
rect 15010 7284 15016 7296
rect 15068 7284 15074 7336
rect 16942 7284 16948 7336
rect 17000 7324 17006 7336
rect 17586 7324 17592 7336
rect 17000 7296 17592 7324
rect 17000 7284 17006 7296
rect 17586 7284 17592 7296
rect 17644 7324 17650 7336
rect 17696 7324 17724 7355
rect 19242 7352 19248 7404
rect 19300 7392 19306 7404
rect 20364 7401 20392 7432
rect 20714 7420 20720 7432
rect 20772 7420 20778 7472
rect 19705 7395 19763 7401
rect 19705 7392 19717 7395
rect 19300 7364 19717 7392
rect 19300 7352 19306 7364
rect 19705 7361 19717 7364
rect 19751 7361 19763 7395
rect 19705 7355 19763 7361
rect 20349 7395 20407 7401
rect 20349 7361 20361 7395
rect 20395 7361 20407 7395
rect 20349 7355 20407 7361
rect 20530 7352 20536 7404
rect 20588 7352 20594 7404
rect 17644 7296 17724 7324
rect 17644 7284 17650 7296
rect 12526 7148 12532 7200
rect 12584 7148 12590 7200
rect 14274 7148 14280 7200
rect 14332 7188 14338 7200
rect 15102 7188 15108 7200
rect 14332 7160 15108 7188
rect 14332 7148 14338 7160
rect 15102 7148 15108 7160
rect 15160 7188 15166 7200
rect 15197 7191 15255 7197
rect 15197 7188 15209 7191
rect 15160 7160 15209 7188
rect 15160 7148 15166 7160
rect 15197 7157 15209 7160
rect 15243 7157 15255 7191
rect 15197 7151 15255 7157
rect 20346 7148 20352 7200
rect 20404 7148 20410 7200
rect 1104 7098 22816 7120
rect 1104 7046 3664 7098
rect 3716 7046 3728 7098
rect 3780 7046 3792 7098
rect 3844 7046 3856 7098
rect 3908 7046 3920 7098
rect 3972 7046 9092 7098
rect 9144 7046 9156 7098
rect 9208 7046 9220 7098
rect 9272 7046 9284 7098
rect 9336 7046 9348 7098
rect 9400 7046 14520 7098
rect 14572 7046 14584 7098
rect 14636 7046 14648 7098
rect 14700 7046 14712 7098
rect 14764 7046 14776 7098
rect 14828 7046 19948 7098
rect 20000 7046 20012 7098
rect 20064 7046 20076 7098
rect 20128 7046 20140 7098
rect 20192 7046 20204 7098
rect 20256 7046 22816 7098
rect 1104 7024 22816 7046
rect 17497 6987 17555 6993
rect 17497 6953 17509 6987
rect 17543 6953 17555 6987
rect 17497 6947 17555 6953
rect 13262 6916 13268 6928
rect 12544 6888 13268 6916
rect 1670 6740 1676 6792
rect 1728 6740 1734 6792
rect 1940 6783 1998 6789
rect 1940 6749 1952 6783
rect 1986 6780 1998 6783
rect 2406 6780 2412 6792
rect 1986 6752 2412 6780
rect 1986 6749 1998 6752
rect 1940 6743 1998 6749
rect 2406 6740 2412 6752
rect 2464 6740 2470 6792
rect 3970 6740 3976 6792
rect 4028 6780 4034 6792
rect 5721 6783 5779 6789
rect 5721 6780 5733 6783
rect 4028 6752 5733 6780
rect 4028 6740 4034 6752
rect 5721 6749 5733 6752
rect 5767 6749 5779 6783
rect 5721 6743 5779 6749
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6780 6975 6783
rect 8938 6780 8944 6792
rect 6963 6752 8944 6780
rect 6963 6749 6975 6752
rect 6917 6743 6975 6749
rect 8938 6740 8944 6752
rect 8996 6740 9002 6792
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 9493 6783 9551 6789
rect 9493 6780 9505 6783
rect 9364 6752 9505 6780
rect 9364 6740 9370 6752
rect 9493 6749 9505 6752
rect 9539 6780 9551 6783
rect 11425 6783 11483 6789
rect 11425 6780 11437 6783
rect 9539 6752 11437 6780
rect 9539 6749 9551 6752
rect 9493 6743 9551 6749
rect 11425 6749 11437 6752
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 11692 6783 11750 6789
rect 11692 6749 11704 6783
rect 11738 6780 11750 6783
rect 12544 6780 12572 6888
rect 13262 6876 13268 6888
rect 13320 6876 13326 6928
rect 13446 6876 13452 6928
rect 13504 6916 13510 6928
rect 15746 6916 15752 6928
rect 13504 6888 15752 6916
rect 13504 6876 13510 6888
rect 15746 6876 15752 6888
rect 15804 6876 15810 6928
rect 17512 6860 17540 6947
rect 17862 6944 17868 6996
rect 17920 6984 17926 6996
rect 18417 6987 18475 6993
rect 18417 6984 18429 6987
rect 17920 6956 18429 6984
rect 17920 6944 17926 6956
rect 18417 6953 18429 6956
rect 18463 6953 18475 6987
rect 19794 6984 19800 6996
rect 18417 6947 18475 6953
rect 19536 6956 19800 6984
rect 18785 6919 18843 6925
rect 17604 6888 17908 6916
rect 17604 6860 17632 6888
rect 13078 6808 13084 6860
rect 13136 6848 13142 6860
rect 13541 6851 13599 6857
rect 13541 6848 13553 6851
rect 13136 6820 13553 6848
rect 13136 6808 13142 6820
rect 13541 6817 13553 6820
rect 13587 6817 13599 6851
rect 13541 6811 13599 6817
rect 13906 6808 13912 6860
rect 13964 6848 13970 6860
rect 14277 6851 14335 6857
rect 14277 6848 14289 6851
rect 13964 6820 14289 6848
rect 13964 6808 13970 6820
rect 14277 6817 14289 6820
rect 14323 6817 14335 6851
rect 14277 6811 14335 6817
rect 15194 6808 15200 6860
rect 15252 6808 15258 6860
rect 16301 6851 16359 6857
rect 16301 6817 16313 6851
rect 16347 6848 16359 6851
rect 16482 6848 16488 6860
rect 16347 6820 16488 6848
rect 16347 6817 16359 6820
rect 16301 6811 16359 6817
rect 16482 6808 16488 6820
rect 16540 6808 16546 6860
rect 17494 6808 17500 6860
rect 17552 6808 17558 6860
rect 17586 6808 17592 6860
rect 17644 6808 17650 6860
rect 17678 6808 17684 6860
rect 17736 6808 17742 6860
rect 17880 6848 17908 6888
rect 18785 6885 18797 6919
rect 18831 6885 18843 6919
rect 18785 6879 18843 6885
rect 18509 6851 18567 6857
rect 18509 6848 18521 6851
rect 17880 6820 18521 6848
rect 18509 6817 18521 6820
rect 18555 6817 18567 6851
rect 18800 6848 18828 6879
rect 19536 6848 19564 6956
rect 19794 6944 19800 6956
rect 19852 6944 19858 6996
rect 19610 6876 19616 6928
rect 19668 6876 19674 6928
rect 18800 6820 19564 6848
rect 19628 6848 19656 6876
rect 19797 6851 19855 6857
rect 19797 6848 19809 6851
rect 19628 6820 19809 6848
rect 18509 6811 18567 6817
rect 19797 6817 19809 6820
rect 19843 6817 19855 6851
rect 19797 6811 19855 6817
rect 19889 6851 19947 6857
rect 19889 6817 19901 6851
rect 19935 6848 19947 6851
rect 20622 6848 20628 6860
rect 19935 6820 20628 6848
rect 19935 6817 19947 6820
rect 19889 6811 19947 6817
rect 20622 6808 20628 6820
rect 20680 6808 20686 6860
rect 11738 6752 12572 6780
rect 11738 6749 11750 6752
rect 11692 6743 11750 6749
rect 12618 6740 12624 6792
rect 12676 6780 12682 6792
rect 13265 6783 13323 6789
rect 13265 6780 13277 6783
rect 12676 6752 13277 6780
rect 12676 6740 12682 6752
rect 13265 6749 13277 6752
rect 13311 6749 13323 6783
rect 13265 6743 13323 6749
rect 13354 6740 13360 6792
rect 13412 6740 13418 6792
rect 15105 6783 15163 6789
rect 15105 6749 15117 6783
rect 15151 6780 15163 6783
rect 15286 6780 15292 6792
rect 15151 6752 15292 6780
rect 15151 6749 15163 6752
rect 15105 6743 15163 6749
rect 15286 6740 15292 6752
rect 15344 6740 15350 6792
rect 16577 6783 16635 6789
rect 16577 6749 16589 6783
rect 16623 6780 16635 6783
rect 17034 6780 17040 6792
rect 16623 6752 17040 6780
rect 16623 6749 16635 6752
rect 16577 6743 16635 6749
rect 17034 6740 17040 6752
rect 17092 6780 17098 6792
rect 17368 6783 17426 6789
rect 17368 6780 17380 6783
rect 17092 6752 17380 6780
rect 17092 6740 17098 6752
rect 17368 6749 17380 6752
rect 17414 6749 17426 6783
rect 17512 6780 17540 6808
rect 18417 6783 18475 6789
rect 18417 6780 18429 6783
rect 17512 6752 18429 6780
rect 17368 6743 17426 6749
rect 18417 6749 18429 6752
rect 18463 6749 18475 6783
rect 18417 6743 18475 6749
rect 19610 6740 19616 6792
rect 19668 6740 19674 6792
rect 19705 6783 19763 6789
rect 19705 6749 19717 6783
rect 19751 6749 19763 6783
rect 19705 6743 19763 6749
rect 5442 6672 5448 6724
rect 5500 6721 5506 6724
rect 9766 6721 9772 6724
rect 5500 6675 5512 6721
rect 7184 6715 7242 6721
rect 7184 6681 7196 6715
rect 7230 6712 7242 6715
rect 7230 6684 9720 6712
rect 7230 6681 7242 6684
rect 7184 6675 7242 6681
rect 5500 6672 5506 6675
rect 2498 6604 2504 6656
rect 2556 6644 2562 6656
rect 3053 6647 3111 6653
rect 3053 6644 3065 6647
rect 2556 6616 3065 6644
rect 2556 6604 2562 6616
rect 3053 6613 3065 6616
rect 3099 6613 3111 6647
rect 3053 6607 3111 6613
rect 4341 6647 4399 6653
rect 4341 6613 4353 6647
rect 4387 6644 4399 6647
rect 4982 6644 4988 6656
rect 4387 6616 4988 6644
rect 4387 6613 4399 6616
rect 4341 6607 4399 6613
rect 4982 6604 4988 6616
rect 5040 6604 5046 6656
rect 8294 6604 8300 6656
rect 8352 6604 8358 6656
rect 9692 6644 9720 6684
rect 9760 6675 9772 6721
rect 9766 6672 9772 6675
rect 9824 6672 9830 6724
rect 12710 6712 12716 6724
rect 10796 6684 12716 6712
rect 10796 6644 10824 6684
rect 12710 6672 12716 6684
rect 12768 6672 12774 6724
rect 12820 6684 13492 6712
rect 9692 6616 10824 6644
rect 10873 6647 10931 6653
rect 10873 6613 10885 6647
rect 10919 6644 10931 6647
rect 12434 6644 12440 6656
rect 10919 6616 12440 6644
rect 10919 6613 10931 6616
rect 10873 6607 10931 6613
rect 12434 6604 12440 6616
rect 12492 6604 12498 6656
rect 12820 6653 12848 6684
rect 12805 6647 12863 6653
rect 12805 6613 12817 6647
rect 12851 6613 12863 6647
rect 12805 6607 12863 6613
rect 13262 6604 13268 6656
rect 13320 6604 13326 6656
rect 13464 6644 13492 6684
rect 16758 6672 16764 6724
rect 16816 6712 16822 6724
rect 17221 6715 17279 6721
rect 17221 6712 17233 6715
rect 16816 6684 17233 6712
rect 16816 6672 16822 6684
rect 17221 6681 17233 6684
rect 17267 6681 17279 6715
rect 17221 6675 17279 6681
rect 18598 6672 18604 6724
rect 18656 6712 18662 6724
rect 19720 6712 19748 6743
rect 18656 6684 19748 6712
rect 18656 6672 18662 6684
rect 16022 6644 16028 6656
rect 13464 6616 16028 6644
rect 16022 6604 16028 6616
rect 16080 6604 16086 6656
rect 19426 6604 19432 6656
rect 19484 6604 19490 6656
rect 1104 6554 22976 6576
rect 1104 6502 6378 6554
rect 6430 6502 6442 6554
rect 6494 6502 6506 6554
rect 6558 6502 6570 6554
rect 6622 6502 6634 6554
rect 6686 6502 11806 6554
rect 11858 6502 11870 6554
rect 11922 6502 11934 6554
rect 11986 6502 11998 6554
rect 12050 6502 12062 6554
rect 12114 6502 17234 6554
rect 17286 6502 17298 6554
rect 17350 6502 17362 6554
rect 17414 6502 17426 6554
rect 17478 6502 17490 6554
rect 17542 6502 22662 6554
rect 22714 6502 22726 6554
rect 22778 6502 22790 6554
rect 22842 6502 22854 6554
rect 22906 6502 22918 6554
rect 22970 6502 22976 6554
rect 1104 6480 22976 6502
rect 3142 6400 3148 6452
rect 3200 6400 3206 6452
rect 12636 6412 15332 6440
rect 1670 6332 1676 6384
rect 1728 6372 1734 6384
rect 10965 6375 11023 6381
rect 1728 6344 3188 6372
rect 1728 6332 1734 6344
rect 1780 6313 1808 6344
rect 3160 6316 3188 6344
rect 10965 6341 10977 6375
rect 11011 6372 11023 6375
rect 12250 6372 12256 6384
rect 11011 6344 12256 6372
rect 11011 6341 11023 6344
rect 10965 6335 11023 6341
rect 12250 6332 12256 6344
rect 12308 6372 12314 6384
rect 12636 6372 12664 6412
rect 15304 6384 15332 6412
rect 16942 6400 16948 6452
rect 17000 6440 17006 6452
rect 17000 6412 17080 6440
rect 17000 6400 17006 6412
rect 12308 6344 12664 6372
rect 12308 6332 12314 6344
rect 15286 6332 15292 6384
rect 15344 6372 15350 6384
rect 17052 6372 17080 6412
rect 17126 6400 17132 6452
rect 17184 6440 17190 6452
rect 17405 6443 17463 6449
rect 17405 6440 17417 6443
rect 17184 6412 17417 6440
rect 17184 6400 17190 6412
rect 17405 6409 17417 6412
rect 17451 6409 17463 6443
rect 17405 6403 17463 6409
rect 18509 6443 18567 6449
rect 18509 6409 18521 6443
rect 18555 6440 18567 6443
rect 18598 6440 18604 6452
rect 18555 6412 18604 6440
rect 18555 6409 18567 6412
rect 18509 6403 18567 6409
rect 18598 6400 18604 6412
rect 18656 6400 18662 6452
rect 19610 6400 19616 6452
rect 19668 6440 19674 6452
rect 19705 6443 19763 6449
rect 19705 6440 19717 6443
rect 19668 6412 19717 6440
rect 19668 6400 19674 6412
rect 19705 6409 19717 6412
rect 19751 6409 19763 6443
rect 19705 6403 19763 6409
rect 15344 6344 15884 6372
rect 17052 6344 17172 6372
rect 15344 6332 15350 6344
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6273 1823 6307
rect 1765 6267 1823 6273
rect 2032 6307 2090 6313
rect 2032 6273 2044 6307
rect 2078 6304 2090 6307
rect 2958 6304 2964 6316
rect 2078 6276 2964 6304
rect 2078 6273 2090 6276
rect 2032 6267 2090 6273
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 3142 6264 3148 6316
rect 3200 6304 3206 6316
rect 3970 6304 3976 6316
rect 3200 6276 3976 6304
rect 3200 6264 3206 6276
rect 3970 6264 3976 6276
rect 4028 6264 4034 6316
rect 6816 6307 6874 6313
rect 6816 6273 6828 6307
rect 6862 6304 6874 6307
rect 6862 6276 9260 6304
rect 6862 6273 6874 6276
rect 6816 6267 6874 6273
rect 4249 6239 4307 6245
rect 4249 6236 4261 6239
rect 2792 6208 4261 6236
rect 2682 6060 2688 6112
rect 2740 6100 2746 6112
rect 2792 6100 2820 6208
rect 4249 6205 4261 6208
rect 4295 6205 4307 6239
rect 4249 6199 4307 6205
rect 6546 6196 6552 6248
rect 6604 6196 6610 6248
rect 9232 6236 9260 6276
rect 9306 6264 9312 6316
rect 9364 6264 9370 6316
rect 9585 6307 9643 6313
rect 9585 6273 9597 6307
rect 9631 6304 9643 6307
rect 11698 6304 11704 6316
rect 9631 6276 11704 6304
rect 9631 6273 9643 6276
rect 9585 6267 9643 6273
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 12802 6264 12808 6316
rect 12860 6264 12866 6316
rect 13078 6264 13084 6316
rect 13136 6264 13142 6316
rect 13265 6307 13323 6313
rect 13265 6273 13277 6307
rect 13311 6273 13323 6307
rect 13265 6267 13323 6273
rect 12526 6236 12532 6248
rect 9232 6208 12532 6236
rect 12526 6196 12532 6208
rect 12584 6196 12590 6248
rect 12618 6196 12624 6248
rect 12676 6196 12682 6248
rect 13280 6236 13308 6267
rect 13814 6264 13820 6316
rect 13872 6304 13878 6316
rect 13872 6276 13952 6304
rect 13872 6264 13878 6276
rect 13924 6236 13952 6276
rect 14090 6264 14096 6316
rect 14148 6304 14154 6316
rect 15102 6304 15108 6316
rect 14148 6276 15108 6304
rect 14148 6264 14154 6276
rect 15102 6264 15108 6276
rect 15160 6264 15166 6316
rect 15194 6264 15200 6316
rect 15252 6304 15258 6316
rect 15654 6304 15660 6316
rect 15252 6276 15660 6304
rect 15252 6264 15258 6276
rect 15654 6264 15660 6276
rect 15712 6264 15718 6316
rect 15856 6313 15884 6344
rect 17144 6316 17172 6344
rect 15841 6307 15899 6313
rect 15841 6273 15853 6307
rect 15887 6304 15899 6307
rect 15930 6304 15936 6316
rect 15887 6276 15936 6304
rect 15887 6273 15899 6276
rect 15841 6267 15899 6273
rect 15930 6264 15936 6276
rect 15988 6264 15994 6316
rect 16117 6307 16175 6313
rect 16117 6273 16129 6307
rect 16163 6304 16175 6307
rect 16758 6304 16764 6316
rect 16163 6276 16764 6304
rect 16163 6273 16175 6276
rect 16117 6267 16175 6273
rect 16758 6264 16764 6276
rect 16816 6304 16822 6316
rect 16945 6307 17003 6313
rect 16945 6304 16957 6307
rect 16816 6276 16957 6304
rect 16816 6264 16822 6276
rect 16945 6273 16957 6276
rect 16991 6273 17003 6307
rect 16945 6267 17003 6273
rect 17126 6264 17132 6316
rect 17184 6304 17190 6316
rect 17221 6307 17279 6313
rect 17221 6304 17233 6307
rect 17184 6276 17233 6304
rect 17184 6264 17190 6276
rect 17221 6273 17233 6276
rect 17267 6273 17279 6307
rect 17221 6267 17279 6273
rect 17770 6264 17776 6316
rect 17828 6304 17834 6316
rect 18141 6307 18199 6313
rect 18141 6304 18153 6307
rect 17828 6276 18153 6304
rect 17828 6264 17834 6276
rect 18141 6273 18153 6276
rect 18187 6273 18199 6307
rect 18141 6267 18199 6273
rect 18230 6264 18236 6316
rect 18288 6264 18294 6316
rect 19334 6264 19340 6316
rect 19392 6264 19398 6316
rect 19475 6307 19533 6313
rect 19475 6273 19487 6307
rect 19521 6304 19533 6307
rect 19702 6304 19708 6316
rect 19521 6276 19708 6304
rect 19521 6273 19533 6276
rect 19475 6267 19533 6273
rect 19702 6264 19708 6276
rect 19760 6264 19766 6316
rect 19797 6307 19855 6313
rect 19797 6273 19809 6307
rect 19843 6304 19855 6307
rect 20438 6304 20444 6316
rect 19843 6276 20444 6304
rect 19843 6273 19855 6276
rect 19797 6267 19855 6273
rect 20438 6264 20444 6276
rect 20496 6264 20502 6316
rect 14918 6236 14924 6248
rect 13280 6208 13860 6236
rect 13924 6208 14924 6236
rect 13832 6180 13860 6208
rect 14918 6196 14924 6208
rect 14976 6196 14982 6248
rect 15746 6196 15752 6248
rect 15804 6236 15810 6248
rect 16209 6239 16267 6245
rect 16209 6236 16221 6239
rect 15804 6208 16221 6236
rect 15804 6196 15810 6208
rect 16209 6205 16221 6208
rect 16255 6205 16267 6239
rect 16209 6199 16267 6205
rect 19613 6239 19671 6245
rect 19613 6205 19625 6239
rect 19659 6236 19671 6239
rect 20346 6236 20352 6248
rect 19659 6208 20352 6236
rect 19659 6205 19671 6208
rect 19613 6199 19671 6205
rect 20346 6196 20352 6208
rect 20404 6196 20410 6248
rect 13814 6128 13820 6180
rect 13872 6128 13878 6180
rect 17034 6128 17040 6180
rect 17092 6128 17098 6180
rect 2740 6072 2820 6100
rect 5537 6103 5595 6109
rect 2740 6060 2746 6072
rect 5537 6069 5549 6103
rect 5583 6100 5595 6103
rect 5626 6100 5632 6112
rect 5583 6072 5632 6100
rect 5583 6069 5595 6072
rect 5537 6063 5595 6069
rect 5626 6060 5632 6072
rect 5684 6060 5690 6112
rect 7929 6103 7987 6109
rect 7929 6069 7941 6103
rect 7975 6100 7987 6103
rect 8754 6100 8760 6112
rect 7975 6072 8760 6100
rect 7975 6069 7987 6072
rect 7929 6063 7987 6069
rect 8754 6060 8760 6072
rect 8812 6060 8818 6112
rect 18138 6060 18144 6112
rect 18196 6060 18202 6112
rect 1104 6010 22816 6032
rect 1104 5958 3664 6010
rect 3716 5958 3728 6010
rect 3780 5958 3792 6010
rect 3844 5958 3856 6010
rect 3908 5958 3920 6010
rect 3972 5958 9092 6010
rect 9144 5958 9156 6010
rect 9208 5958 9220 6010
rect 9272 5958 9284 6010
rect 9336 5958 9348 6010
rect 9400 5958 14520 6010
rect 14572 5958 14584 6010
rect 14636 5958 14648 6010
rect 14700 5958 14712 6010
rect 14764 5958 14776 6010
rect 14828 5958 19948 6010
rect 20000 5958 20012 6010
rect 20064 5958 20076 6010
rect 20128 5958 20140 6010
rect 20192 5958 20204 6010
rect 20256 5958 22816 6010
rect 1104 5936 22816 5958
rect 2406 5856 2412 5908
rect 2464 5896 2470 5908
rect 4341 5899 4399 5905
rect 4341 5896 4353 5899
rect 2464 5868 4353 5896
rect 2464 5856 2470 5868
rect 4341 5865 4353 5868
rect 4387 5896 4399 5899
rect 12802 5896 12808 5908
rect 4387 5868 12808 5896
rect 4387 5865 4399 5868
rect 4341 5859 4399 5865
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 13354 5856 13360 5908
rect 13412 5896 13418 5908
rect 14461 5899 14519 5905
rect 14461 5896 14473 5899
rect 13412 5868 14473 5896
rect 13412 5856 13418 5868
rect 14461 5865 14473 5868
rect 14507 5865 14519 5899
rect 14461 5859 14519 5865
rect 15930 5856 15936 5908
rect 15988 5856 15994 5908
rect 16117 5899 16175 5905
rect 16117 5865 16129 5899
rect 16163 5896 16175 5899
rect 17034 5896 17040 5908
rect 16163 5868 17040 5896
rect 16163 5865 16175 5868
rect 16117 5859 16175 5865
rect 17034 5856 17040 5868
rect 17092 5856 17098 5908
rect 10965 5831 11023 5837
rect 10965 5797 10977 5831
rect 11011 5828 11023 5831
rect 13446 5828 13452 5840
rect 11011 5800 13452 5828
rect 11011 5797 11023 5800
rect 10965 5791 11023 5797
rect 13446 5788 13452 5800
rect 13504 5788 13510 5840
rect 15194 5828 15200 5840
rect 14660 5800 15200 5828
rect 3142 5720 3148 5772
rect 3200 5720 3206 5772
rect 5721 5763 5779 5769
rect 5721 5729 5733 5763
rect 5767 5760 5779 5763
rect 6546 5760 6552 5772
rect 5767 5732 6552 5760
rect 5767 5729 5779 5732
rect 5721 5723 5779 5729
rect 6546 5720 6552 5732
rect 6604 5760 6610 5772
rect 7006 5760 7012 5772
rect 6604 5732 7012 5760
rect 6604 5720 6610 5732
rect 7006 5720 7012 5732
rect 7064 5720 7070 5772
rect 13262 5760 13268 5772
rect 9324 5732 13268 5760
rect 5465 5695 5523 5701
rect 5465 5661 5477 5695
rect 5511 5692 5523 5695
rect 9324 5692 9352 5732
rect 13262 5720 13268 5732
rect 13320 5720 13326 5772
rect 14660 5769 14688 5800
rect 15194 5788 15200 5800
rect 15252 5788 15258 5840
rect 14645 5763 14703 5769
rect 14645 5729 14657 5763
rect 14691 5729 14703 5763
rect 14645 5723 14703 5729
rect 15102 5720 15108 5772
rect 15160 5720 15166 5772
rect 5511 5664 9352 5692
rect 9401 5695 9459 5701
rect 5511 5661 5523 5664
rect 5465 5655 5523 5661
rect 9401 5661 9413 5695
rect 9447 5692 9459 5695
rect 9490 5692 9496 5704
rect 9447 5664 9496 5692
rect 9447 5661 9459 5664
rect 9401 5655 9459 5661
rect 9490 5652 9496 5664
rect 9548 5652 9554 5704
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5692 9735 5695
rect 9723 5664 12434 5692
rect 9723 5661 9735 5664
rect 9677 5655 9735 5661
rect 2900 5627 2958 5633
rect 2900 5593 2912 5627
rect 2946 5624 2958 5627
rect 4430 5624 4436 5636
rect 2946 5596 4436 5624
rect 2946 5593 2958 5596
rect 2900 5587 2958 5593
rect 4430 5584 4436 5596
rect 4488 5584 4494 5636
rect 12406 5624 12434 5664
rect 12986 5652 12992 5704
rect 13044 5652 13050 5704
rect 13173 5695 13231 5701
rect 13173 5661 13185 5695
rect 13219 5692 13231 5695
rect 13814 5692 13820 5704
rect 13219 5664 13820 5692
rect 13219 5661 13231 5664
rect 13173 5655 13231 5661
rect 13814 5652 13820 5664
rect 13872 5652 13878 5704
rect 14737 5695 14795 5701
rect 14737 5661 14749 5695
rect 14783 5661 14795 5695
rect 14737 5655 14795 5661
rect 14752 5624 14780 5655
rect 14826 5652 14832 5704
rect 14884 5652 14890 5704
rect 14921 5695 14979 5701
rect 14921 5661 14933 5695
rect 14967 5692 14979 5695
rect 15120 5692 15148 5720
rect 14967 5664 15148 5692
rect 14967 5661 14979 5664
rect 14921 5655 14979 5661
rect 15102 5624 15108 5636
rect 12406 5596 13860 5624
rect 14752 5596 15108 5624
rect 1762 5516 1768 5568
rect 1820 5516 1826 5568
rect 12802 5516 12808 5568
rect 12860 5516 12866 5568
rect 13832 5556 13860 5596
rect 15102 5584 15108 5596
rect 15160 5584 15166 5636
rect 15746 5584 15752 5636
rect 15804 5584 15810 5636
rect 14274 5556 14280 5568
rect 13832 5528 14280 5556
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 15654 5516 15660 5568
rect 15712 5556 15718 5568
rect 15949 5559 16007 5565
rect 15949 5556 15961 5559
rect 15712 5528 15961 5556
rect 15712 5516 15718 5528
rect 15949 5525 15961 5528
rect 15995 5525 16007 5559
rect 15949 5519 16007 5525
rect 1104 5466 22976 5488
rect 1104 5414 6378 5466
rect 6430 5414 6442 5466
rect 6494 5414 6506 5466
rect 6558 5414 6570 5466
rect 6622 5414 6634 5466
rect 6686 5414 11806 5466
rect 11858 5414 11870 5466
rect 11922 5414 11934 5466
rect 11986 5414 11998 5466
rect 12050 5414 12062 5466
rect 12114 5414 17234 5466
rect 17286 5414 17298 5466
rect 17350 5414 17362 5466
rect 17414 5414 17426 5466
rect 17478 5414 17490 5466
rect 17542 5414 22662 5466
rect 22714 5414 22726 5466
rect 22778 5414 22790 5466
rect 22842 5414 22854 5466
rect 22906 5414 22918 5466
rect 22970 5414 22976 5466
rect 1104 5392 22976 5414
rect 3053 5355 3111 5361
rect 3053 5321 3065 5355
rect 3099 5352 3111 5355
rect 3142 5352 3148 5364
rect 3099 5324 3148 5352
rect 3099 5321 3111 5324
rect 3053 5315 3111 5321
rect 3142 5312 3148 5324
rect 3200 5312 3206 5364
rect 13078 5312 13084 5364
rect 13136 5352 13142 5364
rect 13633 5355 13691 5361
rect 13633 5352 13645 5355
rect 13136 5324 13645 5352
rect 13136 5312 13142 5324
rect 13633 5321 13645 5324
rect 13679 5321 13691 5355
rect 13633 5315 13691 5321
rect 13722 5312 13728 5364
rect 13780 5352 13786 5364
rect 14090 5352 14096 5364
rect 13780 5324 14096 5352
rect 13780 5312 13786 5324
rect 14090 5312 14096 5324
rect 14148 5312 14154 5364
rect 18141 5355 18199 5361
rect 18141 5321 18153 5355
rect 18187 5352 18199 5355
rect 19702 5352 19708 5364
rect 18187 5324 19708 5352
rect 18187 5321 18199 5324
rect 18141 5315 18199 5321
rect 19702 5312 19708 5324
rect 19760 5312 19766 5364
rect 4338 5244 4344 5296
rect 4396 5244 4402 5296
rect 7834 5244 7840 5296
rect 7892 5244 7898 5296
rect 9490 5244 9496 5296
rect 9548 5244 9554 5296
rect 15102 5284 15108 5296
rect 13648 5256 15108 5284
rect 13538 5176 13544 5228
rect 13596 5176 13602 5228
rect 13648 5218 13676 5256
rect 15102 5244 15108 5256
rect 15160 5244 15166 5296
rect 15654 5244 15660 5296
rect 15712 5284 15718 5296
rect 15712 5256 17540 5284
rect 15712 5244 15718 5256
rect 13737 5219 13795 5225
rect 13737 5218 13749 5219
rect 13648 5190 13749 5218
rect 13734 5188 13749 5190
rect 13737 5185 13749 5188
rect 13783 5185 13795 5219
rect 13737 5179 13795 5185
rect 14918 5176 14924 5228
rect 14976 5176 14982 5228
rect 16853 5219 16911 5225
rect 16853 5185 16865 5219
rect 16899 5185 16911 5219
rect 16853 5179 16911 5185
rect 12986 5108 12992 5160
rect 13044 5148 13050 5160
rect 14553 5151 14611 5157
rect 14553 5148 14565 5151
rect 13044 5120 14565 5148
rect 13044 5108 13050 5120
rect 14553 5117 14565 5120
rect 14599 5148 14611 5151
rect 16868 5148 16896 5179
rect 17218 5176 17224 5228
rect 17276 5176 17282 5228
rect 17512 5225 17540 5256
rect 17497 5219 17555 5225
rect 17497 5185 17509 5219
rect 17543 5185 17555 5219
rect 17497 5179 17555 5185
rect 17126 5148 17132 5160
rect 14599 5120 16804 5148
rect 16868 5120 17132 5148
rect 14599 5117 14611 5120
rect 14553 5111 14611 5117
rect 13814 5040 13820 5092
rect 13872 5080 13878 5092
rect 14645 5083 14703 5089
rect 14645 5080 14657 5083
rect 13872 5052 14657 5080
rect 13872 5040 13878 5052
rect 14645 5049 14657 5052
rect 14691 5049 14703 5083
rect 14645 5043 14703 5049
rect 14734 5040 14740 5092
rect 14792 5089 14798 5092
rect 14792 5083 14814 5089
rect 14802 5049 14814 5083
rect 16776 5080 16804 5120
rect 17126 5108 17132 5120
rect 17184 5108 17190 5160
rect 17236 5080 17264 5176
rect 16776 5052 17264 5080
rect 14792 5043 14814 5049
rect 14792 5040 14798 5043
rect 13906 4972 13912 5024
rect 13964 5012 13970 5024
rect 14277 5015 14335 5021
rect 14277 5012 14289 5015
rect 13964 4984 14289 5012
rect 13964 4972 13970 4984
rect 14277 4981 14289 4984
rect 14323 4981 14335 5015
rect 14277 4975 14335 4981
rect 1104 4922 22816 4944
rect 1104 4870 3664 4922
rect 3716 4870 3728 4922
rect 3780 4870 3792 4922
rect 3844 4870 3856 4922
rect 3908 4870 3920 4922
rect 3972 4870 9092 4922
rect 9144 4870 9156 4922
rect 9208 4870 9220 4922
rect 9272 4870 9284 4922
rect 9336 4870 9348 4922
rect 9400 4870 14520 4922
rect 14572 4870 14584 4922
rect 14636 4870 14648 4922
rect 14700 4870 14712 4922
rect 14764 4870 14776 4922
rect 14828 4870 19948 4922
rect 20000 4870 20012 4922
rect 20064 4870 20076 4922
rect 20128 4870 20140 4922
rect 20192 4870 20204 4922
rect 20256 4870 22816 4922
rect 1104 4848 22816 4870
rect 8018 4768 8024 4820
rect 8076 4808 8082 4820
rect 8389 4811 8447 4817
rect 8389 4808 8401 4811
rect 8076 4780 8401 4808
rect 8076 4768 8082 4780
rect 8389 4777 8401 4780
rect 8435 4808 8447 4811
rect 8435 4780 12434 4808
rect 8435 4777 8447 4780
rect 8389 4771 8447 4777
rect 12406 4740 12434 4780
rect 15654 4768 15660 4820
rect 15712 4808 15718 4820
rect 15749 4811 15807 4817
rect 15749 4808 15761 4811
rect 15712 4780 15761 4808
rect 15712 4768 15718 4780
rect 15749 4777 15761 4780
rect 15795 4777 15807 4811
rect 15749 4771 15807 4777
rect 17313 4811 17371 4817
rect 17313 4777 17325 4811
rect 17359 4808 17371 4811
rect 17586 4808 17592 4820
rect 17359 4780 17592 4808
rect 17359 4777 17371 4780
rect 17313 4771 17371 4777
rect 13081 4743 13139 4749
rect 13081 4740 13093 4743
rect 12406 4712 13093 4740
rect 13081 4709 13093 4712
rect 13127 4709 13139 4743
rect 13081 4703 13139 4709
rect 3142 4632 3148 4684
rect 3200 4672 3206 4684
rect 4246 4672 4252 4684
rect 3200 4644 4252 4672
rect 3200 4632 3206 4644
rect 4246 4632 4252 4644
rect 4304 4672 4310 4684
rect 5169 4675 5227 4681
rect 5169 4672 5181 4675
rect 4304 4644 5181 4672
rect 4304 4632 4310 4644
rect 5169 4641 5181 4644
rect 5215 4641 5227 4675
rect 5169 4635 5227 4641
rect 9490 4632 9496 4684
rect 9548 4672 9554 4684
rect 9585 4675 9643 4681
rect 9585 4672 9597 4675
rect 9548 4644 9597 4672
rect 9548 4632 9554 4644
rect 9585 4641 9597 4644
rect 9631 4641 9643 4675
rect 9585 4635 9643 4641
rect 1670 4564 1676 4616
rect 1728 4604 1734 4616
rect 1857 4607 1915 4613
rect 1857 4604 1869 4607
rect 1728 4576 1869 4604
rect 1728 4564 1734 4576
rect 1857 4573 1869 4576
rect 1903 4604 1915 4607
rect 3160 4604 3188 4632
rect 13096 4616 13124 4703
rect 14090 4700 14096 4752
rect 14148 4740 14154 4752
rect 14826 4740 14832 4752
rect 14148 4712 14832 4740
rect 14148 4700 14154 4712
rect 14826 4700 14832 4712
rect 14884 4740 14890 4752
rect 14884 4712 15332 4740
rect 14884 4700 14890 4712
rect 1903 4576 3188 4604
rect 1903 4573 1915 4576
rect 1857 4567 1915 4573
rect 7006 4564 7012 4616
rect 7064 4564 7070 4616
rect 12710 4564 12716 4616
rect 12768 4604 12774 4616
rect 12805 4607 12863 4613
rect 12805 4604 12817 4607
rect 12768 4576 12817 4604
rect 12768 4564 12774 4576
rect 12805 4573 12817 4576
rect 12851 4573 12863 4607
rect 12805 4567 12863 4573
rect 12897 4607 12955 4613
rect 12897 4573 12909 4607
rect 12943 4604 12955 4607
rect 12986 4604 12992 4616
rect 12943 4576 12992 4604
rect 12943 4573 12955 4576
rect 12897 4567 12955 4573
rect 12986 4564 12992 4576
rect 13044 4564 13050 4616
rect 13078 4564 13084 4616
rect 13136 4564 13142 4616
rect 13170 4564 13176 4616
rect 13228 4604 13234 4616
rect 14108 4604 14136 4700
rect 14734 4632 14740 4684
rect 14792 4672 14798 4684
rect 15010 4672 15016 4684
rect 14792 4644 15016 4672
rect 14792 4632 14798 4644
rect 15010 4632 15016 4644
rect 15068 4672 15074 4684
rect 15197 4675 15255 4681
rect 15197 4672 15209 4675
rect 15068 4644 15209 4672
rect 15068 4632 15074 4644
rect 15197 4641 15209 4644
rect 15243 4641 15255 4675
rect 15197 4635 15255 4641
rect 13228 4576 14136 4604
rect 13228 4564 13234 4576
rect 14458 4564 14464 4616
rect 14516 4564 14522 4616
rect 14829 4607 14887 4613
rect 14829 4573 14841 4607
rect 14875 4573 14887 4607
rect 14829 4567 14887 4573
rect 2124 4539 2182 4545
rect 2124 4505 2136 4539
rect 2170 4536 2182 4539
rect 2498 4536 2504 4548
rect 2170 4508 2504 4536
rect 2170 4505 2182 4508
rect 2124 4499 2182 4505
rect 2498 4496 2504 4508
rect 2556 4496 2562 4548
rect 5436 4539 5494 4545
rect 5436 4505 5448 4539
rect 5482 4536 5494 4539
rect 7098 4536 7104 4548
rect 5482 4508 7104 4536
rect 5482 4505 5494 4508
rect 5436 4499 5494 4505
rect 7098 4496 7104 4508
rect 7156 4496 7162 4548
rect 7276 4539 7334 4545
rect 7276 4505 7288 4539
rect 7322 4536 7334 4539
rect 7650 4536 7656 4548
rect 7322 4508 7656 4536
rect 7322 4505 7334 4508
rect 7276 4499 7334 4505
rect 7650 4496 7656 4508
rect 7708 4496 7714 4548
rect 9852 4539 9910 4545
rect 9852 4505 9864 4539
rect 9898 4536 9910 4539
rect 12250 4536 12256 4548
rect 9898 4508 12256 4536
rect 9898 4505 9910 4508
rect 9852 4499 9910 4505
rect 12250 4496 12256 4508
rect 12308 4496 12314 4548
rect 14844 4536 14872 4567
rect 14918 4564 14924 4616
rect 14976 4564 14982 4616
rect 15304 4613 15332 4712
rect 15764 4672 15792 4771
rect 17586 4768 17592 4780
rect 17644 4768 17650 4820
rect 17126 4700 17132 4752
rect 17184 4700 17190 4752
rect 16853 4675 16911 4681
rect 16853 4672 16865 4675
rect 15764 4644 16865 4672
rect 16853 4641 16865 4644
rect 16899 4641 16911 4675
rect 16853 4635 16911 4641
rect 15289 4607 15347 4613
rect 15289 4573 15301 4607
rect 15335 4573 15347 4607
rect 15289 4567 15347 4573
rect 15010 4536 15016 4548
rect 14844 4508 15016 4536
rect 15010 4496 15016 4508
rect 15068 4496 15074 4548
rect 3234 4428 3240 4480
rect 3292 4428 3298 4480
rect 6549 4471 6607 4477
rect 6549 4437 6561 4471
rect 6595 4468 6607 4471
rect 7558 4468 7564 4480
rect 6595 4440 7564 4468
rect 6595 4437 6607 4440
rect 6549 4431 6607 4437
rect 7558 4428 7564 4440
rect 7616 4428 7622 4480
rect 10965 4471 11023 4477
rect 10965 4437 10977 4471
rect 11011 4468 11023 4471
rect 12526 4468 12532 4480
rect 11011 4440 12532 4468
rect 11011 4437 11023 4440
rect 10965 4431 11023 4437
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 12618 4428 12624 4480
rect 12676 4428 12682 4480
rect 1104 4378 22976 4400
rect 1104 4326 6378 4378
rect 6430 4326 6442 4378
rect 6494 4326 6506 4378
rect 6558 4326 6570 4378
rect 6622 4326 6634 4378
rect 6686 4326 11806 4378
rect 11858 4326 11870 4378
rect 11922 4326 11934 4378
rect 11986 4326 11998 4378
rect 12050 4326 12062 4378
rect 12114 4326 17234 4378
rect 17286 4326 17298 4378
rect 17350 4326 17362 4378
rect 17414 4326 17426 4378
rect 17478 4326 17490 4378
rect 17542 4326 22662 4378
rect 22714 4326 22726 4378
rect 22778 4326 22790 4378
rect 22842 4326 22854 4378
rect 22906 4326 22918 4378
rect 22970 4326 22976 4378
rect 1104 4304 22976 4326
rect 12250 4224 12256 4276
rect 12308 4224 12314 4276
rect 12618 4224 12624 4276
rect 12676 4264 12682 4276
rect 12713 4267 12771 4273
rect 12713 4264 12725 4267
rect 12676 4236 12725 4264
rect 12676 4224 12682 4236
rect 12713 4233 12725 4236
rect 12759 4233 12771 4267
rect 12713 4227 12771 4233
rect 14734 4224 14740 4276
rect 14792 4224 14798 4276
rect 7006 4156 7012 4208
rect 7064 4196 7070 4208
rect 9944 4199 10002 4205
rect 7064 4168 9536 4196
rect 7064 4156 7070 4168
rect 1670 4088 1676 4140
rect 1728 4088 1734 4140
rect 1940 4131 1998 4137
rect 1940 4097 1952 4131
rect 1986 4128 1998 4131
rect 2314 4128 2320 4140
rect 1986 4100 2320 4128
rect 1986 4097 1998 4100
rect 1940 4091 1998 4097
rect 2314 4088 2320 4100
rect 2372 4088 2378 4140
rect 4246 4088 4252 4140
rect 4304 4088 4310 4140
rect 4516 4131 4574 4137
rect 4516 4097 4528 4131
rect 4562 4128 4574 4131
rect 4798 4128 4804 4140
rect 4562 4100 4804 4128
rect 4562 4097 4574 4100
rect 4516 4091 4574 4097
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 7116 4137 7144 4168
rect 9508 4140 9536 4168
rect 9944 4165 9956 4199
rect 9990 4196 10002 4199
rect 12158 4196 12164 4208
rect 9990 4168 12164 4196
rect 9990 4165 10002 4168
rect 9944 4159 10002 4165
rect 12158 4156 12164 4168
rect 12216 4156 12222 4208
rect 14752 4196 14780 4224
rect 14752 4168 15056 4196
rect 7101 4131 7159 4137
rect 7101 4097 7113 4131
rect 7147 4097 7159 4131
rect 7101 4091 7159 4097
rect 7368 4131 7426 4137
rect 7368 4097 7380 4131
rect 7414 4128 7426 4131
rect 8938 4128 8944 4140
rect 7414 4100 8944 4128
rect 7414 4097 7426 4100
rect 7368 4091 7426 4097
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 9490 4088 9496 4140
rect 9548 4128 9554 4140
rect 9677 4131 9735 4137
rect 9677 4128 9689 4131
rect 9548 4100 9689 4128
rect 9548 4088 9554 4100
rect 9677 4097 9689 4100
rect 9723 4097 9735 4131
rect 9677 4091 9735 4097
rect 12526 4088 12532 4140
rect 12584 4128 12590 4140
rect 12621 4131 12679 4137
rect 12621 4128 12633 4131
rect 12584 4100 12633 4128
rect 12584 4088 12590 4100
rect 12621 4097 12633 4100
rect 12667 4128 12679 4131
rect 13262 4128 13268 4140
rect 12667 4100 13268 4128
rect 12667 4097 12679 4100
rect 12621 4091 12679 4097
rect 13262 4088 13268 4100
rect 13320 4088 13326 4140
rect 14458 4128 14464 4140
rect 13832 4100 14464 4128
rect 12802 4020 12808 4072
rect 12860 4020 12866 4072
rect 9582 3952 9588 4004
rect 9640 3992 9646 4004
rect 11057 3995 11115 4001
rect 9640 3964 9720 3992
rect 9640 3952 9646 3964
rect 2866 3884 2872 3936
rect 2924 3924 2930 3936
rect 3053 3927 3111 3933
rect 3053 3924 3065 3927
rect 2924 3896 3065 3924
rect 2924 3884 2930 3896
rect 3053 3893 3065 3896
rect 3099 3893 3111 3927
rect 3053 3887 3111 3893
rect 3142 3884 3148 3936
rect 3200 3924 3206 3936
rect 5534 3924 5540 3936
rect 3200 3896 5540 3924
rect 3200 3884 3206 3896
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 5629 3927 5687 3933
rect 5629 3893 5641 3927
rect 5675 3924 5687 3927
rect 5902 3924 5908 3936
rect 5675 3896 5908 3924
rect 5675 3893 5687 3896
rect 5629 3887 5687 3893
rect 5902 3884 5908 3896
rect 5960 3884 5966 3936
rect 8478 3884 8484 3936
rect 8536 3884 8542 3936
rect 9692 3924 9720 3964
rect 11057 3961 11069 3995
rect 11103 3992 11115 3995
rect 13832 3992 13860 4100
rect 14458 4088 14464 4100
rect 14516 4128 14522 4140
rect 14737 4131 14795 4137
rect 14737 4128 14749 4131
rect 14516 4100 14749 4128
rect 14516 4088 14522 4100
rect 14737 4097 14749 4100
rect 14783 4097 14795 4131
rect 14737 4091 14795 4097
rect 14826 4088 14832 4140
rect 14884 4088 14890 4140
rect 15028 4137 15056 4168
rect 15013 4131 15071 4137
rect 15013 4097 15025 4131
rect 15059 4097 15071 4131
rect 15013 4091 15071 4097
rect 15102 4088 15108 4140
rect 15160 4088 15166 4140
rect 15194 4088 15200 4140
rect 15252 4088 15258 4140
rect 11103 3964 13860 3992
rect 15381 3995 15439 4001
rect 11103 3961 11115 3964
rect 11057 3955 11115 3961
rect 15381 3961 15393 3995
rect 15427 3992 15439 3995
rect 17126 3992 17132 4004
rect 15427 3964 17132 3992
rect 15427 3961 15439 3964
rect 15381 3955 15439 3961
rect 17126 3952 17132 3964
rect 17184 3952 17190 4004
rect 15010 3924 15016 3936
rect 9692 3896 15016 3924
rect 15010 3884 15016 3896
rect 15068 3884 15074 3936
rect 1104 3834 22816 3856
rect 1104 3782 3664 3834
rect 3716 3782 3728 3834
rect 3780 3782 3792 3834
rect 3844 3782 3856 3834
rect 3908 3782 3920 3834
rect 3972 3782 9092 3834
rect 9144 3782 9156 3834
rect 9208 3782 9220 3834
rect 9272 3782 9284 3834
rect 9336 3782 9348 3834
rect 9400 3782 14520 3834
rect 14572 3782 14584 3834
rect 14636 3782 14648 3834
rect 14700 3782 14712 3834
rect 14764 3782 14776 3834
rect 14828 3782 19948 3834
rect 20000 3782 20012 3834
rect 20064 3782 20076 3834
rect 20128 3782 20140 3834
rect 20192 3782 20204 3834
rect 20256 3782 22816 3834
rect 1104 3760 22816 3782
rect 4798 3680 4804 3732
rect 4856 3680 4862 3732
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 5592 3692 6914 3720
rect 5592 3680 5598 3692
rect 2866 3652 2872 3664
rect 2332 3624 2872 3652
rect 2332 3593 2360 3624
rect 2866 3612 2872 3624
rect 2924 3612 2930 3664
rect 6886 3652 6914 3692
rect 8202 3680 8208 3732
rect 8260 3720 8266 3732
rect 12802 3720 12808 3732
rect 8260 3692 12808 3720
rect 8260 3680 8266 3692
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 14553 3723 14611 3729
rect 14553 3689 14565 3723
rect 14599 3720 14611 3723
rect 14918 3720 14924 3732
rect 14599 3692 14924 3720
rect 14599 3689 14611 3692
rect 14553 3683 14611 3689
rect 14918 3680 14924 3692
rect 14976 3680 14982 3732
rect 15194 3680 15200 3732
rect 15252 3680 15258 3732
rect 9858 3652 9864 3664
rect 6886 3624 9864 3652
rect 9858 3612 9864 3624
rect 9916 3612 9922 3664
rect 10870 3612 10876 3664
rect 10928 3612 10934 3664
rect 11606 3612 11612 3664
rect 11664 3612 11670 3664
rect 2317 3587 2375 3593
rect 2317 3553 2329 3587
rect 2363 3553 2375 3587
rect 2317 3547 2375 3553
rect 2593 3587 2651 3593
rect 2593 3553 2605 3587
rect 2639 3584 2651 3587
rect 2774 3584 2780 3596
rect 2639 3556 2780 3584
rect 2639 3553 2651 3556
rect 2593 3547 2651 3553
rect 2774 3544 2780 3556
rect 2832 3544 2838 3596
rect 4154 3544 4160 3596
rect 4212 3584 4218 3596
rect 4985 3587 5043 3593
rect 4985 3584 4997 3587
rect 4212 3556 4997 3584
rect 4212 3544 4218 3556
rect 4985 3553 4997 3556
rect 5031 3584 5043 3587
rect 5997 3587 6055 3593
rect 5997 3584 6009 3587
rect 5031 3556 6009 3584
rect 5031 3553 5043 3556
rect 4985 3547 5043 3553
rect 5997 3553 6009 3556
rect 6043 3553 6055 3587
rect 5997 3547 6055 3553
rect 8113 3587 8171 3593
rect 8113 3553 8125 3587
rect 8159 3584 8171 3587
rect 9582 3584 9588 3596
rect 8159 3556 9588 3584
rect 8159 3553 8171 3556
rect 8113 3547 8171 3553
rect 9582 3544 9588 3556
rect 9640 3544 9646 3596
rect 10888 3584 10916 3612
rect 13170 3584 13176 3596
rect 10888 3556 13176 3584
rect 1762 3476 1768 3528
rect 1820 3516 1826 3528
rect 2225 3519 2283 3525
rect 2225 3516 2237 3519
rect 1820 3488 2237 3516
rect 1820 3476 1826 3488
rect 2225 3485 2237 3488
rect 2271 3485 2283 3519
rect 2225 3479 2283 3485
rect 2240 3448 2268 3479
rect 5074 3476 5080 3528
rect 5132 3516 5138 3528
rect 5132 3488 5856 3516
rect 5132 3476 5138 3488
rect 2590 3448 2596 3460
rect 2240 3420 2596 3448
rect 2590 3408 2596 3420
rect 2648 3408 2654 3460
rect 3234 3408 3240 3460
rect 3292 3448 3298 3460
rect 5353 3451 5411 3457
rect 5353 3448 5365 3451
rect 3292 3420 5365 3448
rect 3292 3408 3298 3420
rect 5353 3417 5365 3420
rect 5399 3417 5411 3451
rect 5353 3411 5411 3417
rect 5445 3451 5503 3457
rect 5445 3417 5457 3451
rect 5491 3448 5503 3451
rect 5718 3448 5724 3460
rect 5491 3420 5724 3448
rect 5491 3417 5503 3420
rect 5445 3411 5503 3417
rect 5718 3408 5724 3420
rect 5776 3408 5782 3460
rect 5828 3448 5856 3488
rect 5902 3476 5908 3528
rect 5960 3476 5966 3528
rect 7929 3519 7987 3525
rect 7929 3485 7941 3519
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 7745 3451 7803 3457
rect 7745 3448 7757 3451
rect 5828 3420 7757 3448
rect 7745 3417 7757 3420
rect 7791 3417 7803 3451
rect 7944 3448 7972 3479
rect 9490 3476 9496 3528
rect 9548 3516 9554 3528
rect 10873 3519 10931 3525
rect 10873 3516 10885 3519
rect 9548 3488 10885 3516
rect 9548 3476 9554 3488
rect 10873 3485 10885 3488
rect 10919 3485 10931 3519
rect 10873 3479 10931 3485
rect 11330 3476 11336 3528
rect 11388 3476 11394 3528
rect 11624 3525 11652 3556
rect 13170 3544 13176 3556
rect 13228 3544 13234 3596
rect 11609 3519 11667 3525
rect 11609 3485 11621 3519
rect 11655 3485 11667 3519
rect 11609 3479 11667 3485
rect 12710 3476 12716 3528
rect 12768 3516 12774 3528
rect 13265 3519 13323 3525
rect 13265 3516 13277 3519
rect 12768 3488 13277 3516
rect 12768 3476 12774 3488
rect 13265 3485 13277 3488
rect 13311 3485 13323 3519
rect 13265 3479 13323 3485
rect 14366 3476 14372 3528
rect 14424 3516 14430 3528
rect 14461 3519 14519 3525
rect 14461 3516 14473 3519
rect 14424 3488 14473 3516
rect 14424 3476 14430 3488
rect 14461 3485 14473 3488
rect 14507 3485 14519 3519
rect 14461 3479 14519 3485
rect 14645 3519 14703 3525
rect 14645 3485 14657 3519
rect 14691 3516 14703 3519
rect 15105 3519 15163 3525
rect 15105 3516 15117 3519
rect 14691 3488 15117 3516
rect 14691 3485 14703 3488
rect 14645 3479 14703 3485
rect 15105 3485 15117 3488
rect 15151 3485 15163 3519
rect 15105 3479 15163 3485
rect 8202 3448 8208 3460
rect 7944 3420 8208 3448
rect 7745 3411 7803 3417
rect 8202 3408 8208 3420
rect 8260 3408 8266 3460
rect 10226 3448 10232 3460
rect 9508 3420 10232 3448
rect 9508 3389 9536 3420
rect 10226 3408 10232 3420
rect 10284 3408 10290 3460
rect 10628 3451 10686 3457
rect 10628 3417 10640 3451
rect 10674 3448 10686 3451
rect 10962 3448 10968 3460
rect 10674 3420 10968 3448
rect 10674 3417 10686 3420
rect 10628 3411 10686 3417
rect 10962 3408 10968 3420
rect 11020 3408 11026 3460
rect 12434 3408 12440 3460
rect 12492 3448 12498 3460
rect 13081 3451 13139 3457
rect 13081 3448 13093 3451
rect 12492 3420 13093 3448
rect 12492 3408 12498 3420
rect 13081 3417 13093 3420
rect 13127 3417 13139 3451
rect 13081 3411 13139 3417
rect 13354 3408 13360 3460
rect 13412 3448 13418 3460
rect 14660 3448 14688 3479
rect 13412 3420 14688 3448
rect 13412 3408 13418 3420
rect 9493 3383 9551 3389
rect 9493 3349 9505 3383
rect 9539 3349 9551 3383
rect 9493 3343 9551 3349
rect 10134 3340 10140 3392
rect 10192 3380 10198 3392
rect 10870 3380 10876 3392
rect 10192 3352 10876 3380
rect 10192 3340 10198 3352
rect 10870 3340 10876 3352
rect 10928 3380 10934 3392
rect 11425 3383 11483 3389
rect 11425 3380 11437 3383
rect 10928 3352 11437 3380
rect 10928 3340 10934 3352
rect 11425 3349 11437 3352
rect 11471 3349 11483 3383
rect 11425 3343 11483 3349
rect 13446 3340 13452 3392
rect 13504 3340 13510 3392
rect 1104 3290 22976 3312
rect 1104 3238 6378 3290
rect 6430 3238 6442 3290
rect 6494 3238 6506 3290
rect 6558 3238 6570 3290
rect 6622 3238 6634 3290
rect 6686 3238 11806 3290
rect 11858 3238 11870 3290
rect 11922 3238 11934 3290
rect 11986 3238 11998 3290
rect 12050 3238 12062 3290
rect 12114 3238 17234 3290
rect 17286 3238 17298 3290
rect 17350 3238 17362 3290
rect 17414 3238 17426 3290
rect 17478 3238 17490 3290
rect 17542 3238 22662 3290
rect 22714 3238 22726 3290
rect 22778 3238 22790 3290
rect 22842 3238 22854 3290
rect 22906 3238 22918 3290
rect 22970 3238 22976 3290
rect 1104 3216 22976 3238
rect 2498 3136 2504 3188
rect 2556 3136 2562 3188
rect 7650 3136 7656 3188
rect 7708 3136 7714 3188
rect 8018 3136 8024 3188
rect 8076 3136 8082 3188
rect 8113 3179 8171 3185
rect 8113 3145 8125 3179
rect 8159 3176 8171 3179
rect 10045 3179 10103 3185
rect 10045 3176 10057 3179
rect 8159 3148 10057 3176
rect 8159 3145 8171 3148
rect 8113 3139 8171 3145
rect 10045 3145 10057 3148
rect 10091 3145 10103 3179
rect 13354 3176 13360 3188
rect 10045 3139 10103 3145
rect 10612 3148 13360 3176
rect 5721 3111 5779 3117
rect 5721 3077 5733 3111
rect 5767 3108 5779 3111
rect 10612 3108 10640 3148
rect 13354 3136 13360 3148
rect 13412 3136 13418 3188
rect 13446 3136 13452 3188
rect 13504 3136 13510 3188
rect 15102 3136 15108 3188
rect 15160 3176 15166 3188
rect 15289 3179 15347 3185
rect 15289 3176 15301 3179
rect 15160 3148 15301 3176
rect 15160 3136 15166 3148
rect 15289 3145 15301 3148
rect 15335 3145 15347 3179
rect 15289 3139 15347 3145
rect 5767 3080 10640 3108
rect 10689 3111 10747 3117
rect 5767 3077 5779 3080
rect 5721 3071 5779 3077
rect 10689 3077 10701 3111
rect 10735 3108 10747 3111
rect 11606 3108 11612 3120
rect 10735 3080 11612 3108
rect 10735 3077 10747 3080
rect 10689 3071 10747 3077
rect 11606 3068 11612 3080
rect 11664 3068 11670 3120
rect 13464 3108 13492 3136
rect 13096 3080 13492 3108
rect 2682 3000 2688 3052
rect 2740 3000 2746 3052
rect 2774 3000 2780 3052
rect 2832 3000 2838 3052
rect 3053 3043 3111 3049
rect 3053 3009 3065 3043
rect 3099 3040 3111 3043
rect 3234 3040 3240 3052
rect 3099 3012 3240 3040
rect 3099 3009 3111 3012
rect 3053 3003 3111 3009
rect 3234 3000 3240 3012
rect 3292 3000 3298 3052
rect 4154 3000 4160 3052
rect 4212 3000 4218 3052
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3040 4399 3043
rect 5534 3040 5540 3052
rect 4387 3012 5540 3040
rect 4387 3009 4399 3012
rect 4341 3003 4399 3009
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3040 9091 3043
rect 9490 3040 9496 3052
rect 9079 3012 9496 3040
rect 9079 3009 9091 3012
rect 9033 3003 9091 3009
rect 9490 3000 9496 3012
rect 9548 3040 9554 3052
rect 10321 3043 10379 3049
rect 10321 3040 10333 3043
rect 9548 3012 10333 3040
rect 9548 3000 9554 3012
rect 10321 3009 10333 3012
rect 10367 3009 10379 3043
rect 10321 3003 10379 3009
rect 10870 3000 10876 3052
rect 10928 3040 10934 3052
rect 13096 3049 13124 3080
rect 12069 3043 12127 3049
rect 12069 3040 12081 3043
rect 10928 3012 12081 3040
rect 10928 3000 10934 3012
rect 12069 3009 12081 3012
rect 12115 3009 12127 3043
rect 12069 3003 12127 3009
rect 12161 3043 12219 3049
rect 12161 3009 12173 3043
rect 12207 3040 12219 3043
rect 12897 3043 12955 3049
rect 12897 3040 12909 3043
rect 12207 3012 12909 3040
rect 12207 3009 12219 3012
rect 12161 3003 12219 3009
rect 12897 3009 12909 3012
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3009 13139 3043
rect 13081 3003 13139 3009
rect 13170 3000 13176 3052
rect 13228 3000 13234 3052
rect 13265 3043 13323 3049
rect 13265 3009 13277 3043
rect 13311 3009 13323 3043
rect 13265 3003 13323 3009
rect 3252 2972 3280 3000
rect 4801 2975 4859 2981
rect 4801 2972 4813 2975
rect 3252 2944 4813 2972
rect 4801 2941 4813 2944
rect 4847 2941 4859 2975
rect 4801 2935 4859 2941
rect 5353 2975 5411 2981
rect 5353 2941 5365 2975
rect 5399 2972 5411 2975
rect 5902 2972 5908 2984
rect 5399 2944 5908 2972
rect 5399 2941 5411 2944
rect 5353 2935 5411 2941
rect 5902 2932 5908 2944
rect 5960 2932 5966 2984
rect 8202 2932 8208 2984
rect 8260 2932 8266 2984
rect 8478 2932 8484 2984
rect 8536 2972 8542 2984
rect 9309 2975 9367 2981
rect 9309 2972 9321 2975
rect 8536 2944 9321 2972
rect 8536 2932 8542 2944
rect 9309 2941 9321 2944
rect 9355 2972 9367 2975
rect 10134 2972 10140 2984
rect 9355 2944 10140 2972
rect 9355 2941 9367 2944
rect 9309 2935 9367 2941
rect 10134 2932 10140 2944
rect 10192 2932 10198 2984
rect 10226 2932 10232 2984
rect 10284 2932 10290 2984
rect 10594 2932 10600 2984
rect 10652 2932 10658 2984
rect 12345 2975 12403 2981
rect 12345 2941 12357 2975
rect 12391 2941 12403 2975
rect 12345 2935 12403 2941
rect 2866 2864 2872 2916
rect 2924 2904 2930 2916
rect 5169 2907 5227 2913
rect 5169 2904 5181 2907
rect 2924 2876 5181 2904
rect 2924 2864 2930 2876
rect 5169 2873 5181 2876
rect 5215 2873 5227 2907
rect 5169 2867 5227 2873
rect 8938 2864 8944 2916
rect 8996 2904 9002 2916
rect 11701 2907 11759 2913
rect 11701 2904 11713 2907
rect 8996 2876 11713 2904
rect 8996 2864 9002 2876
rect 11701 2873 11713 2876
rect 11747 2873 11759 2907
rect 12360 2904 12388 2935
rect 12802 2904 12808 2916
rect 12360 2876 12808 2904
rect 11701 2867 11759 2873
rect 12802 2864 12808 2876
rect 12860 2864 12866 2916
rect 13280 2904 13308 3003
rect 13354 3000 13360 3052
rect 13412 3049 13418 3052
rect 13412 3043 13441 3049
rect 13429 3009 13441 3043
rect 13412 3003 13441 3009
rect 13541 3043 13599 3049
rect 13541 3009 13553 3043
rect 13587 3040 13599 3043
rect 14366 3040 14372 3052
rect 13587 3012 14372 3040
rect 13587 3009 13599 3012
rect 13541 3003 13599 3009
rect 13412 3000 13418 3003
rect 14366 3000 14372 3012
rect 14424 3040 14430 3052
rect 14461 3043 14519 3049
rect 14461 3040 14473 3043
rect 14424 3012 14473 3040
rect 14424 3000 14430 3012
rect 14461 3009 14473 3012
rect 14507 3009 14519 3043
rect 14461 3003 14519 3009
rect 14645 3043 14703 3049
rect 14645 3009 14657 3043
rect 14691 3040 14703 3043
rect 15197 3043 15255 3049
rect 15197 3040 15209 3043
rect 14691 3012 15209 3040
rect 14691 3009 14703 3012
rect 14645 3003 14703 3009
rect 15197 3009 15209 3012
rect 15243 3009 15255 3043
rect 15197 3003 15255 3009
rect 14274 2932 14280 2984
rect 14332 2972 14338 2984
rect 14660 2972 14688 3003
rect 14332 2944 14688 2972
rect 14332 2932 14338 2944
rect 14645 2907 14703 2913
rect 14645 2904 14657 2907
rect 13280 2876 14657 2904
rect 14645 2873 14657 2876
rect 14691 2904 14703 2907
rect 15010 2904 15016 2916
rect 14691 2876 15016 2904
rect 14691 2873 14703 2876
rect 14645 2867 14703 2873
rect 15010 2864 15016 2876
rect 15068 2864 15074 2916
rect 2958 2796 2964 2848
rect 3016 2796 3022 2848
rect 4338 2796 4344 2848
rect 4396 2796 4402 2848
rect 5258 2796 5264 2848
rect 5316 2796 5322 2848
rect 8846 2796 8852 2848
rect 8904 2796 8910 2848
rect 9217 2839 9275 2845
rect 9217 2805 9229 2839
rect 9263 2836 9275 2839
rect 9582 2836 9588 2848
rect 9263 2808 9588 2836
rect 9263 2805 9275 2808
rect 9217 2799 9275 2805
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 10226 2796 10232 2848
rect 10284 2836 10290 2848
rect 12618 2836 12624 2848
rect 10284 2808 12624 2836
rect 10284 2796 10290 2808
rect 12618 2796 12624 2808
rect 12676 2796 12682 2848
rect 1104 2746 22816 2768
rect 1104 2694 3664 2746
rect 3716 2694 3728 2746
rect 3780 2694 3792 2746
rect 3844 2694 3856 2746
rect 3908 2694 3920 2746
rect 3972 2694 9092 2746
rect 9144 2694 9156 2746
rect 9208 2694 9220 2746
rect 9272 2694 9284 2746
rect 9336 2694 9348 2746
rect 9400 2694 14520 2746
rect 14572 2694 14584 2746
rect 14636 2694 14648 2746
rect 14700 2694 14712 2746
rect 14764 2694 14776 2746
rect 14828 2694 19948 2746
rect 20000 2694 20012 2746
rect 20064 2694 20076 2746
rect 20128 2694 20140 2746
rect 20192 2694 20204 2746
rect 20256 2694 22816 2746
rect 1104 2672 22816 2694
rect 2314 2592 2320 2644
rect 2372 2592 2378 2644
rect 4341 2635 4399 2641
rect 4341 2601 4353 2635
rect 4387 2632 4399 2635
rect 4430 2632 4436 2644
rect 4387 2604 4436 2632
rect 4387 2601 4399 2604
rect 4341 2595 4399 2601
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 5718 2592 5724 2644
rect 5776 2592 5782 2644
rect 7098 2592 7104 2644
rect 7156 2632 7162 2644
rect 7193 2635 7251 2641
rect 7193 2632 7205 2635
rect 7156 2604 7205 2632
rect 7156 2592 7162 2604
rect 7193 2601 7205 2604
rect 7239 2601 7251 2635
rect 7193 2595 7251 2601
rect 9217 2635 9275 2641
rect 9217 2601 9229 2635
rect 9263 2632 9275 2635
rect 9490 2632 9496 2644
rect 9263 2604 9496 2632
rect 9263 2601 9275 2604
rect 9217 2595 9275 2601
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 12529 2635 12587 2641
rect 12529 2601 12541 2635
rect 12575 2632 12587 2635
rect 13170 2632 13176 2644
rect 12575 2604 13176 2632
rect 12575 2601 12587 2604
rect 12529 2595 12587 2601
rect 13170 2592 13176 2604
rect 13228 2592 13234 2644
rect 13354 2592 13360 2644
rect 13412 2632 13418 2644
rect 13449 2635 13507 2641
rect 13449 2632 13461 2635
rect 13412 2604 13461 2632
rect 13412 2592 13418 2604
rect 13449 2601 13461 2604
rect 13495 2601 13507 2635
rect 13449 2595 13507 2601
rect 2777 2567 2835 2573
rect 2777 2533 2789 2567
rect 2823 2564 2835 2567
rect 2958 2564 2964 2576
rect 2823 2536 2964 2564
rect 2823 2533 2835 2536
rect 2777 2527 2835 2533
rect 2958 2524 2964 2536
rect 3016 2564 3022 2576
rect 12434 2564 12440 2576
rect 3016 2536 5028 2564
rect 3016 2524 3022 2536
rect 2608 2468 4200 2496
rect 2608 2440 2636 2468
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 2516 2360 2544 2391
rect 2590 2388 2596 2440
rect 2648 2388 2654 2440
rect 2866 2388 2872 2440
rect 2924 2388 2930 2440
rect 4172 2428 4200 2468
rect 4338 2456 4344 2508
rect 4396 2496 4402 2508
rect 5000 2505 5028 2536
rect 9140 2536 12440 2564
rect 4801 2499 4859 2505
rect 4801 2496 4813 2499
rect 4396 2468 4813 2496
rect 4396 2456 4402 2468
rect 4801 2465 4813 2468
rect 4847 2465 4859 2499
rect 4801 2459 4859 2465
rect 4985 2499 5043 2505
rect 4985 2465 4997 2499
rect 5031 2496 5043 2499
rect 5074 2496 5080 2508
rect 5031 2468 5080 2496
rect 5031 2465 5043 2468
rect 4985 2459 5043 2465
rect 5074 2456 5080 2468
rect 5132 2456 5138 2508
rect 7837 2499 7895 2505
rect 7837 2465 7849 2499
rect 7883 2496 7895 2499
rect 8202 2496 8208 2508
rect 7883 2468 8208 2496
rect 7883 2465 7895 2468
rect 7837 2459 7895 2465
rect 8202 2456 8208 2468
rect 8260 2456 8266 2508
rect 8754 2456 8760 2508
rect 8812 2496 8818 2508
rect 9140 2496 9168 2536
rect 12434 2524 12440 2536
rect 12492 2524 12498 2576
rect 8812 2468 9168 2496
rect 8812 2456 8818 2468
rect 4709 2431 4767 2437
rect 4709 2428 4721 2431
rect 4172 2400 4721 2428
rect 4709 2397 4721 2400
rect 4755 2428 4767 2431
rect 5258 2428 5264 2440
rect 4755 2400 5264 2428
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2428 5871 2431
rect 5859 2400 6914 2428
rect 5859 2397 5871 2400
rect 5813 2391 5871 2397
rect 2682 2360 2688 2372
rect 2516 2332 2688 2360
rect 2682 2320 2688 2332
rect 2740 2360 2746 2372
rect 5828 2360 5856 2391
rect 2740 2332 5856 2360
rect 2740 2320 2746 2332
rect 6886 2292 6914 2400
rect 7558 2388 7564 2440
rect 7616 2388 7622 2440
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2428 7711 2431
rect 8846 2428 8852 2440
rect 7699 2400 8852 2428
rect 7699 2397 7711 2400
rect 7653 2391 7711 2397
rect 8846 2388 8852 2400
rect 8904 2388 8910 2440
rect 9140 2437 9168 2468
rect 10594 2456 10600 2508
rect 10652 2496 10658 2508
rect 10781 2499 10839 2505
rect 10781 2496 10793 2499
rect 10652 2468 10793 2496
rect 10652 2456 10658 2468
rect 10781 2465 10793 2468
rect 10827 2496 10839 2499
rect 13449 2499 13507 2505
rect 13449 2496 13461 2499
rect 10827 2468 13461 2496
rect 10827 2465 10839 2468
rect 10781 2459 10839 2465
rect 13449 2465 13461 2468
rect 13495 2465 13507 2499
rect 13449 2459 13507 2465
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 9582 2428 9588 2440
rect 9355 2400 9588 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 9582 2388 9588 2400
rect 9640 2388 9646 2440
rect 10134 2388 10140 2440
rect 10192 2428 10198 2440
rect 10965 2431 11023 2437
rect 10965 2428 10977 2431
rect 10192 2400 10977 2428
rect 10192 2388 10198 2400
rect 10965 2397 10977 2400
rect 11011 2397 11023 2431
rect 10965 2391 11023 2397
rect 12434 2388 12440 2440
rect 12492 2388 12498 2440
rect 12618 2388 12624 2440
rect 12676 2388 12682 2440
rect 13078 2388 13084 2440
rect 13136 2388 13142 2440
rect 7576 2360 7604 2388
rect 11149 2363 11207 2369
rect 11149 2360 11161 2363
rect 7576 2332 11161 2360
rect 11149 2329 11161 2332
rect 11195 2360 11207 2363
rect 11330 2360 11336 2372
rect 11195 2332 11336 2360
rect 11195 2329 11207 2332
rect 11149 2323 11207 2329
rect 11330 2320 11336 2332
rect 11388 2320 11394 2372
rect 13906 2360 13912 2372
rect 11440 2332 13912 2360
rect 11440 2292 11468 2332
rect 13906 2320 13912 2332
rect 13964 2320 13970 2372
rect 6886 2264 11468 2292
rect 13265 2295 13323 2301
rect 13265 2261 13277 2295
rect 13311 2292 13323 2295
rect 14274 2292 14280 2304
rect 13311 2264 14280 2292
rect 13311 2261 13323 2264
rect 13265 2255 13323 2261
rect 14274 2252 14280 2264
rect 14332 2252 14338 2304
rect 1104 2202 22976 2224
rect 1104 2150 6378 2202
rect 6430 2150 6442 2202
rect 6494 2150 6506 2202
rect 6558 2150 6570 2202
rect 6622 2150 6634 2202
rect 6686 2150 11806 2202
rect 11858 2150 11870 2202
rect 11922 2150 11934 2202
rect 11986 2150 11998 2202
rect 12050 2150 12062 2202
rect 12114 2150 17234 2202
rect 17286 2150 17298 2202
rect 17350 2150 17362 2202
rect 17414 2150 17426 2202
rect 17478 2150 17490 2202
rect 17542 2150 22662 2202
rect 22714 2150 22726 2202
rect 22778 2150 22790 2202
rect 22842 2150 22854 2202
rect 22906 2150 22918 2202
rect 22970 2150 22976 2202
rect 1104 2128 22976 2150
<< via1 >>
rect 6378 21734 6430 21786
rect 6442 21734 6494 21786
rect 6506 21734 6558 21786
rect 6570 21734 6622 21786
rect 6634 21734 6686 21786
rect 11806 21734 11858 21786
rect 11870 21734 11922 21786
rect 11934 21734 11986 21786
rect 11998 21734 12050 21786
rect 12062 21734 12114 21786
rect 17234 21734 17286 21786
rect 17298 21734 17350 21786
rect 17362 21734 17414 21786
rect 17426 21734 17478 21786
rect 17490 21734 17542 21786
rect 22662 21734 22714 21786
rect 22726 21734 22778 21786
rect 22790 21734 22842 21786
rect 22854 21734 22906 21786
rect 22918 21734 22970 21786
rect 3664 21190 3716 21242
rect 3728 21190 3780 21242
rect 3792 21190 3844 21242
rect 3856 21190 3908 21242
rect 3920 21190 3972 21242
rect 9092 21190 9144 21242
rect 9156 21190 9208 21242
rect 9220 21190 9272 21242
rect 9284 21190 9336 21242
rect 9348 21190 9400 21242
rect 14520 21190 14572 21242
rect 14584 21190 14636 21242
rect 14648 21190 14700 21242
rect 14712 21190 14764 21242
rect 14776 21190 14828 21242
rect 19948 21190 20000 21242
rect 20012 21190 20064 21242
rect 20076 21190 20128 21242
rect 20140 21190 20192 21242
rect 20204 21190 20256 21242
rect 6378 20646 6430 20698
rect 6442 20646 6494 20698
rect 6506 20646 6558 20698
rect 6570 20646 6622 20698
rect 6634 20646 6686 20698
rect 11806 20646 11858 20698
rect 11870 20646 11922 20698
rect 11934 20646 11986 20698
rect 11998 20646 12050 20698
rect 12062 20646 12114 20698
rect 17234 20646 17286 20698
rect 17298 20646 17350 20698
rect 17362 20646 17414 20698
rect 17426 20646 17478 20698
rect 17490 20646 17542 20698
rect 22662 20646 22714 20698
rect 22726 20646 22778 20698
rect 22790 20646 22842 20698
rect 22854 20646 22906 20698
rect 22918 20646 22970 20698
rect 3664 20102 3716 20154
rect 3728 20102 3780 20154
rect 3792 20102 3844 20154
rect 3856 20102 3908 20154
rect 3920 20102 3972 20154
rect 9092 20102 9144 20154
rect 9156 20102 9208 20154
rect 9220 20102 9272 20154
rect 9284 20102 9336 20154
rect 9348 20102 9400 20154
rect 14520 20102 14572 20154
rect 14584 20102 14636 20154
rect 14648 20102 14700 20154
rect 14712 20102 14764 20154
rect 14776 20102 14828 20154
rect 19948 20102 20000 20154
rect 20012 20102 20064 20154
rect 20076 20102 20128 20154
rect 20140 20102 20192 20154
rect 20204 20102 20256 20154
rect 940 19796 992 19848
rect 1584 19728 1636 19780
rect 6378 19558 6430 19610
rect 6442 19558 6494 19610
rect 6506 19558 6558 19610
rect 6570 19558 6622 19610
rect 6634 19558 6686 19610
rect 11806 19558 11858 19610
rect 11870 19558 11922 19610
rect 11934 19558 11986 19610
rect 11998 19558 12050 19610
rect 12062 19558 12114 19610
rect 17234 19558 17286 19610
rect 17298 19558 17350 19610
rect 17362 19558 17414 19610
rect 17426 19558 17478 19610
rect 17490 19558 17542 19610
rect 22662 19558 22714 19610
rect 22726 19558 22778 19610
rect 22790 19558 22842 19610
rect 22854 19558 22906 19610
rect 22918 19558 22970 19610
rect 3664 19014 3716 19066
rect 3728 19014 3780 19066
rect 3792 19014 3844 19066
rect 3856 19014 3908 19066
rect 3920 19014 3972 19066
rect 9092 19014 9144 19066
rect 9156 19014 9208 19066
rect 9220 19014 9272 19066
rect 9284 19014 9336 19066
rect 9348 19014 9400 19066
rect 14520 19014 14572 19066
rect 14584 19014 14636 19066
rect 14648 19014 14700 19066
rect 14712 19014 14764 19066
rect 14776 19014 14828 19066
rect 19948 19014 20000 19066
rect 20012 19014 20064 19066
rect 20076 19014 20128 19066
rect 20140 19014 20192 19066
rect 20204 19014 20256 19066
rect 6378 18470 6430 18522
rect 6442 18470 6494 18522
rect 6506 18470 6558 18522
rect 6570 18470 6622 18522
rect 6634 18470 6686 18522
rect 11806 18470 11858 18522
rect 11870 18470 11922 18522
rect 11934 18470 11986 18522
rect 11998 18470 12050 18522
rect 12062 18470 12114 18522
rect 17234 18470 17286 18522
rect 17298 18470 17350 18522
rect 17362 18470 17414 18522
rect 17426 18470 17478 18522
rect 17490 18470 17542 18522
rect 22662 18470 22714 18522
rect 22726 18470 22778 18522
rect 22790 18470 22842 18522
rect 22854 18470 22906 18522
rect 22918 18470 22970 18522
rect 8852 18275 8904 18284
rect 8852 18241 8861 18275
rect 8861 18241 8895 18275
rect 8895 18241 8904 18275
rect 8852 18232 8904 18241
rect 8392 18164 8444 18216
rect 8944 18071 8996 18080
rect 8944 18037 8953 18071
rect 8953 18037 8987 18071
rect 8987 18037 8996 18071
rect 8944 18028 8996 18037
rect 3664 17926 3716 17978
rect 3728 17926 3780 17978
rect 3792 17926 3844 17978
rect 3856 17926 3908 17978
rect 3920 17926 3972 17978
rect 9092 17926 9144 17978
rect 9156 17926 9208 17978
rect 9220 17926 9272 17978
rect 9284 17926 9336 17978
rect 9348 17926 9400 17978
rect 14520 17926 14572 17978
rect 14584 17926 14636 17978
rect 14648 17926 14700 17978
rect 14712 17926 14764 17978
rect 14776 17926 14828 17978
rect 19948 17926 20000 17978
rect 20012 17926 20064 17978
rect 20076 17926 20128 17978
rect 20140 17926 20192 17978
rect 20204 17926 20256 17978
rect 5724 17688 5776 17740
rect 7012 17663 7064 17672
rect 7012 17629 7021 17663
rect 7021 17629 7055 17663
rect 7055 17629 7064 17663
rect 7012 17620 7064 17629
rect 8944 17756 8996 17808
rect 9312 17756 9364 17808
rect 9404 17688 9456 17740
rect 10876 17688 10928 17740
rect 7196 17663 7248 17672
rect 7196 17629 7205 17663
rect 7205 17629 7239 17663
rect 7239 17629 7248 17663
rect 7196 17620 7248 17629
rect 8208 17663 8260 17672
rect 8208 17629 8217 17663
rect 8217 17629 8251 17663
rect 8251 17629 8260 17663
rect 8208 17620 8260 17629
rect 8300 17663 8352 17672
rect 8300 17629 8309 17663
rect 8309 17629 8343 17663
rect 8343 17629 8352 17663
rect 8300 17620 8352 17629
rect 8852 17620 8904 17672
rect 9312 17663 9364 17672
rect 9312 17629 9321 17663
rect 9321 17629 9355 17663
rect 9355 17629 9364 17663
rect 9312 17620 9364 17629
rect 9956 17620 10008 17672
rect 10600 17620 10652 17672
rect 4712 17527 4764 17536
rect 4712 17493 4721 17527
rect 4721 17493 4755 17527
rect 4755 17493 4764 17527
rect 4712 17484 4764 17493
rect 4896 17484 4948 17536
rect 7104 17484 7156 17536
rect 9496 17484 9548 17536
rect 10600 17484 10652 17536
rect 6378 17382 6430 17434
rect 6442 17382 6494 17434
rect 6506 17382 6558 17434
rect 6570 17382 6622 17434
rect 6634 17382 6686 17434
rect 11806 17382 11858 17434
rect 11870 17382 11922 17434
rect 11934 17382 11986 17434
rect 11998 17382 12050 17434
rect 12062 17382 12114 17434
rect 17234 17382 17286 17434
rect 17298 17382 17350 17434
rect 17362 17382 17414 17434
rect 17426 17382 17478 17434
rect 17490 17382 17542 17434
rect 22662 17382 22714 17434
rect 22726 17382 22778 17434
rect 22790 17382 22842 17434
rect 22854 17382 22906 17434
rect 22918 17382 22970 17434
rect 8116 17280 8168 17332
rect 8852 17280 8904 17332
rect 9404 17323 9456 17332
rect 9404 17289 9413 17323
rect 9413 17289 9447 17323
rect 9447 17289 9456 17323
rect 9404 17280 9456 17289
rect 7012 17212 7064 17264
rect 3332 17144 3384 17196
rect 5080 17144 5132 17196
rect 3240 17119 3292 17128
rect 3240 17085 3249 17119
rect 3249 17085 3283 17119
rect 3283 17085 3292 17119
rect 3240 17076 3292 17085
rect 5724 17076 5776 17128
rect 7196 17187 7248 17196
rect 7196 17153 7205 17187
rect 7205 17153 7239 17187
rect 7239 17153 7248 17187
rect 7196 17144 7248 17153
rect 8116 17187 8168 17196
rect 8116 17153 8125 17187
rect 8125 17153 8159 17187
rect 8159 17153 8168 17187
rect 8116 17144 8168 17153
rect 8392 17144 8444 17196
rect 8944 17144 8996 17196
rect 9680 17187 9732 17196
rect 9680 17153 9689 17187
rect 9689 17153 9723 17187
rect 9723 17153 9732 17187
rect 9680 17144 9732 17153
rect 9956 17187 10008 17196
rect 9956 17153 9965 17187
rect 9965 17153 9999 17187
rect 9999 17153 10008 17187
rect 9956 17144 10008 17153
rect 10692 17144 10744 17196
rect 10876 17076 10928 17128
rect 2688 16983 2740 16992
rect 2688 16949 2697 16983
rect 2697 16949 2731 16983
rect 2731 16949 2740 16983
rect 2688 16940 2740 16949
rect 4804 16983 4856 16992
rect 4804 16949 4813 16983
rect 4813 16949 4847 16983
rect 4847 16949 4856 16983
rect 4804 16940 4856 16949
rect 8300 17008 8352 17060
rect 10508 16940 10560 16992
rect 3664 16838 3716 16890
rect 3728 16838 3780 16890
rect 3792 16838 3844 16890
rect 3856 16838 3908 16890
rect 3920 16838 3972 16890
rect 9092 16838 9144 16890
rect 9156 16838 9208 16890
rect 9220 16838 9272 16890
rect 9284 16838 9336 16890
rect 9348 16838 9400 16890
rect 14520 16838 14572 16890
rect 14584 16838 14636 16890
rect 14648 16838 14700 16890
rect 14712 16838 14764 16890
rect 14776 16838 14828 16890
rect 19948 16838 20000 16890
rect 20012 16838 20064 16890
rect 20076 16838 20128 16890
rect 20140 16838 20192 16890
rect 20204 16838 20256 16890
rect 4896 16600 4948 16652
rect 5724 16643 5776 16652
rect 5724 16609 5733 16643
rect 5733 16609 5767 16643
rect 5767 16609 5776 16643
rect 5724 16600 5776 16609
rect 6736 16600 6788 16652
rect 5080 16532 5132 16584
rect 5632 16575 5684 16584
rect 5632 16541 5641 16575
rect 5641 16541 5675 16575
rect 5675 16541 5684 16575
rect 5632 16532 5684 16541
rect 7472 16736 7524 16788
rect 8300 16736 8352 16788
rect 10508 16736 10560 16788
rect 7196 16668 7248 16720
rect 9956 16668 10008 16720
rect 9680 16600 9732 16652
rect 7288 16575 7340 16584
rect 7288 16541 7323 16575
rect 7323 16541 7340 16575
rect 7288 16532 7340 16541
rect 7472 16575 7524 16584
rect 7472 16541 7481 16575
rect 7481 16541 7515 16575
rect 7515 16541 7524 16575
rect 7472 16532 7524 16541
rect 8116 16575 8168 16584
rect 8116 16541 8125 16575
rect 8125 16541 8159 16575
rect 8159 16541 8168 16575
rect 8116 16532 8168 16541
rect 9496 16532 9548 16584
rect 10600 16575 10652 16584
rect 10600 16541 10609 16575
rect 10609 16541 10643 16575
rect 10643 16541 10652 16575
rect 10600 16532 10652 16541
rect 10968 16532 11020 16584
rect 5172 16464 5224 16516
rect 2596 16439 2648 16448
rect 2596 16405 2605 16439
rect 2605 16405 2639 16439
rect 2639 16405 2648 16439
rect 2596 16396 2648 16405
rect 3332 16396 3384 16448
rect 7196 16507 7248 16516
rect 7196 16473 7205 16507
rect 7205 16473 7239 16507
rect 7239 16473 7248 16507
rect 7196 16464 7248 16473
rect 8392 16464 8444 16516
rect 10416 16464 10468 16516
rect 6378 16294 6430 16346
rect 6442 16294 6494 16346
rect 6506 16294 6558 16346
rect 6570 16294 6622 16346
rect 6634 16294 6686 16346
rect 11806 16294 11858 16346
rect 11870 16294 11922 16346
rect 11934 16294 11986 16346
rect 11998 16294 12050 16346
rect 12062 16294 12114 16346
rect 17234 16294 17286 16346
rect 17298 16294 17350 16346
rect 17362 16294 17414 16346
rect 17426 16294 17478 16346
rect 17490 16294 17542 16346
rect 22662 16294 22714 16346
rect 22726 16294 22778 16346
rect 22790 16294 22842 16346
rect 22854 16294 22906 16346
rect 22918 16294 22970 16346
rect 2688 16192 2740 16244
rect 4804 16192 4856 16244
rect 6920 16192 6972 16244
rect 7196 16192 7248 16244
rect 7472 16192 7524 16244
rect 14372 16192 14424 16244
rect 10140 16124 10192 16176
rect 10692 16124 10744 16176
rect 3056 16056 3108 16108
rect 5264 16056 5316 16108
rect 9496 16056 9548 16108
rect 9680 16056 9732 16108
rect 2688 16031 2740 16040
rect 2688 15997 2697 16031
rect 2697 15997 2731 16031
rect 2731 15997 2740 16031
rect 2688 15988 2740 15997
rect 5172 15988 5224 16040
rect 8116 15988 8168 16040
rect 8392 16031 8444 16040
rect 8392 15997 8401 16031
rect 8401 15997 8435 16031
rect 8435 15997 8444 16031
rect 8392 15988 8444 15997
rect 11060 16056 11112 16108
rect 10324 15988 10376 16040
rect 2044 15852 2096 15904
rect 4528 15852 4580 15904
rect 7196 15852 7248 15904
rect 3664 15750 3716 15802
rect 3728 15750 3780 15802
rect 3792 15750 3844 15802
rect 3856 15750 3908 15802
rect 3920 15750 3972 15802
rect 9092 15750 9144 15802
rect 9156 15750 9208 15802
rect 9220 15750 9272 15802
rect 9284 15750 9336 15802
rect 9348 15750 9400 15802
rect 14520 15750 14572 15802
rect 14584 15750 14636 15802
rect 14648 15750 14700 15802
rect 14712 15750 14764 15802
rect 14776 15750 14828 15802
rect 19948 15750 20000 15802
rect 20012 15750 20064 15802
rect 20076 15750 20128 15802
rect 20140 15750 20192 15802
rect 20204 15750 20256 15802
rect 10416 15691 10468 15700
rect 10416 15657 10425 15691
rect 10425 15657 10459 15691
rect 10459 15657 10468 15691
rect 10416 15648 10468 15657
rect 10968 15623 11020 15632
rect 10968 15589 10977 15623
rect 10977 15589 11011 15623
rect 11011 15589 11020 15623
rect 10968 15580 11020 15589
rect 4712 15512 4764 15564
rect 5172 15512 5224 15564
rect 6920 15444 6972 15496
rect 7196 15487 7248 15496
rect 7196 15453 7205 15487
rect 7205 15453 7239 15487
rect 7239 15453 7248 15487
rect 7196 15444 7248 15453
rect 10324 15487 10376 15496
rect 10324 15453 10333 15487
rect 10333 15453 10367 15487
rect 10367 15453 10376 15487
rect 10324 15444 10376 15453
rect 11060 15444 11112 15496
rect 10876 15376 10928 15428
rect 4436 15308 4488 15360
rect 5080 15308 5132 15360
rect 5540 15308 5592 15360
rect 9220 15351 9272 15360
rect 9220 15317 9229 15351
rect 9229 15317 9263 15351
rect 9263 15317 9272 15351
rect 9220 15308 9272 15317
rect 6378 15206 6430 15258
rect 6442 15206 6494 15258
rect 6506 15206 6558 15258
rect 6570 15206 6622 15258
rect 6634 15206 6686 15258
rect 11806 15206 11858 15258
rect 11870 15206 11922 15258
rect 11934 15206 11986 15258
rect 11998 15206 12050 15258
rect 12062 15206 12114 15258
rect 17234 15206 17286 15258
rect 17298 15206 17350 15258
rect 17362 15206 17414 15258
rect 17426 15206 17478 15258
rect 17490 15206 17542 15258
rect 22662 15206 22714 15258
rect 22726 15206 22778 15258
rect 22790 15206 22842 15258
rect 22854 15206 22906 15258
rect 22918 15206 22970 15258
rect 8116 15104 8168 15156
rect 8208 15104 8260 15156
rect 2412 15036 2464 15088
rect 1860 15011 1912 15020
rect 1860 14977 1869 15011
rect 1869 14977 1903 15011
rect 1903 14977 1912 15011
rect 1860 14968 1912 14977
rect 2136 15011 2188 15020
rect 2136 14977 2145 15011
rect 2145 14977 2179 15011
rect 2179 14977 2188 15011
rect 3240 15036 3292 15088
rect 5540 15036 5592 15088
rect 2136 14968 2188 14977
rect 3056 14968 3108 15020
rect 3332 14968 3384 15020
rect 4068 14968 4120 15020
rect 4804 15011 4856 15020
rect 4804 14977 4813 15011
rect 4813 14977 4847 15011
rect 4847 14977 4856 15011
rect 4804 14968 4856 14977
rect 4896 15011 4948 15020
rect 4896 14977 4905 15011
rect 4905 14977 4939 15011
rect 4939 14977 4948 15011
rect 4896 14968 4948 14977
rect 5264 14968 5316 15020
rect 8300 14968 8352 15020
rect 8944 15011 8996 15020
rect 8944 14977 8953 15011
rect 8953 14977 8987 15011
rect 8987 14977 8996 15011
rect 8944 14968 8996 14977
rect 9220 14968 9272 15020
rect 10140 15011 10192 15020
rect 10140 14977 10149 15011
rect 10149 14977 10183 15011
rect 10183 14977 10192 15011
rect 10140 14968 10192 14977
rect 7012 14900 7064 14952
rect 8852 14943 8904 14952
rect 8852 14909 8861 14943
rect 8861 14909 8895 14943
rect 8895 14909 8904 14943
rect 8852 14900 8904 14909
rect 8116 14832 8168 14884
rect 9496 14900 9548 14952
rect 10876 15011 10928 15020
rect 10876 14977 10885 15011
rect 10885 14977 10919 15011
rect 10919 14977 10928 15011
rect 10876 14968 10928 14977
rect 11060 15011 11112 15020
rect 11060 14977 11069 15011
rect 11069 14977 11103 15011
rect 11103 14977 11112 15011
rect 11060 14968 11112 14977
rect 10968 14900 11020 14952
rect 1768 14764 1820 14816
rect 3424 14764 3476 14816
rect 5540 14764 5592 14816
rect 6644 14764 6696 14816
rect 3664 14662 3716 14714
rect 3728 14662 3780 14714
rect 3792 14662 3844 14714
rect 3856 14662 3908 14714
rect 3920 14662 3972 14714
rect 9092 14662 9144 14714
rect 9156 14662 9208 14714
rect 9220 14662 9272 14714
rect 9284 14662 9336 14714
rect 9348 14662 9400 14714
rect 14520 14662 14572 14714
rect 14584 14662 14636 14714
rect 14648 14662 14700 14714
rect 14712 14662 14764 14714
rect 14776 14662 14828 14714
rect 19948 14662 20000 14714
rect 20012 14662 20064 14714
rect 20076 14662 20128 14714
rect 20140 14662 20192 14714
rect 20204 14662 20256 14714
rect 1584 14560 1636 14612
rect 4068 14560 4120 14612
rect 3516 14492 3568 14544
rect 5172 14560 5224 14612
rect 4344 14467 4396 14476
rect 4344 14433 4353 14467
rect 4353 14433 4387 14467
rect 4387 14433 4396 14467
rect 4344 14424 4396 14433
rect 9496 14603 9548 14612
rect 9496 14569 9505 14603
rect 9505 14569 9539 14603
rect 9539 14569 9548 14603
rect 9496 14560 9548 14569
rect 8852 14492 8904 14544
rect 2412 14356 2464 14408
rect 2688 14356 2740 14408
rect 2320 14288 2372 14340
rect 3056 14288 3108 14340
rect 3332 14288 3384 14340
rect 5264 14356 5316 14408
rect 5356 14356 5408 14408
rect 5816 14288 5868 14340
rect 6644 14467 6696 14476
rect 6644 14433 6653 14467
rect 6653 14433 6687 14467
rect 6687 14433 6696 14467
rect 6644 14424 6696 14433
rect 8300 14424 8352 14476
rect 9680 14424 9732 14476
rect 10324 14424 10376 14476
rect 7380 14288 7432 14340
rect 8024 14288 8076 14340
rect 8944 14356 8996 14408
rect 9496 14356 9548 14408
rect 11520 14356 11572 14408
rect 10508 14288 10560 14340
rect 10784 14331 10836 14340
rect 10784 14297 10793 14331
rect 10793 14297 10827 14331
rect 10827 14297 10836 14331
rect 10784 14288 10836 14297
rect 5172 14220 5224 14272
rect 5632 14220 5684 14272
rect 7288 14220 7340 14272
rect 6378 14118 6430 14170
rect 6442 14118 6494 14170
rect 6506 14118 6558 14170
rect 6570 14118 6622 14170
rect 6634 14118 6686 14170
rect 11806 14118 11858 14170
rect 11870 14118 11922 14170
rect 11934 14118 11986 14170
rect 11998 14118 12050 14170
rect 12062 14118 12114 14170
rect 17234 14118 17286 14170
rect 17298 14118 17350 14170
rect 17362 14118 17414 14170
rect 17426 14118 17478 14170
rect 17490 14118 17542 14170
rect 22662 14118 22714 14170
rect 22726 14118 22778 14170
rect 22790 14118 22842 14170
rect 22854 14118 22906 14170
rect 22918 14118 22970 14170
rect 1860 14016 1912 14068
rect 2412 13948 2464 14000
rect 2136 13923 2188 13932
rect 2136 13889 2145 13923
rect 2145 13889 2179 13923
rect 2179 13889 2188 13923
rect 4344 13948 4396 14000
rect 2136 13880 2188 13889
rect 3424 13923 3476 13932
rect 3424 13889 3433 13923
rect 3433 13889 3467 13923
rect 3467 13889 3476 13923
rect 3424 13880 3476 13889
rect 3516 13923 3568 13932
rect 3516 13889 3525 13923
rect 3525 13889 3559 13923
rect 3559 13889 3568 13923
rect 3516 13880 3568 13889
rect 2688 13812 2740 13864
rect 4988 13948 5040 14000
rect 5448 13880 5500 13932
rect 6828 13991 6880 14000
rect 6828 13957 6837 13991
rect 6837 13957 6871 13991
rect 6871 13957 6880 13991
rect 6828 13948 6880 13957
rect 8208 13948 8260 14000
rect 4988 13812 5040 13864
rect 5356 13812 5408 13864
rect 7104 13880 7156 13932
rect 8116 13855 8168 13864
rect 8116 13821 8125 13855
rect 8125 13821 8159 13855
rect 8159 13821 8168 13855
rect 8116 13812 8168 13821
rect 8760 13923 8812 13932
rect 8760 13889 8769 13923
rect 8769 13889 8803 13923
rect 8803 13889 8812 13923
rect 8760 13880 8812 13889
rect 9496 13880 9548 13932
rect 8944 13812 8996 13864
rect 10784 13923 10836 13932
rect 10784 13889 10793 13923
rect 10793 13889 10827 13923
rect 10827 13889 10836 13923
rect 10784 13880 10836 13889
rect 13084 13923 13136 13932
rect 13084 13889 13093 13923
rect 13093 13889 13127 13923
rect 13127 13889 13136 13923
rect 13084 13880 13136 13889
rect 13268 13923 13320 13932
rect 13268 13889 13277 13923
rect 13277 13889 13311 13923
rect 13311 13889 13320 13923
rect 13268 13880 13320 13889
rect 13452 13880 13504 13932
rect 13544 13812 13596 13864
rect 13636 13855 13688 13864
rect 13636 13821 13645 13855
rect 13645 13821 13679 13855
rect 13679 13821 13688 13855
rect 13636 13812 13688 13821
rect 15200 13855 15252 13864
rect 15200 13821 15209 13855
rect 15209 13821 15243 13855
rect 15243 13821 15252 13855
rect 15200 13812 15252 13821
rect 16764 13744 16816 13796
rect 4804 13676 4856 13728
rect 10508 13676 10560 13728
rect 3664 13574 3716 13626
rect 3728 13574 3780 13626
rect 3792 13574 3844 13626
rect 3856 13574 3908 13626
rect 3920 13574 3972 13626
rect 9092 13574 9144 13626
rect 9156 13574 9208 13626
rect 9220 13574 9272 13626
rect 9284 13574 9336 13626
rect 9348 13574 9400 13626
rect 14520 13574 14572 13626
rect 14584 13574 14636 13626
rect 14648 13574 14700 13626
rect 14712 13574 14764 13626
rect 14776 13574 14828 13626
rect 19948 13574 20000 13626
rect 20012 13574 20064 13626
rect 20076 13574 20128 13626
rect 20140 13574 20192 13626
rect 20204 13574 20256 13626
rect 13268 13515 13320 13524
rect 13268 13481 13277 13515
rect 13277 13481 13311 13515
rect 13311 13481 13320 13515
rect 13268 13472 13320 13481
rect 14372 13515 14424 13524
rect 14372 13481 14381 13515
rect 14381 13481 14415 13515
rect 14415 13481 14424 13515
rect 14372 13472 14424 13481
rect 19800 13472 19852 13524
rect 15844 13404 15896 13456
rect 17592 13404 17644 13456
rect 2688 13336 2740 13388
rect 1860 13268 1912 13320
rect 3148 13311 3200 13320
rect 3148 13277 3157 13311
rect 3157 13277 3191 13311
rect 3191 13277 3200 13311
rect 3148 13268 3200 13277
rect 3608 13268 3660 13320
rect 8944 13268 8996 13320
rect 9496 13336 9548 13388
rect 13820 13336 13872 13388
rect 13912 13336 13964 13388
rect 17040 13336 17092 13388
rect 10508 13311 10560 13320
rect 10508 13277 10517 13311
rect 10517 13277 10551 13311
rect 10551 13277 10560 13311
rect 10508 13268 10560 13277
rect 10692 13311 10744 13320
rect 10692 13277 10701 13311
rect 10701 13277 10735 13311
rect 10735 13277 10744 13311
rect 10692 13268 10744 13277
rect 11612 13311 11664 13320
rect 4804 13200 4856 13252
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 10968 13200 11020 13252
rect 12440 13268 12492 13320
rect 13452 13311 13504 13320
rect 13452 13277 13461 13311
rect 13461 13277 13495 13311
rect 13495 13277 13504 13311
rect 13452 13268 13504 13277
rect 13728 13268 13780 13320
rect 14004 13268 14056 13320
rect 13268 13243 13320 13252
rect 13268 13209 13277 13243
rect 13277 13209 13311 13243
rect 13311 13209 13320 13243
rect 13268 13200 13320 13209
rect 15200 13200 15252 13252
rect 16028 13311 16080 13320
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 16488 13311 16540 13320
rect 16488 13277 16497 13311
rect 16497 13277 16531 13311
rect 16531 13277 16540 13311
rect 16488 13268 16540 13277
rect 17776 13404 17828 13456
rect 18236 13404 18288 13456
rect 2228 13132 2280 13184
rect 2964 13132 3016 13184
rect 8392 13132 8444 13184
rect 9772 13132 9824 13184
rect 15844 13175 15896 13184
rect 15844 13141 15853 13175
rect 15853 13141 15887 13175
rect 15887 13141 15896 13175
rect 15844 13132 15896 13141
rect 17684 13200 17736 13252
rect 16488 13132 16540 13184
rect 16856 13175 16908 13184
rect 16856 13141 16865 13175
rect 16865 13141 16899 13175
rect 16899 13141 16908 13175
rect 16856 13132 16908 13141
rect 18328 13132 18380 13184
rect 18512 13200 18564 13252
rect 19432 13268 19484 13320
rect 19524 13311 19576 13320
rect 19524 13277 19533 13311
rect 19533 13277 19567 13311
rect 19567 13277 19576 13311
rect 19524 13268 19576 13277
rect 19340 13200 19392 13252
rect 20628 13132 20680 13184
rect 6378 13030 6430 13082
rect 6442 13030 6494 13082
rect 6506 13030 6558 13082
rect 6570 13030 6622 13082
rect 6634 13030 6686 13082
rect 11806 13030 11858 13082
rect 11870 13030 11922 13082
rect 11934 13030 11986 13082
rect 11998 13030 12050 13082
rect 12062 13030 12114 13082
rect 17234 13030 17286 13082
rect 17298 13030 17350 13082
rect 17362 13030 17414 13082
rect 17426 13030 17478 13082
rect 17490 13030 17542 13082
rect 22662 13030 22714 13082
rect 22726 13030 22778 13082
rect 22790 13030 22842 13082
rect 22854 13030 22906 13082
rect 22918 13030 22970 13082
rect 3608 12971 3660 12980
rect 3608 12937 3617 12971
rect 3617 12937 3651 12971
rect 3651 12937 3660 12971
rect 3608 12928 3660 12937
rect 4160 12928 4212 12980
rect 2872 12860 2924 12912
rect 3424 12903 3476 12912
rect 3424 12869 3449 12903
rect 3449 12869 3476 12903
rect 3424 12860 3476 12869
rect 2688 12835 2740 12844
rect 2688 12801 2697 12835
rect 2697 12801 2731 12835
rect 2731 12801 2740 12835
rect 2688 12792 2740 12801
rect 5724 12903 5776 12912
rect 5724 12869 5733 12903
rect 5733 12869 5767 12903
rect 5767 12869 5776 12903
rect 5724 12860 5776 12869
rect 4712 12792 4764 12844
rect 4804 12835 4856 12844
rect 4804 12801 4813 12835
rect 4813 12801 4847 12835
rect 4847 12801 4856 12835
rect 8944 12928 8996 12980
rect 7932 12860 7984 12912
rect 10324 12928 10376 12980
rect 11612 12928 11664 12980
rect 12440 12971 12492 12980
rect 12440 12937 12449 12971
rect 12449 12937 12483 12971
rect 12483 12937 12492 12971
rect 12440 12928 12492 12937
rect 15384 12928 15436 12980
rect 16028 12928 16080 12980
rect 19432 12928 19484 12980
rect 4804 12792 4856 12801
rect 2228 12724 2280 12776
rect 7012 12792 7064 12844
rect 7104 12792 7156 12844
rect 8392 12835 8444 12844
rect 8392 12801 8401 12835
rect 8401 12801 8435 12835
rect 8435 12801 8444 12835
rect 8392 12792 8444 12801
rect 10324 12835 10376 12844
rect 10324 12801 10333 12835
rect 10333 12801 10367 12835
rect 10367 12801 10376 12835
rect 10324 12792 10376 12801
rect 10416 12792 10468 12844
rect 10876 12835 10928 12844
rect 10876 12801 10885 12835
rect 10885 12801 10919 12835
rect 10919 12801 10928 12835
rect 10876 12792 10928 12801
rect 10968 12835 11020 12844
rect 10968 12801 10977 12835
rect 10977 12801 11011 12835
rect 11011 12801 11020 12835
rect 10968 12792 11020 12801
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 11612 12792 11664 12844
rect 12348 12835 12400 12844
rect 12348 12801 12357 12835
rect 12357 12801 12391 12835
rect 12391 12801 12400 12835
rect 12348 12792 12400 12801
rect 12624 12792 12676 12844
rect 15108 12792 15160 12844
rect 16764 12860 16816 12912
rect 16948 12860 17000 12912
rect 3240 12588 3292 12640
rect 4620 12631 4672 12640
rect 4620 12597 4629 12631
rect 4629 12597 4663 12631
rect 4663 12597 4672 12631
rect 4620 12588 4672 12597
rect 5632 12588 5684 12640
rect 5724 12588 5776 12640
rect 8668 12767 8720 12776
rect 8668 12733 8677 12767
rect 8677 12733 8711 12767
rect 8711 12733 8720 12767
rect 8668 12724 8720 12733
rect 9588 12724 9640 12776
rect 15476 12835 15528 12844
rect 15476 12801 15485 12835
rect 15485 12801 15519 12835
rect 15519 12801 15528 12835
rect 15476 12792 15528 12801
rect 17040 12835 17092 12844
rect 17040 12801 17049 12835
rect 17049 12801 17083 12835
rect 17083 12801 17092 12835
rect 17040 12792 17092 12801
rect 17868 12792 17920 12844
rect 19524 12860 19576 12912
rect 20536 12928 20588 12980
rect 20352 12860 20404 12912
rect 18236 12835 18288 12844
rect 18236 12801 18245 12835
rect 18245 12801 18279 12835
rect 18279 12801 18288 12835
rect 18236 12792 18288 12801
rect 18328 12835 18380 12844
rect 18328 12801 18337 12835
rect 18337 12801 18371 12835
rect 18371 12801 18380 12835
rect 18328 12792 18380 12801
rect 7748 12656 7800 12708
rect 7196 12588 7248 12640
rect 7932 12588 7984 12640
rect 8208 12631 8260 12640
rect 8208 12597 8217 12631
rect 8217 12597 8251 12631
rect 8251 12597 8260 12631
rect 8208 12588 8260 12597
rect 8944 12588 8996 12640
rect 13728 12588 13780 12640
rect 15384 12767 15436 12776
rect 15384 12733 15393 12767
rect 15393 12733 15427 12767
rect 15427 12733 15436 12767
rect 15384 12724 15436 12733
rect 15844 12724 15896 12776
rect 19340 12835 19392 12844
rect 19340 12801 19349 12835
rect 19349 12801 19383 12835
rect 19383 12801 19392 12835
rect 19340 12792 19392 12801
rect 19432 12835 19484 12844
rect 19432 12801 19441 12835
rect 19441 12801 19475 12835
rect 19475 12801 19484 12835
rect 19432 12792 19484 12801
rect 18604 12724 18656 12776
rect 17684 12656 17736 12708
rect 20628 12835 20680 12844
rect 20628 12801 20637 12835
rect 20637 12801 20671 12835
rect 20671 12801 20680 12835
rect 20628 12792 20680 12801
rect 22192 12835 22244 12844
rect 22192 12801 22201 12835
rect 22201 12801 22235 12835
rect 22235 12801 22244 12835
rect 22192 12792 22244 12801
rect 20444 12724 20496 12776
rect 21732 12724 21784 12776
rect 16028 12588 16080 12640
rect 17224 12588 17276 12640
rect 18144 12588 18196 12640
rect 19524 12631 19576 12640
rect 19524 12597 19533 12631
rect 19533 12597 19567 12631
rect 19567 12597 19576 12631
rect 19524 12588 19576 12597
rect 3664 12486 3716 12538
rect 3728 12486 3780 12538
rect 3792 12486 3844 12538
rect 3856 12486 3908 12538
rect 3920 12486 3972 12538
rect 9092 12486 9144 12538
rect 9156 12486 9208 12538
rect 9220 12486 9272 12538
rect 9284 12486 9336 12538
rect 9348 12486 9400 12538
rect 14520 12486 14572 12538
rect 14584 12486 14636 12538
rect 14648 12486 14700 12538
rect 14712 12486 14764 12538
rect 14776 12486 14828 12538
rect 19948 12486 20000 12538
rect 20012 12486 20064 12538
rect 20076 12486 20128 12538
rect 20140 12486 20192 12538
rect 20204 12486 20256 12538
rect 3148 12427 3200 12436
rect 3148 12393 3157 12427
rect 3157 12393 3191 12427
rect 3191 12393 3200 12427
rect 3148 12384 3200 12393
rect 7012 12427 7064 12436
rect 7012 12393 7021 12427
rect 7021 12393 7055 12427
rect 7055 12393 7064 12427
rect 7012 12384 7064 12393
rect 7748 12427 7800 12436
rect 7748 12393 7757 12427
rect 7757 12393 7791 12427
rect 7791 12393 7800 12427
rect 7748 12384 7800 12393
rect 10692 12384 10744 12436
rect 13084 12427 13136 12436
rect 13084 12393 13093 12427
rect 13093 12393 13127 12427
rect 13127 12393 13136 12427
rect 13084 12384 13136 12393
rect 13176 12384 13228 12436
rect 13544 12384 13596 12436
rect 13636 12384 13688 12436
rect 17868 12384 17920 12436
rect 18604 12384 18656 12436
rect 21088 12384 21140 12436
rect 2872 12316 2924 12368
rect 2780 12248 2832 12300
rect 2136 12223 2188 12232
rect 2136 12189 2145 12223
rect 2145 12189 2179 12223
rect 2179 12189 2188 12223
rect 2136 12180 2188 12189
rect 2504 12180 2556 12232
rect 4712 12291 4764 12300
rect 4712 12257 4721 12291
rect 4721 12257 4755 12291
rect 4755 12257 4764 12291
rect 4712 12248 4764 12257
rect 5724 12248 5776 12300
rect 3424 12180 3476 12232
rect 3148 12155 3200 12164
rect 3148 12121 3157 12155
rect 3157 12121 3191 12155
rect 3191 12121 3200 12155
rect 3148 12112 3200 12121
rect 5632 12223 5684 12232
rect 5632 12189 5641 12223
rect 5641 12189 5675 12223
rect 5675 12189 5684 12223
rect 5632 12180 5684 12189
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 2872 12044 2924 12096
rect 4252 12087 4304 12096
rect 4252 12053 4261 12087
rect 4261 12053 4295 12087
rect 4295 12053 4304 12087
rect 4252 12044 4304 12053
rect 5356 12044 5408 12096
rect 9864 12316 9916 12368
rect 11520 12316 11572 12368
rect 8944 12248 8996 12300
rect 10324 12291 10376 12300
rect 10324 12257 10333 12291
rect 10333 12257 10367 12291
rect 10367 12257 10376 12291
rect 10324 12248 10376 12257
rect 7932 12223 7984 12232
rect 7932 12189 7941 12223
rect 7941 12189 7975 12223
rect 7975 12189 7984 12223
rect 7932 12180 7984 12189
rect 7104 12112 7156 12164
rect 9588 12180 9640 12232
rect 11152 12248 11204 12300
rect 13728 12248 13780 12300
rect 10876 12180 10928 12232
rect 13360 12223 13412 12232
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 13452 12223 13504 12232
rect 13452 12189 13461 12223
rect 13461 12189 13495 12223
rect 13495 12189 13504 12223
rect 13452 12180 13504 12189
rect 16764 12316 16816 12368
rect 19708 12316 19760 12368
rect 19800 12316 19852 12368
rect 20720 12316 20772 12368
rect 16856 12248 16908 12300
rect 13912 12180 13964 12232
rect 14924 12180 14976 12232
rect 10416 12155 10468 12164
rect 10416 12121 10425 12155
rect 10425 12121 10459 12155
rect 10459 12121 10468 12155
rect 10416 12112 10468 12121
rect 15384 12223 15436 12232
rect 15384 12189 15393 12223
rect 15393 12189 15427 12223
rect 15427 12189 15436 12223
rect 15384 12180 15436 12189
rect 16488 12180 16540 12232
rect 16580 12223 16632 12232
rect 16580 12189 16589 12223
rect 16589 12189 16623 12223
rect 16623 12189 16632 12223
rect 16580 12180 16632 12189
rect 16672 12180 16724 12232
rect 17224 12223 17276 12232
rect 17224 12189 17233 12223
rect 17233 12189 17267 12223
rect 17267 12189 17276 12223
rect 17224 12180 17276 12189
rect 17316 12180 17368 12232
rect 17684 12223 17736 12232
rect 17684 12189 17693 12223
rect 17693 12189 17727 12223
rect 17727 12189 17736 12223
rect 17684 12180 17736 12189
rect 20168 12248 20220 12300
rect 20444 12291 20496 12300
rect 20444 12257 20453 12291
rect 20453 12257 20487 12291
rect 20487 12257 20496 12291
rect 20444 12248 20496 12257
rect 20996 12248 21048 12300
rect 19340 12180 19392 12232
rect 20352 12223 20404 12232
rect 20352 12189 20361 12223
rect 20361 12189 20395 12223
rect 20395 12189 20404 12223
rect 20352 12180 20404 12189
rect 20720 12180 20772 12232
rect 20812 12180 20864 12232
rect 21732 12223 21784 12232
rect 21732 12189 21741 12223
rect 21741 12189 21775 12223
rect 21775 12189 21784 12223
rect 21732 12180 21784 12189
rect 6276 12044 6328 12096
rect 8484 12044 8536 12096
rect 8760 12044 8812 12096
rect 11612 12044 11664 12096
rect 11704 12044 11756 12096
rect 12348 12044 12400 12096
rect 13544 12044 13596 12096
rect 15752 12087 15804 12096
rect 15752 12053 15761 12087
rect 15761 12053 15795 12087
rect 15795 12053 15804 12087
rect 15752 12044 15804 12053
rect 17684 12044 17736 12096
rect 18696 12044 18748 12096
rect 20076 12087 20128 12096
rect 20076 12053 20085 12087
rect 20085 12053 20119 12087
rect 20119 12053 20128 12087
rect 20076 12044 20128 12053
rect 21272 12044 21324 12096
rect 6378 11942 6430 11994
rect 6442 11942 6494 11994
rect 6506 11942 6558 11994
rect 6570 11942 6622 11994
rect 6634 11942 6686 11994
rect 11806 11942 11858 11994
rect 11870 11942 11922 11994
rect 11934 11942 11986 11994
rect 11998 11942 12050 11994
rect 12062 11942 12114 11994
rect 17234 11942 17286 11994
rect 17298 11942 17350 11994
rect 17362 11942 17414 11994
rect 17426 11942 17478 11994
rect 17490 11942 17542 11994
rect 22662 11942 22714 11994
rect 22726 11942 22778 11994
rect 22790 11942 22842 11994
rect 22854 11942 22906 11994
rect 22918 11942 22970 11994
rect 15384 11840 15436 11892
rect 16580 11840 16632 11892
rect 17500 11840 17552 11892
rect 17776 11840 17828 11892
rect 2504 11772 2556 11824
rect 2228 11704 2280 11756
rect 2780 11704 2832 11756
rect 4160 11704 4212 11756
rect 4620 11747 4672 11756
rect 4620 11713 4629 11747
rect 4629 11713 4663 11747
rect 4663 11713 4672 11747
rect 4620 11704 4672 11713
rect 16764 11704 16816 11756
rect 16856 11704 16908 11756
rect 4344 11679 4396 11688
rect 4344 11645 4353 11679
rect 4353 11645 4387 11679
rect 4387 11645 4396 11679
rect 4344 11636 4396 11645
rect 2136 11611 2188 11620
rect 2136 11577 2145 11611
rect 2145 11577 2179 11611
rect 2179 11577 2188 11611
rect 2136 11568 2188 11577
rect 4804 11543 4856 11552
rect 4804 11509 4813 11543
rect 4813 11509 4847 11543
rect 4847 11509 4856 11543
rect 4804 11500 4856 11509
rect 14924 11500 14976 11552
rect 16488 11636 16540 11688
rect 17408 11747 17460 11756
rect 17408 11713 17417 11747
rect 17417 11713 17451 11747
rect 17451 11713 17460 11747
rect 17408 11704 17460 11713
rect 17684 11704 17736 11756
rect 20812 11840 20864 11892
rect 19524 11772 19576 11824
rect 20076 11815 20128 11824
rect 20076 11781 20085 11815
rect 20085 11781 20119 11815
rect 20119 11781 20128 11815
rect 20076 11772 20128 11781
rect 20996 11704 21048 11756
rect 15936 11568 15988 11620
rect 19524 11636 19576 11688
rect 18236 11568 18288 11620
rect 19340 11568 19392 11620
rect 20720 11636 20772 11688
rect 17868 11500 17920 11552
rect 19616 11500 19668 11552
rect 21180 11543 21232 11552
rect 21180 11509 21189 11543
rect 21189 11509 21223 11543
rect 21223 11509 21232 11543
rect 21180 11500 21232 11509
rect 3664 11398 3716 11450
rect 3728 11398 3780 11450
rect 3792 11398 3844 11450
rect 3856 11398 3908 11450
rect 3920 11398 3972 11450
rect 9092 11398 9144 11450
rect 9156 11398 9208 11450
rect 9220 11398 9272 11450
rect 9284 11398 9336 11450
rect 9348 11398 9400 11450
rect 14520 11398 14572 11450
rect 14584 11398 14636 11450
rect 14648 11398 14700 11450
rect 14712 11398 14764 11450
rect 14776 11398 14828 11450
rect 19948 11398 20000 11450
rect 20012 11398 20064 11450
rect 20076 11398 20128 11450
rect 20140 11398 20192 11450
rect 20204 11398 20256 11450
rect 6276 11296 6328 11348
rect 7104 11296 7156 11348
rect 14556 11296 14608 11348
rect 15384 11296 15436 11348
rect 17408 11296 17460 11348
rect 21272 11339 21324 11348
rect 21272 11305 21281 11339
rect 21281 11305 21315 11339
rect 21315 11305 21324 11339
rect 21272 11296 21324 11305
rect 1860 11271 1912 11280
rect 1860 11237 1869 11271
rect 1869 11237 1903 11271
rect 1903 11237 1912 11271
rect 1860 11228 1912 11237
rect 940 11092 992 11144
rect 4160 11092 4212 11144
rect 5356 11135 5408 11144
rect 5356 11101 5390 11135
rect 5390 11101 5408 11135
rect 5356 11092 5408 11101
rect 6920 11135 6972 11144
rect 6920 11101 6929 11135
rect 6929 11101 6963 11135
rect 6963 11101 6972 11135
rect 6920 11092 6972 11101
rect 7196 11135 7248 11144
rect 7196 11101 7230 11135
rect 7230 11101 7248 11135
rect 7196 11092 7248 11101
rect 14188 11228 14240 11280
rect 14280 11160 14332 11212
rect 16396 11228 16448 11280
rect 21180 11271 21232 11280
rect 21180 11237 21189 11271
rect 21189 11237 21223 11271
rect 21223 11237 21232 11271
rect 21180 11228 21232 11237
rect 15660 11160 15712 11212
rect 13728 11135 13780 11144
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 13728 11092 13780 11101
rect 14464 11135 14516 11144
rect 14464 11101 14473 11135
rect 14473 11101 14507 11135
rect 14507 11101 14516 11135
rect 14464 11092 14516 11101
rect 14556 11135 14608 11144
rect 14556 11101 14565 11135
rect 14565 11101 14599 11135
rect 14599 11101 14608 11135
rect 14556 11092 14608 11101
rect 14004 11024 14056 11076
rect 14188 11024 14240 11076
rect 14924 11092 14976 11144
rect 15476 11135 15528 11144
rect 15476 11101 15485 11135
rect 15485 11101 15519 11135
rect 15519 11101 15528 11135
rect 15476 11092 15528 11101
rect 15292 11067 15344 11076
rect 15292 11033 15301 11067
rect 15301 11033 15335 11067
rect 15335 11033 15344 11067
rect 15292 11024 15344 11033
rect 15752 11135 15804 11144
rect 15752 11101 15761 11135
rect 15761 11101 15795 11135
rect 15795 11101 15804 11135
rect 15752 11092 15804 11101
rect 16672 11092 16724 11144
rect 16764 11135 16816 11144
rect 16764 11101 16773 11135
rect 16773 11101 16807 11135
rect 16807 11101 16816 11135
rect 16764 11092 16816 11101
rect 17684 11203 17736 11212
rect 17684 11169 17693 11203
rect 17693 11169 17727 11203
rect 17727 11169 17736 11203
rect 17684 11160 17736 11169
rect 17868 11203 17920 11212
rect 17868 11169 17877 11203
rect 17877 11169 17911 11203
rect 17911 11169 17920 11203
rect 17868 11160 17920 11169
rect 18144 11203 18196 11212
rect 18144 11169 18153 11203
rect 18153 11169 18187 11203
rect 18187 11169 18196 11203
rect 18144 11160 18196 11169
rect 17776 11092 17828 11144
rect 17960 11135 18012 11144
rect 17960 11101 17969 11135
rect 17969 11101 18003 11135
rect 18003 11101 18012 11135
rect 17960 11092 18012 11101
rect 18236 11092 18288 11144
rect 18696 11135 18748 11144
rect 18696 11101 18705 11135
rect 18705 11101 18739 11135
rect 18739 11101 18748 11135
rect 18696 11092 18748 11101
rect 18880 11135 18932 11144
rect 18880 11101 18889 11135
rect 18889 11101 18923 11135
rect 18923 11101 18932 11135
rect 18880 11092 18932 11101
rect 16488 11067 16540 11076
rect 16488 11033 16497 11067
rect 16497 11033 16531 11067
rect 16531 11033 16540 11067
rect 16488 11024 16540 11033
rect 16856 11024 16908 11076
rect 17868 11024 17920 11076
rect 19800 11160 19852 11212
rect 19616 11135 19668 11144
rect 19616 11101 19625 11135
rect 19625 11101 19659 11135
rect 19659 11101 19668 11135
rect 19616 11092 19668 11101
rect 19708 11135 19760 11144
rect 19708 11101 19717 11135
rect 19717 11101 19751 11135
rect 19751 11101 19760 11135
rect 19708 11092 19760 11101
rect 13176 10999 13228 11008
rect 13176 10965 13185 10999
rect 13185 10965 13219 10999
rect 13219 10965 13228 10999
rect 13176 10956 13228 10965
rect 13912 10956 13964 11008
rect 16672 10956 16724 11008
rect 17500 10956 17552 11008
rect 17776 10956 17828 11008
rect 19800 11067 19852 11076
rect 19800 11033 19809 11067
rect 19809 11033 19843 11067
rect 19843 11033 19852 11067
rect 19800 11024 19852 11033
rect 21088 11135 21140 11144
rect 21088 11101 21097 11135
rect 21097 11101 21131 11135
rect 21131 11101 21140 11135
rect 21088 11092 21140 11101
rect 21180 11092 21232 11144
rect 22008 11092 22060 11144
rect 20444 11024 20496 11076
rect 19248 10956 19300 11008
rect 6378 10854 6430 10906
rect 6442 10854 6494 10906
rect 6506 10854 6558 10906
rect 6570 10854 6622 10906
rect 6634 10854 6686 10906
rect 11806 10854 11858 10906
rect 11870 10854 11922 10906
rect 11934 10854 11986 10906
rect 11998 10854 12050 10906
rect 12062 10854 12114 10906
rect 17234 10854 17286 10906
rect 17298 10854 17350 10906
rect 17362 10854 17414 10906
rect 17426 10854 17478 10906
rect 17490 10854 17542 10906
rect 22662 10854 22714 10906
rect 22726 10854 22778 10906
rect 22790 10854 22842 10906
rect 22854 10854 22906 10906
rect 22918 10854 22970 10906
rect 2780 10752 2832 10804
rect 4896 10752 4948 10804
rect 8668 10752 8720 10804
rect 10876 10795 10928 10804
rect 10876 10761 10885 10795
rect 10885 10761 10919 10795
rect 10919 10761 10928 10795
rect 10876 10752 10928 10761
rect 1952 10727 2004 10736
rect 1952 10693 1986 10727
rect 1986 10693 2004 10727
rect 1952 10684 2004 10693
rect 5540 10684 5592 10736
rect 8208 10684 8260 10736
rect 9772 10727 9824 10736
rect 9772 10693 9806 10727
rect 9806 10693 9824 10727
rect 9772 10684 9824 10693
rect 6920 10616 6972 10668
rect 1676 10591 1728 10600
rect 1676 10557 1685 10591
rect 1685 10557 1719 10591
rect 1719 10557 1728 10591
rect 1676 10548 1728 10557
rect 6736 10548 6788 10600
rect 9496 10591 9548 10600
rect 9496 10557 9505 10591
rect 9505 10557 9539 10591
rect 9539 10557 9548 10591
rect 9496 10548 9548 10557
rect 12164 10659 12216 10668
rect 12164 10625 12173 10659
rect 12173 10625 12207 10659
rect 12207 10625 12216 10659
rect 12164 10616 12216 10625
rect 13728 10752 13780 10804
rect 14464 10752 14516 10804
rect 15476 10752 15528 10804
rect 16028 10752 16080 10804
rect 13176 10684 13228 10736
rect 16672 10684 16724 10736
rect 13912 10616 13964 10668
rect 15936 10616 15988 10668
rect 16212 10659 16264 10668
rect 16212 10625 16221 10659
rect 16221 10625 16255 10659
rect 16255 10625 16264 10659
rect 16212 10616 16264 10625
rect 16948 10616 17000 10668
rect 19340 10752 19392 10804
rect 19432 10752 19484 10804
rect 19616 10752 19668 10804
rect 20996 10795 21048 10804
rect 20996 10761 21005 10795
rect 21005 10761 21039 10795
rect 21039 10761 21048 10795
rect 20996 10752 21048 10761
rect 17960 10684 18012 10736
rect 12348 10548 12400 10600
rect 12900 10591 12952 10600
rect 12900 10557 12909 10591
rect 12909 10557 12943 10591
rect 12943 10557 12952 10591
rect 12900 10548 12952 10557
rect 13084 10480 13136 10532
rect 14004 10591 14056 10600
rect 14004 10557 14013 10591
rect 14013 10557 14047 10591
rect 14047 10557 14056 10591
rect 15016 10591 15068 10600
rect 14004 10548 14056 10557
rect 15016 10557 15025 10591
rect 15025 10557 15059 10591
rect 15059 10557 15068 10591
rect 15016 10548 15068 10557
rect 15108 10591 15160 10600
rect 15108 10557 15117 10591
rect 15117 10557 15151 10591
rect 15151 10557 15160 10591
rect 15108 10548 15160 10557
rect 16304 10548 16356 10600
rect 14188 10480 14240 10532
rect 16948 10480 17000 10532
rect 17408 10616 17460 10668
rect 19432 10659 19484 10668
rect 19432 10625 19441 10659
rect 19441 10625 19475 10659
rect 19475 10625 19484 10659
rect 19432 10616 19484 10625
rect 17868 10548 17920 10600
rect 18420 10591 18472 10600
rect 18420 10557 18429 10591
rect 18429 10557 18463 10591
rect 18463 10557 18472 10591
rect 18420 10548 18472 10557
rect 18880 10548 18932 10600
rect 19708 10659 19760 10668
rect 19708 10625 19717 10659
rect 19717 10625 19751 10659
rect 19751 10625 19760 10659
rect 19708 10616 19760 10625
rect 19616 10548 19668 10600
rect 20628 10616 20680 10668
rect 22192 10659 22244 10668
rect 22192 10625 22201 10659
rect 22201 10625 22235 10659
rect 22235 10625 22244 10659
rect 22192 10616 22244 10625
rect 21272 10548 21324 10600
rect 21548 10548 21600 10600
rect 11244 10412 11296 10464
rect 13268 10412 13320 10464
rect 16764 10412 16816 10464
rect 17408 10412 17460 10464
rect 17500 10455 17552 10464
rect 17500 10421 17509 10455
rect 17509 10421 17543 10455
rect 17543 10421 17552 10455
rect 17500 10412 17552 10421
rect 17868 10412 17920 10464
rect 22008 10455 22060 10464
rect 22008 10421 22017 10455
rect 22017 10421 22051 10455
rect 22051 10421 22060 10455
rect 22008 10412 22060 10421
rect 3664 10310 3716 10362
rect 3728 10310 3780 10362
rect 3792 10310 3844 10362
rect 3856 10310 3908 10362
rect 3920 10310 3972 10362
rect 9092 10310 9144 10362
rect 9156 10310 9208 10362
rect 9220 10310 9272 10362
rect 9284 10310 9336 10362
rect 9348 10310 9400 10362
rect 14520 10310 14572 10362
rect 14584 10310 14636 10362
rect 14648 10310 14700 10362
rect 14712 10310 14764 10362
rect 14776 10310 14828 10362
rect 19948 10310 20000 10362
rect 20012 10310 20064 10362
rect 20076 10310 20128 10362
rect 20140 10310 20192 10362
rect 20204 10310 20256 10362
rect 2412 10208 2464 10260
rect 5080 10208 5132 10260
rect 8484 10251 8536 10260
rect 8484 10217 8493 10251
rect 8493 10217 8527 10251
rect 8527 10217 8536 10251
rect 8484 10208 8536 10217
rect 9680 10208 9732 10260
rect 12900 10208 12952 10260
rect 13636 10208 13688 10260
rect 15660 10251 15712 10260
rect 15660 10217 15669 10251
rect 15669 10217 15703 10251
rect 15703 10217 15712 10251
rect 15660 10208 15712 10217
rect 16212 10208 16264 10260
rect 19616 10251 19668 10260
rect 19616 10217 19625 10251
rect 19625 10217 19659 10251
rect 19659 10217 19668 10251
rect 19616 10208 19668 10217
rect 19800 10208 19852 10260
rect 20536 10208 20588 10260
rect 4160 10115 4212 10124
rect 4160 10081 4169 10115
rect 4169 10081 4203 10115
rect 4203 10081 4212 10115
rect 4160 10072 4212 10081
rect 6736 10072 6788 10124
rect 17500 10140 17552 10192
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 1768 10004 1820 10056
rect 4436 10047 4488 10056
rect 4436 10013 4470 10047
rect 4470 10013 4488 10047
rect 4436 10004 4488 10013
rect 16948 10072 17000 10124
rect 19708 10115 19760 10124
rect 19708 10081 19717 10115
rect 19717 10081 19751 10115
rect 19751 10081 19760 10115
rect 19708 10072 19760 10081
rect 9496 10047 9548 10056
rect 9496 10013 9505 10047
rect 9505 10013 9539 10047
rect 9539 10013 9548 10047
rect 9496 10004 9548 10013
rect 10968 10004 11020 10056
rect 13084 10047 13136 10056
rect 13084 10013 13090 10047
rect 13090 10013 13124 10047
rect 13124 10013 13136 10047
rect 13084 10004 13136 10013
rect 8116 9936 8168 9988
rect 12348 9936 12400 9988
rect 16672 10004 16724 10056
rect 16764 10004 16816 10056
rect 17592 10004 17644 10056
rect 19800 10004 19852 10056
rect 20352 10004 20404 10056
rect 15108 9936 15160 9988
rect 21272 9936 21324 9988
rect 12716 9868 12768 9920
rect 13084 9911 13136 9920
rect 13084 9877 13093 9911
rect 13093 9877 13127 9911
rect 13127 9877 13136 9911
rect 13084 9868 13136 9877
rect 16028 9911 16080 9920
rect 16028 9877 16037 9911
rect 16037 9877 16071 9911
rect 16071 9877 16080 9911
rect 16028 9868 16080 9877
rect 16212 9868 16264 9920
rect 20260 9868 20312 9920
rect 20720 9868 20772 9920
rect 6378 9766 6430 9818
rect 6442 9766 6494 9818
rect 6506 9766 6558 9818
rect 6570 9766 6622 9818
rect 6634 9766 6686 9818
rect 11806 9766 11858 9818
rect 11870 9766 11922 9818
rect 11934 9766 11986 9818
rect 11998 9766 12050 9818
rect 12062 9766 12114 9818
rect 17234 9766 17286 9818
rect 17298 9766 17350 9818
rect 17362 9766 17414 9818
rect 17426 9766 17478 9818
rect 17490 9766 17542 9818
rect 22662 9766 22714 9818
rect 22726 9766 22778 9818
rect 22790 9766 22842 9818
rect 22854 9766 22906 9818
rect 22918 9766 22970 9818
rect 9772 9664 9824 9716
rect 12164 9664 12216 9716
rect 14188 9664 14240 9716
rect 15016 9664 15068 9716
rect 16488 9664 16540 9716
rect 16948 9707 17000 9716
rect 16948 9673 16957 9707
rect 16957 9673 16991 9707
rect 16991 9673 17000 9707
rect 16948 9664 17000 9673
rect 17132 9664 17184 9716
rect 17684 9664 17736 9716
rect 17868 9664 17920 9716
rect 19248 9664 19300 9716
rect 20628 9664 20680 9716
rect 1676 9596 1728 9648
rect 2872 9596 2924 9648
rect 9864 9639 9916 9648
rect 9864 9605 9898 9639
rect 9898 9605 9916 9639
rect 9864 9596 9916 9605
rect 2044 9571 2096 9580
rect 2044 9537 2078 9571
rect 2078 9537 2096 9571
rect 2044 9528 2096 9537
rect 4160 9528 4212 9580
rect 4528 9571 4580 9580
rect 4528 9537 4562 9571
rect 4562 9537 4580 9571
rect 4528 9528 4580 9537
rect 9496 9528 9548 9580
rect 16488 9528 16540 9580
rect 16856 9571 16908 9580
rect 16856 9537 16865 9571
rect 16865 9537 16899 9571
rect 16899 9537 16908 9571
rect 16856 9528 16908 9537
rect 17592 9596 17644 9648
rect 17224 9528 17276 9580
rect 17776 9571 17828 9580
rect 17776 9537 17785 9571
rect 17785 9537 17819 9571
rect 17819 9537 17828 9571
rect 17776 9528 17828 9537
rect 17868 9528 17920 9580
rect 3056 9392 3108 9444
rect 5264 9392 5316 9444
rect 11704 9392 11756 9444
rect 17684 9392 17736 9444
rect 17776 9324 17828 9376
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 18420 9460 18472 9512
rect 18788 9571 18840 9580
rect 18788 9537 18797 9571
rect 18797 9537 18831 9571
rect 18831 9537 18840 9571
rect 18788 9528 18840 9537
rect 20720 9528 20772 9580
rect 20996 9596 21048 9648
rect 21548 9596 21600 9648
rect 18512 9435 18564 9444
rect 18512 9401 18521 9435
rect 18521 9401 18555 9435
rect 18555 9401 18564 9435
rect 18512 9392 18564 9401
rect 20260 9392 20312 9444
rect 20628 9392 20680 9444
rect 21272 9571 21324 9580
rect 21272 9537 21286 9571
rect 21286 9537 21320 9571
rect 21320 9537 21324 9571
rect 21272 9528 21324 9537
rect 22100 9528 22152 9580
rect 20720 9324 20772 9376
rect 21088 9324 21140 9376
rect 21272 9324 21324 9376
rect 22008 9367 22060 9376
rect 22008 9333 22017 9367
rect 22017 9333 22051 9367
rect 22051 9333 22060 9367
rect 22008 9324 22060 9333
rect 3664 9222 3716 9274
rect 3728 9222 3780 9274
rect 3792 9222 3844 9274
rect 3856 9222 3908 9274
rect 3920 9222 3972 9274
rect 9092 9222 9144 9274
rect 9156 9222 9208 9274
rect 9220 9222 9272 9274
rect 9284 9222 9336 9274
rect 9348 9222 9400 9274
rect 14520 9222 14572 9274
rect 14584 9222 14636 9274
rect 14648 9222 14700 9274
rect 14712 9222 14764 9274
rect 14776 9222 14828 9274
rect 19948 9222 20000 9274
rect 20012 9222 20064 9274
rect 20076 9222 20128 9274
rect 20140 9222 20192 9274
rect 20204 9222 20256 9274
rect 3332 9120 3384 9172
rect 11060 9120 11112 9172
rect 13084 9163 13136 9172
rect 13084 9129 13093 9163
rect 13093 9129 13127 9163
rect 13127 9129 13136 9163
rect 13084 9120 13136 9129
rect 15108 9120 15160 9172
rect 19340 9120 19392 9172
rect 1676 8984 1728 9036
rect 9496 9027 9548 9036
rect 9496 8993 9505 9027
rect 9505 8993 9539 9027
rect 9539 8993 9548 9027
rect 9496 8984 9548 8993
rect 2596 8916 2648 8968
rect 16580 9052 16632 9104
rect 20444 9052 20496 9104
rect 12808 8984 12860 9036
rect 13360 8916 13412 8968
rect 14924 8916 14976 8968
rect 16764 8984 16816 9036
rect 16948 8984 17000 9036
rect 18236 8984 18288 9036
rect 13268 8848 13320 8900
rect 13544 8848 13596 8900
rect 16488 8916 16540 8968
rect 16948 8848 17000 8900
rect 17592 8959 17644 8968
rect 17592 8925 17601 8959
rect 17601 8925 17635 8959
rect 17635 8925 17644 8959
rect 17592 8916 17644 8925
rect 19248 8916 19300 8968
rect 17684 8848 17736 8900
rect 18788 8848 18840 8900
rect 22008 8984 22060 9036
rect 21180 8916 21232 8968
rect 21272 8959 21324 8968
rect 21272 8925 21281 8959
rect 21281 8925 21315 8959
rect 21315 8925 21324 8959
rect 21272 8916 21324 8925
rect 15016 8780 15068 8832
rect 16212 8823 16264 8832
rect 16212 8789 16221 8823
rect 16221 8789 16255 8823
rect 16255 8789 16264 8823
rect 16212 8780 16264 8789
rect 16856 8780 16908 8832
rect 17224 8780 17276 8832
rect 17592 8780 17644 8832
rect 19340 8780 19392 8832
rect 20628 8823 20680 8832
rect 20628 8789 20637 8823
rect 20637 8789 20671 8823
rect 20671 8789 20680 8823
rect 20628 8780 20680 8789
rect 6378 8678 6430 8730
rect 6442 8678 6494 8730
rect 6506 8678 6558 8730
rect 6570 8678 6622 8730
rect 6634 8678 6686 8730
rect 11806 8678 11858 8730
rect 11870 8678 11922 8730
rect 11934 8678 11986 8730
rect 11998 8678 12050 8730
rect 12062 8678 12114 8730
rect 17234 8678 17286 8730
rect 17298 8678 17350 8730
rect 17362 8678 17414 8730
rect 17426 8678 17478 8730
rect 17490 8678 17542 8730
rect 22662 8678 22714 8730
rect 22726 8678 22778 8730
rect 22790 8678 22842 8730
rect 22854 8678 22906 8730
rect 22918 8678 22970 8730
rect 4344 8619 4396 8628
rect 4344 8585 4353 8619
rect 4353 8585 4387 8619
rect 4387 8585 4396 8619
rect 4344 8576 4396 8585
rect 8024 8619 8076 8628
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 10784 8576 10836 8628
rect 12808 8619 12860 8628
rect 12808 8585 12817 8619
rect 12817 8585 12851 8619
rect 12851 8585 12860 8619
rect 12808 8576 12860 8585
rect 13360 8619 13412 8628
rect 13360 8585 13369 8619
rect 13369 8585 13403 8619
rect 13403 8585 13412 8619
rect 13360 8576 13412 8585
rect 15292 8576 15344 8628
rect 4804 8508 4856 8560
rect 7288 8508 7340 8560
rect 6736 8440 6788 8492
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 11244 8440 11296 8492
rect 12256 8440 12308 8492
rect 13728 8440 13780 8492
rect 17592 8576 17644 8628
rect 18052 8576 18104 8628
rect 19524 8619 19576 8628
rect 19524 8585 19533 8619
rect 19533 8585 19567 8619
rect 19567 8585 19576 8619
rect 19524 8576 19576 8585
rect 20444 8619 20496 8628
rect 20444 8585 20453 8619
rect 20453 8585 20487 8619
rect 20487 8585 20496 8619
rect 20444 8576 20496 8585
rect 15752 8508 15804 8560
rect 13544 8415 13596 8424
rect 13544 8381 13553 8415
rect 13553 8381 13587 8415
rect 13587 8381 13596 8415
rect 13544 8372 13596 8381
rect 13912 8415 13964 8424
rect 13912 8381 13921 8415
rect 13921 8381 13955 8415
rect 13955 8381 13964 8415
rect 13912 8372 13964 8381
rect 14188 8372 14240 8424
rect 15384 8440 15436 8492
rect 15844 8483 15896 8492
rect 15844 8449 15853 8483
rect 15853 8449 15887 8483
rect 15887 8449 15896 8483
rect 15844 8440 15896 8449
rect 16488 8508 16540 8560
rect 16856 8483 16908 8492
rect 16856 8449 16865 8483
rect 16865 8449 16899 8483
rect 16899 8449 16908 8483
rect 16856 8440 16908 8449
rect 17500 8483 17552 8492
rect 17500 8449 17509 8483
rect 17509 8449 17543 8483
rect 17543 8449 17552 8483
rect 17500 8440 17552 8449
rect 17684 8440 17736 8492
rect 15108 8372 15160 8424
rect 15476 8372 15528 8424
rect 16948 8415 17000 8424
rect 16948 8381 16957 8415
rect 16957 8381 16991 8415
rect 16991 8381 17000 8415
rect 16948 8372 17000 8381
rect 17408 8372 17460 8424
rect 19156 8483 19208 8492
rect 19156 8449 19165 8483
rect 19165 8449 19199 8483
rect 19199 8449 19208 8483
rect 19156 8440 19208 8449
rect 19340 8440 19392 8492
rect 20720 8508 20772 8560
rect 20812 8551 20864 8560
rect 20812 8517 20821 8551
rect 20821 8517 20855 8551
rect 20855 8517 20864 8551
rect 20812 8508 20864 8517
rect 19708 8372 19760 8424
rect 20536 8372 20588 8424
rect 17960 8304 18012 8356
rect 14924 8236 14976 8288
rect 15752 8236 15804 8288
rect 15936 8279 15988 8288
rect 15936 8245 15945 8279
rect 15945 8245 15979 8279
rect 15979 8245 15988 8279
rect 15936 8236 15988 8245
rect 17592 8279 17644 8288
rect 17592 8245 17601 8279
rect 17601 8245 17635 8279
rect 17635 8245 17644 8279
rect 17592 8236 17644 8245
rect 20536 8236 20588 8288
rect 3664 8134 3716 8186
rect 3728 8134 3780 8186
rect 3792 8134 3844 8186
rect 3856 8134 3908 8186
rect 3920 8134 3972 8186
rect 9092 8134 9144 8186
rect 9156 8134 9208 8186
rect 9220 8134 9272 8186
rect 9284 8134 9336 8186
rect 9348 8134 9400 8186
rect 14520 8134 14572 8186
rect 14584 8134 14636 8186
rect 14648 8134 14700 8186
rect 14712 8134 14764 8186
rect 14776 8134 14828 8186
rect 19948 8134 20000 8186
rect 20012 8134 20064 8186
rect 20076 8134 20128 8186
rect 20140 8134 20192 8186
rect 20204 8134 20256 8186
rect 13452 8032 13504 8084
rect 15108 8032 15160 8084
rect 15476 8032 15528 8084
rect 15752 8032 15804 8084
rect 17316 8032 17368 8084
rect 17592 8032 17644 8084
rect 19432 8032 19484 8084
rect 12624 7964 12676 8016
rect 13360 7964 13412 8016
rect 16212 7964 16264 8016
rect 9496 7896 9548 7948
rect 2228 7828 2280 7880
rect 2504 7871 2556 7880
rect 2504 7837 2513 7871
rect 2513 7837 2547 7871
rect 2547 7837 2556 7871
rect 2504 7828 2556 7837
rect 12164 7828 12216 7880
rect 14924 7896 14976 7948
rect 13268 7871 13320 7880
rect 13268 7837 13277 7871
rect 13277 7837 13311 7871
rect 13311 7837 13320 7871
rect 13268 7828 13320 7837
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 15292 7939 15344 7948
rect 15292 7905 15301 7939
rect 15301 7905 15335 7939
rect 15335 7905 15344 7939
rect 15292 7896 15344 7905
rect 15844 7896 15896 7948
rect 16948 7896 17000 7948
rect 17408 7896 17460 7948
rect 20352 7828 20404 7880
rect 20996 7964 21048 8016
rect 2688 7760 2740 7812
rect 5540 7760 5592 7812
rect 2412 7735 2464 7744
rect 2412 7701 2421 7735
rect 2421 7701 2455 7735
rect 2455 7701 2464 7735
rect 2412 7692 2464 7701
rect 4344 7692 4396 7744
rect 7840 7760 7892 7812
rect 12348 7760 12400 7812
rect 12808 7760 12860 7812
rect 20444 7760 20496 7812
rect 12900 7692 12952 7744
rect 13452 7692 13504 7744
rect 15108 7692 15160 7744
rect 18144 7692 18196 7744
rect 19708 7692 19760 7744
rect 6378 7590 6430 7642
rect 6442 7590 6494 7642
rect 6506 7590 6558 7642
rect 6570 7590 6622 7642
rect 6634 7590 6686 7642
rect 11806 7590 11858 7642
rect 11870 7590 11922 7642
rect 11934 7590 11986 7642
rect 11998 7590 12050 7642
rect 12062 7590 12114 7642
rect 17234 7590 17286 7642
rect 17298 7590 17350 7642
rect 17362 7590 17414 7642
rect 17426 7590 17478 7642
rect 17490 7590 17542 7642
rect 22662 7590 22714 7642
rect 22726 7590 22778 7642
rect 22790 7590 22842 7642
rect 22854 7590 22906 7642
rect 22918 7590 22970 7642
rect 2872 7531 2924 7540
rect 2872 7497 2881 7531
rect 2881 7497 2915 7531
rect 2915 7497 2924 7531
rect 2872 7488 2924 7497
rect 12440 7488 12492 7540
rect 13452 7488 13504 7540
rect 17592 7531 17644 7540
rect 17592 7497 17601 7531
rect 17601 7497 17635 7531
rect 17635 7497 17644 7531
rect 17592 7488 17644 7497
rect 19248 7488 19300 7540
rect 19340 7488 19392 7540
rect 20352 7488 20404 7540
rect 4344 7463 4396 7472
rect 4344 7429 4353 7463
rect 4353 7429 4387 7463
rect 4387 7429 4396 7463
rect 4344 7420 4396 7429
rect 8944 7420 8996 7472
rect 9496 7463 9548 7472
rect 9496 7429 9505 7463
rect 9505 7429 9539 7463
rect 9539 7429 9548 7463
rect 9496 7420 9548 7429
rect 11704 7420 11756 7472
rect 15384 7420 15436 7472
rect 17868 7463 17920 7472
rect 17868 7429 17877 7463
rect 17877 7429 17911 7463
rect 17911 7429 17920 7463
rect 17868 7420 17920 7429
rect 7840 7395 7892 7404
rect 7840 7361 7849 7395
rect 7849 7361 7883 7395
rect 7883 7361 7892 7395
rect 7840 7352 7892 7361
rect 12348 7352 12400 7404
rect 12900 7395 12952 7404
rect 12900 7361 12909 7395
rect 12909 7361 12943 7395
rect 12943 7361 12952 7395
rect 12900 7352 12952 7361
rect 12992 7395 13044 7404
rect 12992 7361 13001 7395
rect 13001 7361 13035 7395
rect 13035 7361 13044 7395
rect 12992 7352 13044 7361
rect 15568 7352 15620 7404
rect 17132 7352 17184 7404
rect 15016 7284 15068 7336
rect 16948 7284 17000 7336
rect 17592 7284 17644 7336
rect 19248 7352 19300 7404
rect 20720 7420 20772 7472
rect 20536 7395 20588 7404
rect 20536 7361 20545 7395
rect 20545 7361 20579 7395
rect 20579 7361 20588 7395
rect 20536 7352 20588 7361
rect 12532 7191 12584 7200
rect 12532 7157 12541 7191
rect 12541 7157 12575 7191
rect 12575 7157 12584 7191
rect 12532 7148 12584 7157
rect 14280 7148 14332 7200
rect 15108 7148 15160 7200
rect 20352 7191 20404 7200
rect 20352 7157 20361 7191
rect 20361 7157 20395 7191
rect 20395 7157 20404 7191
rect 20352 7148 20404 7157
rect 3664 7046 3716 7098
rect 3728 7046 3780 7098
rect 3792 7046 3844 7098
rect 3856 7046 3908 7098
rect 3920 7046 3972 7098
rect 9092 7046 9144 7098
rect 9156 7046 9208 7098
rect 9220 7046 9272 7098
rect 9284 7046 9336 7098
rect 9348 7046 9400 7098
rect 14520 7046 14572 7098
rect 14584 7046 14636 7098
rect 14648 7046 14700 7098
rect 14712 7046 14764 7098
rect 14776 7046 14828 7098
rect 19948 7046 20000 7098
rect 20012 7046 20064 7098
rect 20076 7046 20128 7098
rect 20140 7046 20192 7098
rect 20204 7046 20256 7098
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 2412 6740 2464 6792
rect 3976 6740 4028 6792
rect 8944 6740 8996 6792
rect 9312 6740 9364 6792
rect 13268 6876 13320 6928
rect 13452 6876 13504 6928
rect 15752 6876 15804 6928
rect 17868 6944 17920 6996
rect 13084 6808 13136 6860
rect 13912 6808 13964 6860
rect 15200 6851 15252 6860
rect 15200 6817 15209 6851
rect 15209 6817 15243 6851
rect 15243 6817 15252 6851
rect 15200 6808 15252 6817
rect 16488 6808 16540 6860
rect 17500 6808 17552 6860
rect 17592 6851 17644 6860
rect 17592 6817 17601 6851
rect 17601 6817 17635 6851
rect 17635 6817 17644 6851
rect 17592 6808 17644 6817
rect 17684 6851 17736 6860
rect 17684 6817 17693 6851
rect 17693 6817 17727 6851
rect 17727 6817 17736 6851
rect 17684 6808 17736 6817
rect 19800 6944 19852 6996
rect 19616 6876 19668 6928
rect 20628 6808 20680 6860
rect 12624 6740 12676 6792
rect 13360 6783 13412 6792
rect 13360 6749 13369 6783
rect 13369 6749 13403 6783
rect 13403 6749 13412 6783
rect 13360 6740 13412 6749
rect 15292 6740 15344 6792
rect 17040 6740 17092 6792
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 5448 6715 5500 6724
rect 5448 6681 5466 6715
rect 5466 6681 5500 6715
rect 5448 6672 5500 6681
rect 2504 6604 2556 6656
rect 4988 6604 5040 6656
rect 8300 6647 8352 6656
rect 8300 6613 8309 6647
rect 8309 6613 8343 6647
rect 8343 6613 8352 6647
rect 8300 6604 8352 6613
rect 9772 6715 9824 6724
rect 9772 6681 9806 6715
rect 9806 6681 9824 6715
rect 9772 6672 9824 6681
rect 12716 6672 12768 6724
rect 12440 6604 12492 6656
rect 13268 6647 13320 6656
rect 13268 6613 13277 6647
rect 13277 6613 13311 6647
rect 13311 6613 13320 6647
rect 13268 6604 13320 6613
rect 16764 6715 16816 6724
rect 16764 6681 16773 6715
rect 16773 6681 16807 6715
rect 16807 6681 16816 6715
rect 16764 6672 16816 6681
rect 18604 6672 18656 6724
rect 16028 6604 16080 6656
rect 19432 6647 19484 6656
rect 19432 6613 19441 6647
rect 19441 6613 19475 6647
rect 19475 6613 19484 6647
rect 19432 6604 19484 6613
rect 6378 6502 6430 6554
rect 6442 6502 6494 6554
rect 6506 6502 6558 6554
rect 6570 6502 6622 6554
rect 6634 6502 6686 6554
rect 11806 6502 11858 6554
rect 11870 6502 11922 6554
rect 11934 6502 11986 6554
rect 11998 6502 12050 6554
rect 12062 6502 12114 6554
rect 17234 6502 17286 6554
rect 17298 6502 17350 6554
rect 17362 6502 17414 6554
rect 17426 6502 17478 6554
rect 17490 6502 17542 6554
rect 22662 6502 22714 6554
rect 22726 6502 22778 6554
rect 22790 6502 22842 6554
rect 22854 6502 22906 6554
rect 22918 6502 22970 6554
rect 3148 6443 3200 6452
rect 3148 6409 3157 6443
rect 3157 6409 3191 6443
rect 3191 6409 3200 6443
rect 3148 6400 3200 6409
rect 1676 6332 1728 6384
rect 12256 6332 12308 6384
rect 16948 6400 17000 6452
rect 15292 6332 15344 6384
rect 17132 6400 17184 6452
rect 18604 6400 18656 6452
rect 19616 6400 19668 6452
rect 2964 6264 3016 6316
rect 3148 6264 3200 6316
rect 3976 6307 4028 6316
rect 3976 6273 3985 6307
rect 3985 6273 4019 6307
rect 4019 6273 4028 6307
rect 3976 6264 4028 6273
rect 2688 6060 2740 6112
rect 6552 6239 6604 6248
rect 6552 6205 6561 6239
rect 6561 6205 6595 6239
rect 6595 6205 6604 6239
rect 6552 6196 6604 6205
rect 9312 6307 9364 6316
rect 9312 6273 9321 6307
rect 9321 6273 9355 6307
rect 9355 6273 9364 6307
rect 9312 6264 9364 6273
rect 11704 6264 11756 6316
rect 12808 6307 12860 6316
rect 12808 6273 12817 6307
rect 12817 6273 12851 6307
rect 12851 6273 12860 6307
rect 12808 6264 12860 6273
rect 13084 6307 13136 6316
rect 13084 6273 13093 6307
rect 13093 6273 13127 6307
rect 13127 6273 13136 6307
rect 13084 6264 13136 6273
rect 12532 6196 12584 6248
rect 12624 6239 12676 6248
rect 12624 6205 12633 6239
rect 12633 6205 12667 6239
rect 12667 6205 12676 6239
rect 12624 6196 12676 6205
rect 13820 6307 13872 6316
rect 13820 6273 13829 6307
rect 13829 6273 13863 6307
rect 13863 6273 13872 6307
rect 13820 6264 13872 6273
rect 14096 6307 14148 6316
rect 14096 6273 14105 6307
rect 14105 6273 14139 6307
rect 14139 6273 14148 6307
rect 14096 6264 14148 6273
rect 15108 6264 15160 6316
rect 15200 6264 15252 6316
rect 15660 6307 15712 6316
rect 15660 6273 15669 6307
rect 15669 6273 15703 6307
rect 15703 6273 15712 6307
rect 15660 6264 15712 6273
rect 15936 6264 15988 6316
rect 16764 6264 16816 6316
rect 17132 6264 17184 6316
rect 17776 6264 17828 6316
rect 18236 6307 18288 6316
rect 18236 6273 18245 6307
rect 18245 6273 18279 6307
rect 18279 6273 18288 6307
rect 18236 6264 18288 6273
rect 19340 6307 19392 6316
rect 19340 6273 19349 6307
rect 19349 6273 19383 6307
rect 19383 6273 19392 6307
rect 19340 6264 19392 6273
rect 19708 6264 19760 6316
rect 20444 6264 20496 6316
rect 14924 6196 14976 6248
rect 15752 6196 15804 6248
rect 20352 6196 20404 6248
rect 13820 6171 13872 6180
rect 13820 6137 13829 6171
rect 13829 6137 13863 6171
rect 13863 6137 13872 6171
rect 13820 6128 13872 6137
rect 17040 6171 17092 6180
rect 17040 6137 17049 6171
rect 17049 6137 17083 6171
rect 17083 6137 17092 6171
rect 17040 6128 17092 6137
rect 5632 6060 5684 6112
rect 8760 6060 8812 6112
rect 18144 6103 18196 6112
rect 18144 6069 18153 6103
rect 18153 6069 18187 6103
rect 18187 6069 18196 6103
rect 18144 6060 18196 6069
rect 3664 5958 3716 6010
rect 3728 5958 3780 6010
rect 3792 5958 3844 6010
rect 3856 5958 3908 6010
rect 3920 5958 3972 6010
rect 9092 5958 9144 6010
rect 9156 5958 9208 6010
rect 9220 5958 9272 6010
rect 9284 5958 9336 6010
rect 9348 5958 9400 6010
rect 14520 5958 14572 6010
rect 14584 5958 14636 6010
rect 14648 5958 14700 6010
rect 14712 5958 14764 6010
rect 14776 5958 14828 6010
rect 19948 5958 20000 6010
rect 20012 5958 20064 6010
rect 20076 5958 20128 6010
rect 20140 5958 20192 6010
rect 20204 5958 20256 6010
rect 2412 5856 2464 5908
rect 12808 5856 12860 5908
rect 13360 5856 13412 5908
rect 15936 5899 15988 5908
rect 15936 5865 15945 5899
rect 15945 5865 15979 5899
rect 15979 5865 15988 5899
rect 15936 5856 15988 5865
rect 17040 5856 17092 5908
rect 13452 5788 13504 5840
rect 3148 5763 3200 5772
rect 3148 5729 3157 5763
rect 3157 5729 3191 5763
rect 3191 5729 3200 5763
rect 3148 5720 3200 5729
rect 6552 5720 6604 5772
rect 7012 5720 7064 5772
rect 13268 5720 13320 5772
rect 15200 5788 15252 5840
rect 15108 5720 15160 5772
rect 9496 5652 9548 5704
rect 4436 5584 4488 5636
rect 12992 5695 13044 5704
rect 12992 5661 13001 5695
rect 13001 5661 13035 5695
rect 13035 5661 13044 5695
rect 12992 5652 13044 5661
rect 13820 5652 13872 5704
rect 14832 5695 14884 5704
rect 14832 5661 14841 5695
rect 14841 5661 14875 5695
rect 14875 5661 14884 5695
rect 14832 5652 14884 5661
rect 1768 5559 1820 5568
rect 1768 5525 1777 5559
rect 1777 5525 1811 5559
rect 1811 5525 1820 5559
rect 1768 5516 1820 5525
rect 12808 5559 12860 5568
rect 12808 5525 12817 5559
rect 12817 5525 12851 5559
rect 12851 5525 12860 5559
rect 12808 5516 12860 5525
rect 15108 5584 15160 5636
rect 15752 5627 15804 5636
rect 15752 5593 15761 5627
rect 15761 5593 15795 5627
rect 15795 5593 15804 5627
rect 15752 5584 15804 5593
rect 14280 5516 14332 5568
rect 15660 5516 15712 5568
rect 6378 5414 6430 5466
rect 6442 5414 6494 5466
rect 6506 5414 6558 5466
rect 6570 5414 6622 5466
rect 6634 5414 6686 5466
rect 11806 5414 11858 5466
rect 11870 5414 11922 5466
rect 11934 5414 11986 5466
rect 11998 5414 12050 5466
rect 12062 5414 12114 5466
rect 17234 5414 17286 5466
rect 17298 5414 17350 5466
rect 17362 5414 17414 5466
rect 17426 5414 17478 5466
rect 17490 5414 17542 5466
rect 22662 5414 22714 5466
rect 22726 5414 22778 5466
rect 22790 5414 22842 5466
rect 22854 5414 22906 5466
rect 22918 5414 22970 5466
rect 3148 5312 3200 5364
rect 13084 5312 13136 5364
rect 13728 5312 13780 5364
rect 14096 5312 14148 5364
rect 19708 5312 19760 5364
rect 4344 5287 4396 5296
rect 4344 5253 4353 5287
rect 4353 5253 4387 5287
rect 4387 5253 4396 5287
rect 4344 5244 4396 5253
rect 7840 5287 7892 5296
rect 7840 5253 7849 5287
rect 7849 5253 7883 5287
rect 7883 5253 7892 5287
rect 7840 5244 7892 5253
rect 9496 5287 9548 5296
rect 9496 5253 9505 5287
rect 9505 5253 9539 5287
rect 9539 5253 9548 5287
rect 9496 5244 9548 5253
rect 13544 5219 13596 5228
rect 13544 5185 13553 5219
rect 13553 5185 13587 5219
rect 13587 5185 13596 5219
rect 13544 5176 13596 5185
rect 15108 5244 15160 5296
rect 15660 5244 15712 5296
rect 14924 5219 14976 5228
rect 14924 5185 14933 5219
rect 14933 5185 14967 5219
rect 14967 5185 14976 5219
rect 14924 5176 14976 5185
rect 12992 5108 13044 5160
rect 17224 5219 17276 5228
rect 17224 5185 17233 5219
rect 17233 5185 17267 5219
rect 17267 5185 17276 5219
rect 17224 5176 17276 5185
rect 13820 5040 13872 5092
rect 14740 5083 14792 5092
rect 14740 5049 14768 5083
rect 14768 5049 14792 5083
rect 17132 5108 17184 5160
rect 14740 5040 14792 5049
rect 13912 4972 13964 5024
rect 3664 4870 3716 4922
rect 3728 4870 3780 4922
rect 3792 4870 3844 4922
rect 3856 4870 3908 4922
rect 3920 4870 3972 4922
rect 9092 4870 9144 4922
rect 9156 4870 9208 4922
rect 9220 4870 9272 4922
rect 9284 4870 9336 4922
rect 9348 4870 9400 4922
rect 14520 4870 14572 4922
rect 14584 4870 14636 4922
rect 14648 4870 14700 4922
rect 14712 4870 14764 4922
rect 14776 4870 14828 4922
rect 19948 4870 20000 4922
rect 20012 4870 20064 4922
rect 20076 4870 20128 4922
rect 20140 4870 20192 4922
rect 20204 4870 20256 4922
rect 8024 4768 8076 4820
rect 15660 4768 15712 4820
rect 3148 4632 3200 4684
rect 4252 4632 4304 4684
rect 9496 4632 9548 4684
rect 1676 4564 1728 4616
rect 14096 4700 14148 4752
rect 14832 4700 14884 4752
rect 7012 4607 7064 4616
rect 7012 4573 7021 4607
rect 7021 4573 7055 4607
rect 7055 4573 7064 4607
rect 7012 4564 7064 4573
rect 12716 4564 12768 4616
rect 12992 4564 13044 4616
rect 13084 4564 13136 4616
rect 13176 4607 13228 4616
rect 13176 4573 13185 4607
rect 13185 4573 13219 4607
rect 13219 4573 13228 4607
rect 14740 4632 14792 4684
rect 15016 4632 15068 4684
rect 13176 4564 13228 4573
rect 14464 4607 14516 4616
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 2504 4496 2556 4548
rect 7104 4496 7156 4548
rect 7656 4496 7708 4548
rect 12256 4496 12308 4548
rect 14924 4607 14976 4616
rect 14924 4573 14933 4607
rect 14933 4573 14967 4607
rect 14967 4573 14976 4607
rect 14924 4564 14976 4573
rect 17592 4768 17644 4820
rect 17132 4743 17184 4752
rect 17132 4709 17141 4743
rect 17141 4709 17175 4743
rect 17175 4709 17184 4743
rect 17132 4700 17184 4709
rect 15016 4496 15068 4548
rect 3240 4471 3292 4480
rect 3240 4437 3249 4471
rect 3249 4437 3283 4471
rect 3283 4437 3292 4471
rect 3240 4428 3292 4437
rect 7564 4428 7616 4480
rect 12532 4428 12584 4480
rect 12624 4471 12676 4480
rect 12624 4437 12633 4471
rect 12633 4437 12667 4471
rect 12667 4437 12676 4471
rect 12624 4428 12676 4437
rect 6378 4326 6430 4378
rect 6442 4326 6494 4378
rect 6506 4326 6558 4378
rect 6570 4326 6622 4378
rect 6634 4326 6686 4378
rect 11806 4326 11858 4378
rect 11870 4326 11922 4378
rect 11934 4326 11986 4378
rect 11998 4326 12050 4378
rect 12062 4326 12114 4378
rect 17234 4326 17286 4378
rect 17298 4326 17350 4378
rect 17362 4326 17414 4378
rect 17426 4326 17478 4378
rect 17490 4326 17542 4378
rect 22662 4326 22714 4378
rect 22726 4326 22778 4378
rect 22790 4326 22842 4378
rect 22854 4326 22906 4378
rect 22918 4326 22970 4378
rect 12256 4267 12308 4276
rect 12256 4233 12265 4267
rect 12265 4233 12299 4267
rect 12299 4233 12308 4267
rect 12256 4224 12308 4233
rect 12624 4224 12676 4276
rect 14740 4224 14792 4276
rect 7012 4156 7064 4208
rect 1676 4131 1728 4140
rect 1676 4097 1685 4131
rect 1685 4097 1719 4131
rect 1719 4097 1728 4131
rect 1676 4088 1728 4097
rect 2320 4088 2372 4140
rect 4252 4131 4304 4140
rect 4252 4097 4261 4131
rect 4261 4097 4295 4131
rect 4295 4097 4304 4131
rect 4252 4088 4304 4097
rect 4804 4088 4856 4140
rect 12164 4156 12216 4208
rect 8944 4088 8996 4140
rect 9496 4088 9548 4140
rect 12532 4088 12584 4140
rect 13268 4088 13320 4140
rect 12808 4063 12860 4072
rect 12808 4029 12817 4063
rect 12817 4029 12851 4063
rect 12851 4029 12860 4063
rect 12808 4020 12860 4029
rect 9588 3952 9640 4004
rect 2872 3884 2924 3936
rect 3148 3884 3200 3936
rect 5540 3884 5592 3936
rect 5908 3884 5960 3936
rect 8484 3927 8536 3936
rect 8484 3893 8493 3927
rect 8493 3893 8527 3927
rect 8527 3893 8536 3927
rect 8484 3884 8536 3893
rect 14464 4088 14516 4140
rect 14832 4131 14884 4140
rect 14832 4097 14841 4131
rect 14841 4097 14875 4131
rect 14875 4097 14884 4131
rect 14832 4088 14884 4097
rect 15108 4131 15160 4140
rect 15108 4097 15117 4131
rect 15117 4097 15151 4131
rect 15151 4097 15160 4131
rect 15108 4088 15160 4097
rect 15200 4131 15252 4140
rect 15200 4097 15209 4131
rect 15209 4097 15243 4131
rect 15243 4097 15252 4131
rect 15200 4088 15252 4097
rect 17132 3952 17184 4004
rect 15016 3884 15068 3936
rect 3664 3782 3716 3834
rect 3728 3782 3780 3834
rect 3792 3782 3844 3834
rect 3856 3782 3908 3834
rect 3920 3782 3972 3834
rect 9092 3782 9144 3834
rect 9156 3782 9208 3834
rect 9220 3782 9272 3834
rect 9284 3782 9336 3834
rect 9348 3782 9400 3834
rect 14520 3782 14572 3834
rect 14584 3782 14636 3834
rect 14648 3782 14700 3834
rect 14712 3782 14764 3834
rect 14776 3782 14828 3834
rect 19948 3782 20000 3834
rect 20012 3782 20064 3834
rect 20076 3782 20128 3834
rect 20140 3782 20192 3834
rect 20204 3782 20256 3834
rect 4804 3723 4856 3732
rect 4804 3689 4813 3723
rect 4813 3689 4847 3723
rect 4847 3689 4856 3723
rect 4804 3680 4856 3689
rect 5540 3680 5592 3732
rect 2872 3612 2924 3664
rect 8208 3680 8260 3732
rect 12808 3680 12860 3732
rect 14924 3680 14976 3732
rect 15200 3723 15252 3732
rect 15200 3689 15209 3723
rect 15209 3689 15243 3723
rect 15243 3689 15252 3723
rect 15200 3680 15252 3689
rect 9864 3612 9916 3664
rect 10876 3612 10928 3664
rect 11612 3655 11664 3664
rect 11612 3621 11621 3655
rect 11621 3621 11655 3655
rect 11655 3621 11664 3655
rect 11612 3612 11664 3621
rect 2780 3544 2832 3596
rect 4160 3544 4212 3596
rect 9588 3544 9640 3596
rect 1768 3476 1820 3528
rect 5080 3519 5132 3528
rect 5080 3485 5089 3519
rect 5089 3485 5123 3519
rect 5123 3485 5132 3519
rect 5080 3476 5132 3485
rect 2596 3408 2648 3460
rect 3240 3408 3292 3460
rect 5724 3408 5776 3460
rect 5908 3519 5960 3528
rect 5908 3485 5917 3519
rect 5917 3485 5951 3519
rect 5951 3485 5960 3519
rect 5908 3476 5960 3485
rect 9496 3476 9548 3528
rect 11336 3519 11388 3528
rect 11336 3485 11345 3519
rect 11345 3485 11379 3519
rect 11379 3485 11388 3519
rect 11336 3476 11388 3485
rect 13176 3544 13228 3596
rect 12716 3476 12768 3528
rect 14372 3476 14424 3528
rect 8208 3408 8260 3460
rect 10232 3408 10284 3460
rect 10968 3408 11020 3460
rect 12440 3408 12492 3460
rect 13360 3408 13412 3460
rect 10140 3340 10192 3392
rect 10876 3340 10928 3392
rect 13452 3383 13504 3392
rect 13452 3349 13461 3383
rect 13461 3349 13495 3383
rect 13495 3349 13504 3383
rect 13452 3340 13504 3349
rect 6378 3238 6430 3290
rect 6442 3238 6494 3290
rect 6506 3238 6558 3290
rect 6570 3238 6622 3290
rect 6634 3238 6686 3290
rect 11806 3238 11858 3290
rect 11870 3238 11922 3290
rect 11934 3238 11986 3290
rect 11998 3238 12050 3290
rect 12062 3238 12114 3290
rect 17234 3238 17286 3290
rect 17298 3238 17350 3290
rect 17362 3238 17414 3290
rect 17426 3238 17478 3290
rect 17490 3238 17542 3290
rect 22662 3238 22714 3290
rect 22726 3238 22778 3290
rect 22790 3238 22842 3290
rect 22854 3238 22906 3290
rect 22918 3238 22970 3290
rect 2504 3179 2556 3188
rect 2504 3145 2513 3179
rect 2513 3145 2547 3179
rect 2547 3145 2556 3179
rect 2504 3136 2556 3145
rect 7656 3179 7708 3188
rect 7656 3145 7665 3179
rect 7665 3145 7699 3179
rect 7699 3145 7708 3179
rect 7656 3136 7708 3145
rect 8024 3179 8076 3188
rect 8024 3145 8033 3179
rect 8033 3145 8067 3179
rect 8067 3145 8076 3179
rect 8024 3136 8076 3145
rect 13360 3136 13412 3188
rect 13452 3136 13504 3188
rect 15108 3136 15160 3188
rect 11612 3068 11664 3120
rect 2688 3043 2740 3052
rect 2688 3009 2697 3043
rect 2697 3009 2731 3043
rect 2731 3009 2740 3043
rect 2688 3000 2740 3009
rect 2780 3043 2832 3052
rect 2780 3009 2789 3043
rect 2789 3009 2823 3043
rect 2823 3009 2832 3043
rect 2780 3000 2832 3009
rect 3240 3000 3292 3052
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 5540 3000 5592 3052
rect 9496 3000 9548 3052
rect 10876 3000 10928 3052
rect 13176 3043 13228 3052
rect 13176 3009 13185 3043
rect 13185 3009 13219 3043
rect 13219 3009 13228 3043
rect 13176 3000 13228 3009
rect 5908 2932 5960 2984
rect 8208 2975 8260 2984
rect 8208 2941 8217 2975
rect 8217 2941 8251 2975
rect 8251 2941 8260 2975
rect 8208 2932 8260 2941
rect 8484 2932 8536 2984
rect 10140 2932 10192 2984
rect 10232 2975 10284 2984
rect 10232 2941 10241 2975
rect 10241 2941 10275 2975
rect 10275 2941 10284 2975
rect 10232 2932 10284 2941
rect 10600 2975 10652 2984
rect 10600 2941 10609 2975
rect 10609 2941 10643 2975
rect 10643 2941 10652 2975
rect 10600 2932 10652 2941
rect 2872 2864 2924 2916
rect 8944 2864 8996 2916
rect 12808 2864 12860 2916
rect 13360 3043 13412 3052
rect 13360 3009 13395 3043
rect 13395 3009 13412 3043
rect 13360 3000 13412 3009
rect 14372 3000 14424 3052
rect 14280 2932 14332 2984
rect 15016 2864 15068 2916
rect 2964 2839 3016 2848
rect 2964 2805 2973 2839
rect 2973 2805 3007 2839
rect 3007 2805 3016 2839
rect 2964 2796 3016 2805
rect 4344 2839 4396 2848
rect 4344 2805 4353 2839
rect 4353 2805 4387 2839
rect 4387 2805 4396 2839
rect 4344 2796 4396 2805
rect 5264 2839 5316 2848
rect 5264 2805 5273 2839
rect 5273 2805 5307 2839
rect 5307 2805 5316 2839
rect 5264 2796 5316 2805
rect 8852 2839 8904 2848
rect 8852 2805 8861 2839
rect 8861 2805 8895 2839
rect 8895 2805 8904 2839
rect 8852 2796 8904 2805
rect 9588 2796 9640 2848
rect 10232 2796 10284 2848
rect 12624 2796 12676 2848
rect 3664 2694 3716 2746
rect 3728 2694 3780 2746
rect 3792 2694 3844 2746
rect 3856 2694 3908 2746
rect 3920 2694 3972 2746
rect 9092 2694 9144 2746
rect 9156 2694 9208 2746
rect 9220 2694 9272 2746
rect 9284 2694 9336 2746
rect 9348 2694 9400 2746
rect 14520 2694 14572 2746
rect 14584 2694 14636 2746
rect 14648 2694 14700 2746
rect 14712 2694 14764 2746
rect 14776 2694 14828 2746
rect 19948 2694 20000 2746
rect 20012 2694 20064 2746
rect 20076 2694 20128 2746
rect 20140 2694 20192 2746
rect 20204 2694 20256 2746
rect 2320 2635 2372 2644
rect 2320 2601 2329 2635
rect 2329 2601 2363 2635
rect 2363 2601 2372 2635
rect 2320 2592 2372 2601
rect 4436 2592 4488 2644
rect 5724 2635 5776 2644
rect 5724 2601 5733 2635
rect 5733 2601 5767 2635
rect 5767 2601 5776 2635
rect 5724 2592 5776 2601
rect 7104 2592 7156 2644
rect 9496 2592 9548 2644
rect 13176 2592 13228 2644
rect 13360 2592 13412 2644
rect 2964 2524 3016 2576
rect 2596 2431 2648 2440
rect 2596 2397 2605 2431
rect 2605 2397 2639 2431
rect 2639 2397 2648 2431
rect 2596 2388 2648 2397
rect 2872 2431 2924 2440
rect 2872 2397 2881 2431
rect 2881 2397 2915 2431
rect 2915 2397 2924 2431
rect 2872 2388 2924 2397
rect 4344 2456 4396 2508
rect 5080 2456 5132 2508
rect 8208 2456 8260 2508
rect 8760 2456 8812 2508
rect 12440 2524 12492 2576
rect 5264 2388 5316 2440
rect 2688 2320 2740 2372
rect 7564 2431 7616 2440
rect 7564 2397 7573 2431
rect 7573 2397 7607 2431
rect 7607 2397 7616 2431
rect 7564 2388 7616 2397
rect 8852 2388 8904 2440
rect 10600 2456 10652 2508
rect 9588 2388 9640 2440
rect 10140 2388 10192 2440
rect 12440 2431 12492 2440
rect 12440 2397 12449 2431
rect 12449 2397 12483 2431
rect 12483 2397 12492 2431
rect 12440 2388 12492 2397
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 13084 2431 13136 2440
rect 13084 2397 13093 2431
rect 13093 2397 13127 2431
rect 13127 2397 13136 2431
rect 13084 2388 13136 2397
rect 11336 2320 11388 2372
rect 13912 2320 13964 2372
rect 14280 2252 14332 2304
rect 6378 2150 6430 2202
rect 6442 2150 6494 2202
rect 6506 2150 6558 2202
rect 6570 2150 6622 2202
rect 6634 2150 6686 2202
rect 11806 2150 11858 2202
rect 11870 2150 11922 2202
rect 11934 2150 11986 2202
rect 11998 2150 12050 2202
rect 12062 2150 12114 2202
rect 17234 2150 17286 2202
rect 17298 2150 17350 2202
rect 17362 2150 17414 2202
rect 17426 2150 17478 2202
rect 17490 2150 17542 2202
rect 22662 2150 22714 2202
rect 22726 2150 22778 2202
rect 22790 2150 22842 2202
rect 22854 2150 22906 2202
rect 22918 2150 22970 2202
<< metal2 >>
rect 6378 21788 6686 21797
rect 6378 21786 6384 21788
rect 6440 21786 6464 21788
rect 6520 21786 6544 21788
rect 6600 21786 6624 21788
rect 6680 21786 6686 21788
rect 6440 21734 6442 21786
rect 6622 21734 6624 21786
rect 6378 21732 6384 21734
rect 6440 21732 6464 21734
rect 6520 21732 6544 21734
rect 6600 21732 6624 21734
rect 6680 21732 6686 21734
rect 6378 21723 6686 21732
rect 11806 21788 12114 21797
rect 11806 21786 11812 21788
rect 11868 21786 11892 21788
rect 11948 21786 11972 21788
rect 12028 21786 12052 21788
rect 12108 21786 12114 21788
rect 11868 21734 11870 21786
rect 12050 21734 12052 21786
rect 11806 21732 11812 21734
rect 11868 21732 11892 21734
rect 11948 21732 11972 21734
rect 12028 21732 12052 21734
rect 12108 21732 12114 21734
rect 11806 21723 12114 21732
rect 17234 21788 17542 21797
rect 17234 21786 17240 21788
rect 17296 21786 17320 21788
rect 17376 21786 17400 21788
rect 17456 21786 17480 21788
rect 17536 21786 17542 21788
rect 17296 21734 17298 21786
rect 17478 21734 17480 21786
rect 17234 21732 17240 21734
rect 17296 21732 17320 21734
rect 17376 21732 17400 21734
rect 17456 21732 17480 21734
rect 17536 21732 17542 21734
rect 17234 21723 17542 21732
rect 22662 21788 22970 21797
rect 22662 21786 22668 21788
rect 22724 21786 22748 21788
rect 22804 21786 22828 21788
rect 22884 21786 22908 21788
rect 22964 21786 22970 21788
rect 22724 21734 22726 21786
rect 22906 21734 22908 21786
rect 22662 21732 22668 21734
rect 22724 21732 22748 21734
rect 22804 21732 22828 21734
rect 22884 21732 22908 21734
rect 22964 21732 22970 21734
rect 22662 21723 22970 21732
rect 3664 21244 3972 21253
rect 3664 21242 3670 21244
rect 3726 21242 3750 21244
rect 3806 21242 3830 21244
rect 3886 21242 3910 21244
rect 3966 21242 3972 21244
rect 3726 21190 3728 21242
rect 3908 21190 3910 21242
rect 3664 21188 3670 21190
rect 3726 21188 3750 21190
rect 3806 21188 3830 21190
rect 3886 21188 3910 21190
rect 3966 21188 3972 21190
rect 3664 21179 3972 21188
rect 9092 21244 9400 21253
rect 9092 21242 9098 21244
rect 9154 21242 9178 21244
rect 9234 21242 9258 21244
rect 9314 21242 9338 21244
rect 9394 21242 9400 21244
rect 9154 21190 9156 21242
rect 9336 21190 9338 21242
rect 9092 21188 9098 21190
rect 9154 21188 9178 21190
rect 9234 21188 9258 21190
rect 9314 21188 9338 21190
rect 9394 21188 9400 21190
rect 9092 21179 9400 21188
rect 14520 21244 14828 21253
rect 14520 21242 14526 21244
rect 14582 21242 14606 21244
rect 14662 21242 14686 21244
rect 14742 21242 14766 21244
rect 14822 21242 14828 21244
rect 14582 21190 14584 21242
rect 14764 21190 14766 21242
rect 14520 21188 14526 21190
rect 14582 21188 14606 21190
rect 14662 21188 14686 21190
rect 14742 21188 14766 21190
rect 14822 21188 14828 21190
rect 14520 21179 14828 21188
rect 19948 21244 20256 21253
rect 19948 21242 19954 21244
rect 20010 21242 20034 21244
rect 20090 21242 20114 21244
rect 20170 21242 20194 21244
rect 20250 21242 20256 21244
rect 20010 21190 20012 21242
rect 20192 21190 20194 21242
rect 19948 21188 19954 21190
rect 20010 21188 20034 21190
rect 20090 21188 20114 21190
rect 20170 21188 20194 21190
rect 20250 21188 20256 21190
rect 19948 21179 20256 21188
rect 6378 20700 6686 20709
rect 6378 20698 6384 20700
rect 6440 20698 6464 20700
rect 6520 20698 6544 20700
rect 6600 20698 6624 20700
rect 6680 20698 6686 20700
rect 6440 20646 6442 20698
rect 6622 20646 6624 20698
rect 6378 20644 6384 20646
rect 6440 20644 6464 20646
rect 6520 20644 6544 20646
rect 6600 20644 6624 20646
rect 6680 20644 6686 20646
rect 6378 20635 6686 20644
rect 11806 20700 12114 20709
rect 11806 20698 11812 20700
rect 11868 20698 11892 20700
rect 11948 20698 11972 20700
rect 12028 20698 12052 20700
rect 12108 20698 12114 20700
rect 11868 20646 11870 20698
rect 12050 20646 12052 20698
rect 11806 20644 11812 20646
rect 11868 20644 11892 20646
rect 11948 20644 11972 20646
rect 12028 20644 12052 20646
rect 12108 20644 12114 20646
rect 11806 20635 12114 20644
rect 17234 20700 17542 20709
rect 17234 20698 17240 20700
rect 17296 20698 17320 20700
rect 17376 20698 17400 20700
rect 17456 20698 17480 20700
rect 17536 20698 17542 20700
rect 17296 20646 17298 20698
rect 17478 20646 17480 20698
rect 17234 20644 17240 20646
rect 17296 20644 17320 20646
rect 17376 20644 17400 20646
rect 17456 20644 17480 20646
rect 17536 20644 17542 20646
rect 17234 20635 17542 20644
rect 22662 20700 22970 20709
rect 22662 20698 22668 20700
rect 22724 20698 22748 20700
rect 22804 20698 22828 20700
rect 22884 20698 22908 20700
rect 22964 20698 22970 20700
rect 22724 20646 22726 20698
rect 22906 20646 22908 20698
rect 22662 20644 22668 20646
rect 22724 20644 22748 20646
rect 22804 20644 22828 20646
rect 22884 20644 22908 20646
rect 22964 20644 22970 20646
rect 22662 20635 22970 20644
rect 3664 20156 3972 20165
rect 3664 20154 3670 20156
rect 3726 20154 3750 20156
rect 3806 20154 3830 20156
rect 3886 20154 3910 20156
rect 3966 20154 3972 20156
rect 3726 20102 3728 20154
rect 3908 20102 3910 20154
rect 3664 20100 3670 20102
rect 3726 20100 3750 20102
rect 3806 20100 3830 20102
rect 3886 20100 3910 20102
rect 3966 20100 3972 20102
rect 3664 20091 3972 20100
rect 9092 20156 9400 20165
rect 9092 20154 9098 20156
rect 9154 20154 9178 20156
rect 9234 20154 9258 20156
rect 9314 20154 9338 20156
rect 9394 20154 9400 20156
rect 9154 20102 9156 20154
rect 9336 20102 9338 20154
rect 9092 20100 9098 20102
rect 9154 20100 9178 20102
rect 9234 20100 9258 20102
rect 9314 20100 9338 20102
rect 9394 20100 9400 20102
rect 9092 20091 9400 20100
rect 14520 20156 14828 20165
rect 14520 20154 14526 20156
rect 14582 20154 14606 20156
rect 14662 20154 14686 20156
rect 14742 20154 14766 20156
rect 14822 20154 14828 20156
rect 14582 20102 14584 20154
rect 14764 20102 14766 20154
rect 14520 20100 14526 20102
rect 14582 20100 14606 20102
rect 14662 20100 14686 20102
rect 14742 20100 14766 20102
rect 14822 20100 14828 20102
rect 14520 20091 14828 20100
rect 19948 20156 20256 20165
rect 19948 20154 19954 20156
rect 20010 20154 20034 20156
rect 20090 20154 20114 20156
rect 20170 20154 20194 20156
rect 20250 20154 20256 20156
rect 20010 20102 20012 20154
rect 20192 20102 20194 20154
rect 19948 20100 19954 20102
rect 20010 20100 20034 20102
rect 20090 20100 20114 20102
rect 20170 20100 20194 20102
rect 20250 20100 20256 20102
rect 19948 20091 20256 20100
rect 940 19848 992 19854
rect 938 19816 940 19825
rect 992 19816 994 19825
rect 938 19751 994 19760
rect 1584 19780 1636 19786
rect 1584 19722 1636 19728
rect 1596 14618 1624 19722
rect 6378 19612 6686 19621
rect 6378 19610 6384 19612
rect 6440 19610 6464 19612
rect 6520 19610 6544 19612
rect 6600 19610 6624 19612
rect 6680 19610 6686 19612
rect 6440 19558 6442 19610
rect 6622 19558 6624 19610
rect 6378 19556 6384 19558
rect 6440 19556 6464 19558
rect 6520 19556 6544 19558
rect 6600 19556 6624 19558
rect 6680 19556 6686 19558
rect 6378 19547 6686 19556
rect 11806 19612 12114 19621
rect 11806 19610 11812 19612
rect 11868 19610 11892 19612
rect 11948 19610 11972 19612
rect 12028 19610 12052 19612
rect 12108 19610 12114 19612
rect 11868 19558 11870 19610
rect 12050 19558 12052 19610
rect 11806 19556 11812 19558
rect 11868 19556 11892 19558
rect 11948 19556 11972 19558
rect 12028 19556 12052 19558
rect 12108 19556 12114 19558
rect 11806 19547 12114 19556
rect 17234 19612 17542 19621
rect 17234 19610 17240 19612
rect 17296 19610 17320 19612
rect 17376 19610 17400 19612
rect 17456 19610 17480 19612
rect 17536 19610 17542 19612
rect 17296 19558 17298 19610
rect 17478 19558 17480 19610
rect 17234 19556 17240 19558
rect 17296 19556 17320 19558
rect 17376 19556 17400 19558
rect 17456 19556 17480 19558
rect 17536 19556 17542 19558
rect 17234 19547 17542 19556
rect 22662 19612 22970 19621
rect 22662 19610 22668 19612
rect 22724 19610 22748 19612
rect 22804 19610 22828 19612
rect 22884 19610 22908 19612
rect 22964 19610 22970 19612
rect 22724 19558 22726 19610
rect 22906 19558 22908 19610
rect 22662 19556 22668 19558
rect 22724 19556 22748 19558
rect 22804 19556 22828 19558
rect 22884 19556 22908 19558
rect 22964 19556 22970 19558
rect 22662 19547 22970 19556
rect 3664 19068 3972 19077
rect 3664 19066 3670 19068
rect 3726 19066 3750 19068
rect 3806 19066 3830 19068
rect 3886 19066 3910 19068
rect 3966 19066 3972 19068
rect 3726 19014 3728 19066
rect 3908 19014 3910 19066
rect 3664 19012 3670 19014
rect 3726 19012 3750 19014
rect 3806 19012 3830 19014
rect 3886 19012 3910 19014
rect 3966 19012 3972 19014
rect 3664 19003 3972 19012
rect 9092 19068 9400 19077
rect 9092 19066 9098 19068
rect 9154 19066 9178 19068
rect 9234 19066 9258 19068
rect 9314 19066 9338 19068
rect 9394 19066 9400 19068
rect 9154 19014 9156 19066
rect 9336 19014 9338 19066
rect 9092 19012 9098 19014
rect 9154 19012 9178 19014
rect 9234 19012 9258 19014
rect 9314 19012 9338 19014
rect 9394 19012 9400 19014
rect 9092 19003 9400 19012
rect 14520 19068 14828 19077
rect 14520 19066 14526 19068
rect 14582 19066 14606 19068
rect 14662 19066 14686 19068
rect 14742 19066 14766 19068
rect 14822 19066 14828 19068
rect 14582 19014 14584 19066
rect 14764 19014 14766 19066
rect 14520 19012 14526 19014
rect 14582 19012 14606 19014
rect 14662 19012 14686 19014
rect 14742 19012 14766 19014
rect 14822 19012 14828 19014
rect 14520 19003 14828 19012
rect 19948 19068 20256 19077
rect 19948 19066 19954 19068
rect 20010 19066 20034 19068
rect 20090 19066 20114 19068
rect 20170 19066 20194 19068
rect 20250 19066 20256 19068
rect 20010 19014 20012 19066
rect 20192 19014 20194 19066
rect 19948 19012 19954 19014
rect 20010 19012 20034 19014
rect 20090 19012 20114 19014
rect 20170 19012 20194 19014
rect 20250 19012 20256 19014
rect 19948 19003 20256 19012
rect 6378 18524 6686 18533
rect 6378 18522 6384 18524
rect 6440 18522 6464 18524
rect 6520 18522 6544 18524
rect 6600 18522 6624 18524
rect 6680 18522 6686 18524
rect 6440 18470 6442 18522
rect 6622 18470 6624 18522
rect 6378 18468 6384 18470
rect 6440 18468 6464 18470
rect 6520 18468 6544 18470
rect 6600 18468 6624 18470
rect 6680 18468 6686 18470
rect 6378 18459 6686 18468
rect 11806 18524 12114 18533
rect 11806 18522 11812 18524
rect 11868 18522 11892 18524
rect 11948 18522 11972 18524
rect 12028 18522 12052 18524
rect 12108 18522 12114 18524
rect 11868 18470 11870 18522
rect 12050 18470 12052 18522
rect 11806 18468 11812 18470
rect 11868 18468 11892 18470
rect 11948 18468 11972 18470
rect 12028 18468 12052 18470
rect 12108 18468 12114 18470
rect 11806 18459 12114 18468
rect 17234 18524 17542 18533
rect 17234 18522 17240 18524
rect 17296 18522 17320 18524
rect 17376 18522 17400 18524
rect 17456 18522 17480 18524
rect 17536 18522 17542 18524
rect 17296 18470 17298 18522
rect 17478 18470 17480 18522
rect 17234 18468 17240 18470
rect 17296 18468 17320 18470
rect 17376 18468 17400 18470
rect 17456 18468 17480 18470
rect 17536 18468 17542 18470
rect 17234 18459 17542 18468
rect 22662 18524 22970 18533
rect 22662 18522 22668 18524
rect 22724 18522 22748 18524
rect 22804 18522 22828 18524
rect 22884 18522 22908 18524
rect 22964 18522 22970 18524
rect 22724 18470 22726 18522
rect 22906 18470 22908 18522
rect 22662 18468 22668 18470
rect 22724 18468 22748 18470
rect 22804 18468 22828 18470
rect 22884 18468 22908 18470
rect 22964 18468 22970 18470
rect 22662 18459 22970 18468
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 3664 17980 3972 17989
rect 3664 17978 3670 17980
rect 3726 17978 3750 17980
rect 3806 17978 3830 17980
rect 3886 17978 3910 17980
rect 3966 17978 3972 17980
rect 3726 17926 3728 17978
rect 3908 17926 3910 17978
rect 3664 17924 3670 17926
rect 3726 17924 3750 17926
rect 3806 17924 3830 17926
rect 3886 17924 3910 17926
rect 3966 17924 3972 17926
rect 3664 17915 3972 17924
rect 5724 17740 5776 17746
rect 5724 17682 5776 17688
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 3240 17128 3292 17134
rect 3240 17070 3292 17076
rect 2688 16992 2740 16998
rect 2688 16934 2740 16940
rect 2596 16448 2648 16454
rect 2596 16390 2648 16396
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1768 14816 1820 14822
rect 1768 14758 1820 14764
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 938 11928 994 11937
rect 938 11863 994 11872
rect 952 11150 980 11863
rect 940 11144 992 11150
rect 940 11086 992 11092
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1688 10062 1716 10542
rect 1780 10062 1808 14758
rect 1872 14074 1900 14962
rect 1860 14068 1912 14074
rect 1860 14010 1912 14016
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1872 11286 1900 13262
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1860 11280 1912 11286
rect 1860 11222 1912 11228
rect 1964 10742 1992 12038
rect 1952 10736 2004 10742
rect 1952 10678 2004 10684
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1688 9654 1716 9998
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 1688 9042 1716 9590
rect 2056 9586 2084 15846
rect 2412 15088 2464 15094
rect 2412 15030 2464 15036
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 2148 13938 2176 14962
rect 2424 14414 2452 15030
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2320 14340 2372 14346
rect 2320 14282 2372 14288
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2240 12782 2268 13126
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2148 11626 2176 12174
rect 2240 11762 2268 12718
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 2136 11620 2188 11626
rect 2136 11562 2188 11568
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 2240 7886 2268 11698
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1688 6390 1716 6734
rect 1676 6384 1728 6390
rect 1676 6326 1728 6332
rect 2332 5930 2360 14282
rect 2424 14006 2452 14350
rect 2412 14000 2464 14006
rect 2412 13942 2464 13948
rect 2424 10266 2452 13942
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2516 11830 2544 12174
rect 2504 11824 2556 11830
rect 2504 11766 2556 11772
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2516 7886 2544 11766
rect 2608 8974 2636 16390
rect 2700 16250 2728 16934
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 3056 16108 3108 16114
rect 3056 16050 3108 16056
rect 2688 16040 2740 16046
rect 2688 15982 2740 15988
rect 2700 14414 2728 15982
rect 3068 15026 3096 16050
rect 3252 15094 3280 17070
rect 3344 16454 3372 17138
rect 3664 16892 3972 16901
rect 3664 16890 3670 16892
rect 3726 16890 3750 16892
rect 3806 16890 3830 16892
rect 3886 16890 3910 16892
rect 3966 16890 3972 16892
rect 3726 16838 3728 16890
rect 3908 16838 3910 16890
rect 3664 16836 3670 16838
rect 3726 16836 3750 16838
rect 3806 16836 3830 16838
rect 3886 16836 3910 16838
rect 3966 16836 3972 16838
rect 3664 16827 3972 16836
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3240 15088 3292 15094
rect 3240 15030 3292 15036
rect 3344 15026 3372 16390
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 3664 15804 3972 15813
rect 3664 15802 3670 15804
rect 3726 15802 3750 15804
rect 3806 15802 3830 15804
rect 3886 15802 3910 15804
rect 3966 15802 3972 15804
rect 3726 15750 3728 15802
rect 3908 15750 3910 15802
rect 3664 15748 3670 15750
rect 3726 15748 3750 15750
rect 3806 15748 3830 15750
rect 3886 15748 3910 15750
rect 3966 15748 3972 15750
rect 3664 15739 3972 15748
rect 4436 15360 4488 15366
rect 4436 15302 4488 15308
rect 3056 15020 3108 15026
rect 3056 14962 3108 14968
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2700 13870 2728 14350
rect 3068 14346 3096 14962
rect 3344 14346 3372 14962
rect 3424 14816 3476 14822
rect 3424 14758 3476 14764
rect 3056 14340 3108 14346
rect 3056 14282 3108 14288
rect 3332 14340 3384 14346
rect 3332 14282 3384 14288
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 2700 12850 2728 13330
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 2884 12374 2912 12854
rect 2872 12368 2924 12374
rect 2872 12310 2924 12316
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2792 11762 2820 12242
rect 2884 12102 2912 12310
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2792 10810 2820 11698
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2424 6798 2452 7686
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 2516 6662 2544 7822
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2700 6118 2728 7754
rect 2884 7546 2912 9590
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2976 6322 3004 13126
rect 3068 9450 3096 14282
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3160 12442 3188 13262
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 3148 12164 3200 12170
rect 3252 12152 3280 12582
rect 3200 12124 3280 12152
rect 3148 12106 3200 12112
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 3160 6458 3188 12106
rect 3344 9178 3372 14282
rect 3436 13938 3464 14758
rect 3664 14716 3972 14725
rect 3664 14714 3670 14716
rect 3726 14714 3750 14716
rect 3806 14714 3830 14716
rect 3886 14714 3910 14716
rect 3966 14714 3972 14716
rect 3726 14662 3728 14714
rect 3908 14662 3910 14714
rect 3664 14660 3670 14662
rect 3726 14660 3750 14662
rect 3806 14660 3830 14662
rect 3886 14660 3910 14662
rect 3966 14660 3972 14662
rect 3664 14651 3972 14660
rect 4080 14618 4108 14962
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 3516 14544 3568 14550
rect 3516 14486 3568 14492
rect 3528 13938 3556 14486
rect 4344 14476 4396 14482
rect 4344 14418 4396 14424
rect 4356 14006 4384 14418
rect 4344 14000 4396 14006
rect 4344 13942 4396 13948
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3664 13628 3972 13637
rect 3664 13626 3670 13628
rect 3726 13626 3750 13628
rect 3806 13626 3830 13628
rect 3886 13626 3910 13628
rect 3966 13626 3972 13628
rect 3726 13574 3728 13626
rect 3908 13574 3910 13626
rect 3664 13572 3670 13574
rect 3726 13572 3750 13574
rect 3806 13572 3830 13574
rect 3886 13572 3910 13574
rect 3966 13572 3972 13574
rect 3664 13563 3972 13572
rect 3608 13320 3660 13326
rect 3608 13262 3660 13268
rect 3620 12986 3648 13262
rect 3608 12980 3660 12986
rect 3608 12922 3660 12928
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 3424 12912 3476 12918
rect 3424 12854 3476 12860
rect 3436 12238 3464 12854
rect 3664 12540 3972 12549
rect 3664 12538 3670 12540
rect 3726 12538 3750 12540
rect 3806 12538 3830 12540
rect 3886 12538 3910 12540
rect 3966 12538 3972 12540
rect 3726 12486 3728 12538
rect 3908 12486 3910 12538
rect 3664 12484 3670 12486
rect 3726 12484 3750 12486
rect 3806 12484 3830 12486
rect 3886 12484 3910 12486
rect 3966 12484 3972 12486
rect 3664 12475 3972 12484
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 4172 11762 4200 12922
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 4264 11778 4292 12038
rect 4160 11756 4212 11762
rect 4264 11750 4384 11778
rect 4160 11698 4212 11704
rect 4356 11694 4384 11750
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 3664 11452 3972 11461
rect 3664 11450 3670 11452
rect 3726 11450 3750 11452
rect 3806 11450 3830 11452
rect 3886 11450 3910 11452
rect 3966 11450 3972 11452
rect 3726 11398 3728 11450
rect 3908 11398 3910 11450
rect 3664 11396 3670 11398
rect 3726 11396 3750 11398
rect 3806 11396 3830 11398
rect 3886 11396 3910 11398
rect 3966 11396 3972 11398
rect 3664 11387 3972 11396
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 3664 10364 3972 10373
rect 3664 10362 3670 10364
rect 3726 10362 3750 10364
rect 3806 10362 3830 10364
rect 3886 10362 3910 10364
rect 3966 10362 3972 10364
rect 3726 10310 3728 10362
rect 3908 10310 3910 10362
rect 3664 10308 3670 10310
rect 3726 10308 3750 10310
rect 3806 10308 3830 10310
rect 3886 10308 3910 10310
rect 3966 10308 3972 10310
rect 3664 10299 3972 10308
rect 4172 10130 4200 11086
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 4172 9586 4200 10066
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 3664 9276 3972 9285
rect 3664 9274 3670 9276
rect 3726 9274 3750 9276
rect 3806 9274 3830 9276
rect 3886 9274 3910 9276
rect 3966 9274 3972 9276
rect 3726 9222 3728 9274
rect 3908 9222 3910 9274
rect 3664 9220 3670 9222
rect 3726 9220 3750 9222
rect 3806 9220 3830 9222
rect 3886 9220 3910 9222
rect 3966 9220 3972 9222
rect 3664 9211 3972 9220
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 4356 8634 4384 11630
rect 4448 10062 4476 15302
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4540 9586 4568 15846
rect 4724 15570 4752 17478
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4816 16250 4844 16934
rect 4908 16658 4936 17478
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 4908 15026 4936 16594
rect 5092 16590 5120 17138
rect 5736 17134 5764 17682
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 6378 17436 6686 17445
rect 6378 17434 6384 17436
rect 6440 17434 6464 17436
rect 6520 17434 6544 17436
rect 6600 17434 6624 17436
rect 6680 17434 6686 17436
rect 6440 17382 6442 17434
rect 6622 17382 6624 17434
rect 6378 17380 6384 17382
rect 6440 17380 6464 17382
rect 6520 17380 6544 17382
rect 6600 17380 6624 17382
rect 6680 17380 6686 17382
rect 6378 17371 6686 17380
rect 7024 17270 7052 17614
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7012 17264 7064 17270
rect 7012 17206 7064 17212
rect 5724 17128 5776 17134
rect 5724 17070 5776 17076
rect 5736 16658 5764 17070
rect 5724 16652 5776 16658
rect 5724 16594 5776 16600
rect 6736 16652 6788 16658
rect 6736 16594 6788 16600
rect 5080 16584 5132 16590
rect 5080 16526 5132 16532
rect 5632 16584 5684 16590
rect 5632 16526 5684 16532
rect 5092 15366 5120 16526
rect 5172 16516 5224 16522
rect 5172 16458 5224 16464
rect 5184 16046 5212 16458
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 5184 15570 5212 15982
rect 5172 15564 5224 15570
rect 5172 15506 5224 15512
rect 5080 15360 5132 15366
rect 5080 15302 5132 15308
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 4896 15020 4948 15026
rect 4896 14962 4948 14968
rect 4816 13734 4844 14962
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4816 13258 4844 13670
rect 4804 13252 4856 13258
rect 4804 13194 4856 13200
rect 4816 12850 4844 13194
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4632 11762 4660 12582
rect 4724 12306 4752 12786
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4816 8566 4844 11494
rect 4908 10810 4936 14962
rect 4988 14000 5040 14006
rect 4988 13942 5040 13948
rect 5000 13870 5028 13942
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4804 8560 4856 8566
rect 4804 8502 4856 8508
rect 3664 8188 3972 8197
rect 3664 8186 3670 8188
rect 3726 8186 3750 8188
rect 3806 8186 3830 8188
rect 3886 8186 3910 8188
rect 3966 8186 3972 8188
rect 3726 8134 3728 8186
rect 3908 8134 3910 8186
rect 3664 8132 3670 8134
rect 3726 8132 3750 8134
rect 3806 8132 3830 8134
rect 3886 8132 3910 8134
rect 3966 8132 3972 8134
rect 3664 8123 3972 8132
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4356 7478 4384 7686
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 3664 7100 3972 7109
rect 3664 7098 3670 7100
rect 3726 7098 3750 7100
rect 3806 7098 3830 7100
rect 3886 7098 3910 7100
rect 3966 7098 3972 7100
rect 3726 7046 3728 7098
rect 3908 7046 3910 7098
rect 3664 7044 3670 7046
rect 3726 7044 3750 7046
rect 3806 7044 3830 7046
rect 3886 7044 3910 7046
rect 3966 7044 3972 7046
rect 3664 7035 3972 7044
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3988 6322 4016 6734
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2332 5914 2452 5930
rect 2332 5908 2464 5914
rect 2332 5902 2412 5908
rect 2412 5850 2464 5856
rect 3160 5778 3188 6258
rect 3664 6012 3972 6021
rect 3664 6010 3670 6012
rect 3726 6010 3750 6012
rect 3806 6010 3830 6012
rect 3886 6010 3910 6012
rect 3966 6010 3972 6012
rect 3726 5958 3728 6010
rect 3908 5958 3910 6010
rect 3664 5956 3670 5958
rect 3726 5956 3750 5958
rect 3806 5956 3830 5958
rect 3886 5956 3910 5958
rect 3966 5956 3972 5958
rect 3664 5947 3972 5956
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 1768 5568 1820 5574
rect 1768 5510 1820 5516
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1688 4146 1716 4558
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1780 3534 1808 5510
rect 3160 5370 3188 5714
rect 3148 5364 3200 5370
rect 3148 5306 3200 5312
rect 3160 4690 3188 5306
rect 4356 5302 4384 7414
rect 5000 6662 5028 13806
rect 5092 10266 5120 15302
rect 5184 14618 5212 15506
rect 5276 15026 5304 16050
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5552 15094 5580 15302
rect 5540 15088 5592 15094
rect 5540 15030 5592 15036
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 5184 14278 5212 14554
rect 5276 14414 5304 14962
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 5276 9450 5304 14350
rect 5368 13870 5396 14350
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5368 11150 5396 12038
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 5264 9444 5316 9450
rect 5264 9386 5316 9392
rect 5460 6730 5488 13874
rect 5552 10742 5580 14758
rect 5644 14278 5672 16526
rect 6378 16348 6686 16357
rect 6378 16346 6384 16348
rect 6440 16346 6464 16348
rect 6520 16346 6544 16348
rect 6600 16346 6624 16348
rect 6680 16346 6686 16348
rect 6440 16294 6442 16346
rect 6622 16294 6624 16346
rect 6378 16292 6384 16294
rect 6440 16292 6464 16294
rect 6520 16292 6544 16294
rect 6600 16292 6624 16294
rect 6680 16292 6686 16294
rect 6378 16283 6686 16292
rect 6748 16232 6776 16594
rect 6920 16244 6972 16250
rect 6748 16204 6920 16232
rect 6748 15586 6776 16204
rect 6920 16186 6972 16192
rect 6748 15558 6960 15586
rect 6932 15502 6960 15558
rect 6920 15496 6972 15502
rect 6920 15438 6972 15444
rect 6378 15260 6686 15269
rect 6378 15258 6384 15260
rect 6440 15258 6464 15260
rect 6520 15258 6544 15260
rect 6600 15258 6624 15260
rect 6680 15258 6686 15260
rect 6440 15206 6442 15258
rect 6622 15206 6624 15258
rect 6378 15204 6384 15206
rect 6440 15204 6464 15206
rect 6520 15204 6544 15206
rect 6600 15204 6624 15206
rect 6680 15204 6686 15206
rect 6378 15195 6686 15204
rect 6932 15042 6960 15438
rect 6932 15014 7052 15042
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6656 14482 6684 14758
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 5816 14340 5868 14346
rect 5816 14282 5868 14288
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5724 12912 5776 12918
rect 5724 12854 5776 12860
rect 5736 12646 5764 12854
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5644 12238 5672 12582
rect 5736 12306 5764 12582
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 4436 5636 4488 5642
rect 4436 5578 4488 5584
rect 4344 5296 4396 5302
rect 4344 5238 4396 5244
rect 3664 4924 3972 4933
rect 3664 4922 3670 4924
rect 3726 4922 3750 4924
rect 3806 4922 3830 4924
rect 3886 4922 3910 4924
rect 3966 4922 3972 4924
rect 3726 4870 3728 4922
rect 3908 4870 3910 4922
rect 3664 4868 3670 4870
rect 3726 4868 3750 4870
rect 3806 4868 3830 4870
rect 3886 4868 3910 4870
rect 3966 4868 3972 4870
rect 3664 4859 3972 4868
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 2504 4548 2556 4554
rect 2504 4490 2556 4496
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 2332 2650 2360 4082
rect 2516 3194 2544 4490
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3146 4040 3202 4049
rect 3146 3975 3202 3984
rect 3160 3942 3188 3975
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 2884 3670 2912 3878
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 2596 3460 2648 3466
rect 2596 3402 2648 3408
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 2608 2446 2636 3402
rect 2792 3058 2820 3538
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 2700 2378 2728 2994
rect 2884 2922 2912 3606
rect 3252 3466 3280 4422
rect 4264 4146 4292 4626
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 3664 3836 3972 3845
rect 3664 3834 3670 3836
rect 3726 3834 3750 3836
rect 3806 3834 3830 3836
rect 3886 3834 3910 3836
rect 3966 3834 3972 3836
rect 3726 3782 3728 3834
rect 3908 3782 3910 3834
rect 3664 3780 3670 3782
rect 3726 3780 3750 3782
rect 3806 3780 3830 3782
rect 3886 3780 3910 3782
rect 3966 3780 3972 3782
rect 3664 3771 3972 3780
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 3240 3460 3292 3466
rect 3240 3402 3292 3408
rect 3252 3058 3280 3402
rect 4172 3058 4200 3538
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 2872 2916 2924 2922
rect 2872 2858 2924 2864
rect 2884 2446 2912 2858
rect 2964 2848 3016 2854
rect 2964 2790 3016 2796
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 2976 2582 3004 2790
rect 3664 2748 3972 2757
rect 3664 2746 3670 2748
rect 3726 2746 3750 2748
rect 3806 2746 3830 2748
rect 3886 2746 3910 2748
rect 3966 2746 3972 2748
rect 3726 2694 3728 2746
rect 3908 2694 3910 2746
rect 3664 2692 3670 2694
rect 3726 2692 3750 2694
rect 3806 2692 3830 2694
rect 3886 2692 3910 2694
rect 3966 2692 3972 2694
rect 3664 2683 3972 2692
rect 2964 2576 3016 2582
rect 2964 2518 3016 2524
rect 4356 2514 4384 2790
rect 4448 2650 4476 5578
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4816 3738 4844 4082
rect 5552 3942 5580 7754
rect 5828 6914 5856 14282
rect 6378 14172 6686 14181
rect 6378 14170 6384 14172
rect 6440 14170 6464 14172
rect 6520 14170 6544 14172
rect 6600 14170 6624 14172
rect 6680 14170 6686 14172
rect 6440 14118 6442 14170
rect 6622 14118 6624 14170
rect 6378 14116 6384 14118
rect 6440 14116 6464 14118
rect 6520 14116 6544 14118
rect 6600 14116 6624 14118
rect 6680 14116 6686 14118
rect 6378 14107 6686 14116
rect 6828 14000 6880 14006
rect 6932 13988 6960 15014
rect 7024 14958 7052 15014
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 6880 13960 6960 13988
rect 6828 13942 6880 13948
rect 7116 13938 7144 17478
rect 7208 17202 7236 17614
rect 8116 17332 8168 17338
rect 8116 17274 8168 17280
rect 8128 17202 8156 17274
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 8116 17196 8168 17202
rect 8116 17138 8168 17144
rect 7208 16726 7236 17138
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7196 16720 7248 16726
rect 7196 16662 7248 16668
rect 7484 16590 7512 16730
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 7196 16516 7248 16522
rect 7196 16458 7248 16464
rect 7208 16250 7236 16458
rect 7300 16436 7328 16526
rect 7300 16408 7420 16436
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7208 15502 7236 15846
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 7392 14346 7420 16408
rect 7484 16250 7512 16526
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 8128 16046 8156 16526
rect 8116 16040 8168 16046
rect 8116 15982 8168 15988
rect 8128 15162 8156 15982
rect 8220 15162 8248 17614
rect 8312 17066 8340 17614
rect 8404 17202 8432 18158
rect 8864 17678 8892 18226
rect 8944 18080 8996 18086
rect 8944 18022 8996 18028
rect 8956 17814 8984 18022
rect 9092 17980 9400 17989
rect 9092 17978 9098 17980
rect 9154 17978 9178 17980
rect 9234 17978 9258 17980
rect 9314 17978 9338 17980
rect 9394 17978 9400 17980
rect 9154 17926 9156 17978
rect 9336 17926 9338 17978
rect 9092 17924 9098 17926
rect 9154 17924 9178 17926
rect 9234 17924 9258 17926
rect 9314 17924 9338 17926
rect 9394 17924 9400 17926
rect 9092 17915 9400 17924
rect 14520 17980 14828 17989
rect 14520 17978 14526 17980
rect 14582 17978 14606 17980
rect 14662 17978 14686 17980
rect 14742 17978 14766 17980
rect 14822 17978 14828 17980
rect 14582 17926 14584 17978
rect 14764 17926 14766 17978
rect 14520 17924 14526 17926
rect 14582 17924 14606 17926
rect 14662 17924 14686 17926
rect 14742 17924 14766 17926
rect 14822 17924 14828 17926
rect 14520 17915 14828 17924
rect 19948 17980 20256 17989
rect 19948 17978 19954 17980
rect 20010 17978 20034 17980
rect 20090 17978 20114 17980
rect 20170 17978 20194 17980
rect 20250 17978 20256 17980
rect 20010 17926 20012 17978
rect 20192 17926 20194 17978
rect 19948 17924 19954 17926
rect 20010 17924 20034 17926
rect 20090 17924 20114 17926
rect 20170 17924 20194 17926
rect 20250 17924 20256 17926
rect 19948 17915 20256 17924
rect 8944 17808 8996 17814
rect 8944 17750 8996 17756
rect 9312 17808 9364 17814
rect 9312 17750 9364 17756
rect 8852 17672 8904 17678
rect 8852 17614 8904 17620
rect 8864 17338 8892 17614
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8956 17202 8984 17750
rect 9324 17678 9352 17750
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 10876 17740 10928 17746
rect 10876 17682 10928 17688
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 9416 17338 9444 17682
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 10600 17672 10652 17678
rect 10652 17620 10732 17626
rect 10600 17614 10732 17620
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 8312 16794 8340 17002
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8404 16522 8432 17138
rect 9092 16892 9400 16901
rect 9092 16890 9098 16892
rect 9154 16890 9178 16892
rect 9234 16890 9258 16892
rect 9314 16890 9338 16892
rect 9394 16890 9400 16892
rect 9154 16838 9156 16890
rect 9336 16838 9338 16890
rect 9092 16836 9098 16838
rect 9154 16836 9178 16838
rect 9234 16836 9258 16838
rect 9314 16836 9338 16838
rect 9394 16836 9400 16838
rect 9092 16827 9400 16836
rect 9508 16590 9536 17478
rect 9968 17202 9996 17614
rect 10612 17598 10732 17614
rect 10600 17536 10652 17542
rect 10600 17478 10652 17484
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9692 16658 9720 17138
rect 9968 16726 9996 17138
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10520 16794 10548 16934
rect 10508 16788 10560 16794
rect 10508 16730 10560 16736
rect 9956 16720 10008 16726
rect 9956 16662 10008 16668
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 8392 16516 8444 16522
rect 8392 16458 8444 16464
rect 8404 16046 8432 16458
rect 9508 16114 9536 16526
rect 9692 16114 9720 16594
rect 10612 16590 10640 17478
rect 10704 17202 10732 17598
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10416 16516 10468 16522
rect 10416 16458 10468 16464
rect 10140 16176 10192 16182
rect 10140 16118 10192 16124
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 9092 15804 9400 15813
rect 9092 15802 9098 15804
rect 9154 15802 9178 15804
rect 9234 15802 9258 15804
rect 9314 15802 9338 15804
rect 9394 15802 9400 15804
rect 9154 15750 9156 15802
rect 9336 15750 9338 15802
rect 9092 15748 9098 15750
rect 9154 15748 9178 15750
rect 9234 15748 9258 15750
rect 9314 15748 9338 15750
rect 9394 15748 9400 15750
rect 9092 15739 9400 15748
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8128 14890 8156 15098
rect 8116 14884 8168 14890
rect 8116 14826 8168 14832
rect 7380 14340 7432 14346
rect 7380 14282 7432 14288
rect 8024 14340 8076 14346
rect 8024 14282 8076 14288
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 6378 13084 6686 13093
rect 6378 13082 6384 13084
rect 6440 13082 6464 13084
rect 6520 13082 6544 13084
rect 6600 13082 6624 13084
rect 6680 13082 6686 13084
rect 6440 13030 6442 13082
rect 6622 13030 6624 13082
rect 6378 13028 6384 13030
rect 6440 13028 6464 13030
rect 6520 13028 6544 13030
rect 6600 13028 6624 13030
rect 6680 13028 6686 13030
rect 6378 13019 6686 13028
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7024 12442 7052 12786
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 7116 12170 7144 12786
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6288 11354 6316 12038
rect 6378 11996 6686 12005
rect 6378 11994 6384 11996
rect 6440 11994 6464 11996
rect 6520 11994 6544 11996
rect 6600 11994 6624 11996
rect 6680 11994 6686 11996
rect 6440 11942 6442 11994
rect 6622 11942 6624 11994
rect 6378 11940 6384 11942
rect 6440 11940 6464 11942
rect 6520 11940 6544 11942
rect 6600 11940 6624 11942
rect 6680 11940 6686 11942
rect 6378 11931 6686 11940
rect 7116 11354 7144 12106
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 7208 11150 7236 12582
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 6378 10908 6686 10917
rect 6378 10906 6384 10908
rect 6440 10906 6464 10908
rect 6520 10906 6544 10908
rect 6600 10906 6624 10908
rect 6680 10906 6686 10908
rect 6440 10854 6442 10906
rect 6622 10854 6624 10906
rect 6378 10852 6384 10854
rect 6440 10852 6464 10854
rect 6520 10852 6544 10854
rect 6600 10852 6624 10854
rect 6680 10852 6686 10854
rect 6378 10843 6686 10852
rect 6932 10674 6960 11086
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 6748 10130 6776 10542
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 6378 9820 6686 9829
rect 6378 9818 6384 9820
rect 6440 9818 6464 9820
rect 6520 9818 6544 9820
rect 6600 9818 6624 9820
rect 6680 9818 6686 9820
rect 6440 9766 6442 9818
rect 6622 9766 6624 9818
rect 6378 9764 6384 9766
rect 6440 9764 6464 9766
rect 6520 9764 6544 9766
rect 6600 9764 6624 9766
rect 6680 9764 6686 9766
rect 6378 9755 6686 9764
rect 6378 8732 6686 8741
rect 6378 8730 6384 8732
rect 6440 8730 6464 8732
rect 6520 8730 6544 8732
rect 6600 8730 6624 8732
rect 6680 8730 6686 8732
rect 6440 8678 6442 8730
rect 6622 8678 6624 8730
rect 6378 8676 6384 8678
rect 6440 8676 6464 8678
rect 6520 8676 6544 8678
rect 6600 8676 6624 8678
rect 6680 8676 6686 8678
rect 6378 8667 6686 8676
rect 6748 8498 6776 10066
rect 7300 8566 7328 14214
rect 7932 12912 7984 12918
rect 7932 12854 7984 12860
rect 7748 12708 7800 12714
rect 7748 12650 7800 12656
rect 7760 12442 7788 12650
rect 7944 12646 7972 12854
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 7944 12238 7972 12582
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 8036 8634 8064 14282
rect 8220 14006 8248 15098
rect 9232 15026 9260 15302
rect 10152 15026 10180 16118
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10336 15502 10364 15982
rect 10428 15706 10456 16458
rect 10704 16182 10732 17138
rect 10888 17134 10916 17682
rect 11806 17436 12114 17445
rect 11806 17434 11812 17436
rect 11868 17434 11892 17436
rect 11948 17434 11972 17436
rect 12028 17434 12052 17436
rect 12108 17434 12114 17436
rect 11868 17382 11870 17434
rect 12050 17382 12052 17434
rect 11806 17380 11812 17382
rect 11868 17380 11892 17382
rect 11948 17380 11972 17382
rect 12028 17380 12052 17382
rect 12108 17380 12114 17382
rect 11806 17371 12114 17380
rect 17234 17436 17542 17445
rect 17234 17434 17240 17436
rect 17296 17434 17320 17436
rect 17376 17434 17400 17436
rect 17456 17434 17480 17436
rect 17536 17434 17542 17436
rect 17296 17382 17298 17434
rect 17478 17382 17480 17434
rect 17234 17380 17240 17382
rect 17296 17380 17320 17382
rect 17376 17380 17400 17382
rect 17456 17380 17480 17382
rect 17536 17380 17542 17382
rect 17234 17371 17542 17380
rect 22662 17436 22970 17445
rect 22662 17434 22668 17436
rect 22724 17434 22748 17436
rect 22804 17434 22828 17436
rect 22884 17434 22908 17436
rect 22964 17434 22970 17436
rect 22724 17382 22726 17434
rect 22906 17382 22908 17434
rect 22662 17380 22668 17382
rect 22724 17380 22748 17382
rect 22804 17380 22828 17382
rect 22884 17380 22908 17382
rect 22964 17380 22970 17382
rect 22662 17371 22970 17380
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10692 16176 10744 16182
rect 10692 16118 10744 16124
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 8312 14482 8340 14962
rect 8852 14952 8904 14958
rect 8852 14894 8904 14900
rect 8864 14550 8892 14894
rect 8852 14544 8904 14550
rect 8852 14486 8904 14492
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 8128 9994 8156 13806
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 8220 10742 8248 12582
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 7840 7812 7892 7818
rect 7840 7754 7892 7760
rect 6378 7644 6686 7653
rect 6378 7642 6384 7644
rect 6440 7642 6464 7644
rect 6520 7642 6544 7644
rect 6600 7642 6624 7644
rect 6680 7642 6686 7644
rect 6440 7590 6442 7642
rect 6622 7590 6624 7642
rect 6378 7588 6384 7590
rect 6440 7588 6464 7590
rect 6520 7588 6544 7590
rect 6600 7588 6624 7590
rect 6680 7588 6686 7590
rect 6378 7579 6686 7588
rect 7852 7410 7880 7754
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 5644 6886 5856 6914
rect 5644 6118 5672 6886
rect 6378 6556 6686 6565
rect 6378 6554 6384 6556
rect 6440 6554 6464 6556
rect 6520 6554 6544 6556
rect 6600 6554 6624 6556
rect 6680 6554 6686 6556
rect 6440 6502 6442 6554
rect 6622 6502 6624 6554
rect 6378 6500 6384 6502
rect 6440 6500 6464 6502
rect 6520 6500 6544 6502
rect 6600 6500 6624 6502
rect 6680 6500 6686 6502
rect 6378 6491 6686 6500
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5644 3754 5672 6054
rect 6564 5778 6592 6190
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 6378 5468 6686 5477
rect 6378 5466 6384 5468
rect 6440 5466 6464 5468
rect 6520 5466 6544 5468
rect 6600 5466 6624 5468
rect 6680 5466 6686 5468
rect 6440 5414 6442 5466
rect 6622 5414 6624 5466
rect 6378 5412 6384 5414
rect 6440 5412 6464 5414
rect 6520 5412 6544 5414
rect 6600 5412 6624 5414
rect 6680 5412 6686 5414
rect 6378 5403 6686 5412
rect 7024 4622 7052 5714
rect 7852 5302 7880 7346
rect 8312 6662 8340 14418
rect 8956 14414 8984 14962
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9092 14716 9400 14725
rect 9092 14714 9098 14716
rect 9154 14714 9178 14716
rect 9234 14714 9258 14716
rect 9314 14714 9338 14716
rect 9394 14714 9400 14716
rect 9154 14662 9156 14714
rect 9336 14662 9338 14714
rect 9092 14660 9098 14662
rect 9154 14660 9178 14662
rect 9234 14660 9258 14662
rect 9314 14660 9338 14662
rect 9394 14660 9400 14662
rect 9092 14651 9400 14660
rect 9508 14618 9536 14894
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 10336 14482 10364 15438
rect 10888 15434 10916 17070
rect 14520 16892 14828 16901
rect 14520 16890 14526 16892
rect 14582 16890 14606 16892
rect 14662 16890 14686 16892
rect 14742 16890 14766 16892
rect 14822 16890 14828 16892
rect 14582 16838 14584 16890
rect 14764 16838 14766 16890
rect 14520 16836 14526 16838
rect 14582 16836 14606 16838
rect 14662 16836 14686 16838
rect 14742 16836 14766 16838
rect 14822 16836 14828 16838
rect 14520 16827 14828 16836
rect 19948 16892 20256 16901
rect 19948 16890 19954 16892
rect 20010 16890 20034 16892
rect 20090 16890 20114 16892
rect 20170 16890 20194 16892
rect 20250 16890 20256 16892
rect 20010 16838 20012 16890
rect 20192 16838 20194 16890
rect 19948 16836 19954 16838
rect 20010 16836 20034 16838
rect 20090 16836 20114 16838
rect 20170 16836 20194 16838
rect 20250 16836 20256 16838
rect 19948 16827 20256 16836
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 10980 15638 11008 16526
rect 11806 16348 12114 16357
rect 11806 16346 11812 16348
rect 11868 16346 11892 16348
rect 11948 16346 11972 16348
rect 12028 16346 12052 16348
rect 12108 16346 12114 16348
rect 11868 16294 11870 16346
rect 12050 16294 12052 16346
rect 11806 16292 11812 16294
rect 11868 16292 11892 16294
rect 11948 16292 11972 16294
rect 12028 16292 12052 16294
rect 12108 16292 12114 16294
rect 11806 16283 12114 16292
rect 17234 16348 17542 16357
rect 17234 16346 17240 16348
rect 17296 16346 17320 16348
rect 17376 16346 17400 16348
rect 17456 16346 17480 16348
rect 17536 16346 17542 16348
rect 17296 16294 17298 16346
rect 17478 16294 17480 16346
rect 17234 16292 17240 16294
rect 17296 16292 17320 16294
rect 17376 16292 17400 16294
rect 17456 16292 17480 16294
rect 17536 16292 17542 16294
rect 17234 16283 17542 16292
rect 22662 16348 22970 16357
rect 22662 16346 22668 16348
rect 22724 16346 22748 16348
rect 22804 16346 22828 16348
rect 22884 16346 22908 16348
rect 22964 16346 22970 16348
rect 22724 16294 22726 16346
rect 22906 16294 22908 16346
rect 22662 16292 22668 16294
rect 22724 16292 22748 16294
rect 22804 16292 22828 16294
rect 22884 16292 22908 16294
rect 22964 16292 22970 16294
rect 22662 16283 22970 16292
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 10968 15632 11020 15638
rect 10968 15574 11020 15580
rect 10876 15428 10928 15434
rect 10876 15370 10928 15376
rect 10888 15026 10916 15370
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 9508 13938 9536 14350
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8404 12850 8432 13126
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8496 10266 8524 12038
rect 8680 10810 8708 12718
rect 8772 12102 8800 13874
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 8956 13326 8984 13806
rect 9092 13628 9400 13637
rect 9092 13626 9098 13628
rect 9154 13626 9178 13628
rect 9234 13626 9258 13628
rect 9314 13626 9338 13628
rect 9394 13626 9400 13628
rect 9154 13574 9156 13626
rect 9336 13574 9338 13626
rect 9092 13572 9098 13574
rect 9154 13572 9178 13574
rect 9234 13572 9258 13574
rect 9314 13572 9338 13574
rect 9394 13572 9400 13574
rect 9092 13563 9400 13572
rect 9508 13394 9536 13874
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 8956 12986 8984 13262
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8956 12306 8984 12582
rect 9092 12540 9400 12549
rect 9092 12538 9098 12540
rect 9154 12538 9178 12540
rect 9234 12538 9258 12540
rect 9314 12538 9338 12540
rect 9394 12538 9400 12540
rect 9154 12486 9156 12538
rect 9336 12486 9338 12538
rect 9092 12484 9098 12486
rect 9154 12484 9178 12486
rect 9234 12484 9258 12486
rect 9314 12484 9338 12486
rect 9394 12484 9400 12486
rect 9092 12475 9400 12484
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 9600 12238 9628 12718
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 9092 11452 9400 11461
rect 9092 11450 9098 11452
rect 9154 11450 9178 11452
rect 9234 11450 9258 11452
rect 9314 11450 9338 11452
rect 9394 11450 9400 11452
rect 9154 11398 9156 11450
rect 9336 11398 9338 11450
rect 9092 11396 9098 11398
rect 9154 11396 9178 11398
rect 9234 11396 9258 11398
rect 9314 11396 9338 11398
rect 9394 11396 9400 11398
rect 9092 11387 9400 11396
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9092 10364 9400 10373
rect 9092 10362 9098 10364
rect 9154 10362 9178 10364
rect 9234 10362 9258 10364
rect 9314 10362 9338 10364
rect 9394 10362 9400 10364
rect 9154 10310 9156 10362
rect 9336 10310 9338 10362
rect 9092 10308 9098 10310
rect 9154 10308 9178 10310
rect 9234 10308 9258 10310
rect 9314 10308 9338 10310
rect 9394 10308 9400 10310
rect 9092 10299 9400 10308
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 9508 10062 9536 10542
rect 9692 10266 9720 14418
rect 10508 14340 10560 14346
rect 10508 14282 10560 14288
rect 10784 14340 10836 14346
rect 10784 14282 10836 14288
rect 10520 13734 10548 14282
rect 10796 13938 10824 14282
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10888 13818 10916 14962
rect 10980 14958 11008 15574
rect 11072 15502 11100 16050
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 11072 15026 11100 15438
rect 11806 15260 12114 15269
rect 11806 15258 11812 15260
rect 11868 15258 11892 15260
rect 11948 15258 11972 15260
rect 12028 15258 12052 15260
rect 12108 15258 12114 15260
rect 11868 15206 11870 15258
rect 12050 15206 12052 15258
rect 11806 15204 11812 15206
rect 11868 15204 11892 15206
rect 11948 15204 11972 15206
rect 12028 15204 12052 15206
rect 12108 15204 12114 15206
rect 11806 15195 12114 15204
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 10968 14952 11020 14958
rect 10968 14894 11020 14900
rect 10796 13790 10916 13818
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10520 13326 10548 13670
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9784 10742 9812 13126
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10336 12850 10364 12922
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 9864 12368 9916 12374
rect 9864 12310 9916 12316
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9508 9586 9536 9998
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9092 9276 9400 9285
rect 9092 9274 9098 9276
rect 9154 9274 9178 9276
rect 9234 9274 9258 9276
rect 9314 9274 9338 9276
rect 9394 9274 9400 9276
rect 9154 9222 9156 9274
rect 9336 9222 9338 9274
rect 9092 9220 9098 9222
rect 9154 9220 9178 9222
rect 9234 9220 9258 9222
rect 9314 9220 9338 9222
rect 9394 9220 9400 9222
rect 9092 9211 9400 9220
rect 9508 9042 9536 9522
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9508 8498 9536 8978
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9092 8188 9400 8197
rect 9092 8186 9098 8188
rect 9154 8186 9178 8188
rect 9234 8186 9258 8188
rect 9314 8186 9338 8188
rect 9394 8186 9400 8188
rect 9154 8134 9156 8186
rect 9336 8134 9338 8186
rect 9092 8132 9098 8134
rect 9154 8132 9178 8134
rect 9234 8132 9258 8134
rect 9314 8132 9338 8134
rect 9394 8132 9400 8134
rect 9092 8123 9400 8132
rect 9508 7954 9536 8434
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9508 7478 9536 7890
rect 8944 7472 8996 7478
rect 8944 7414 8996 7420
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 8956 6798 8984 7414
rect 9092 7100 9400 7109
rect 9092 7098 9098 7100
rect 9154 7098 9178 7100
rect 9234 7098 9258 7100
rect 9314 7098 9338 7100
rect 9394 7098 9400 7100
rect 9154 7046 9156 7098
rect 9336 7046 9338 7098
rect 9092 7044 9098 7046
rect 9154 7044 9178 7046
rect 9234 7044 9258 7046
rect 9314 7044 9338 7046
rect 9394 7044 9400 7046
rect 9092 7035 9400 7044
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 9324 6322 9352 6734
rect 9784 6730 9812 9658
rect 9876 9654 9904 12310
rect 10336 12306 10364 12786
rect 10324 12300 10376 12306
rect 10324 12242 10376 12248
rect 10428 12170 10456 12786
rect 10704 12442 10732 13262
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10416 12164 10468 12170
rect 10416 12106 10468 12112
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 10796 8634 10824 13790
rect 10968 13252 11020 13258
rect 10968 13194 11020 13200
rect 10980 12850 11008 13194
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 10888 12238 10916 12786
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10888 10810 10916 12174
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10966 10160 11022 10169
rect 10966 10095 11022 10104
rect 10980 10062 11008 10095
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 11072 9178 11100 14962
rect 11520 14408 11572 14414
rect 11520 14350 11572 14356
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11164 12306 11192 12786
rect 11532 12374 11560 14350
rect 11806 14172 12114 14181
rect 11806 14170 11812 14172
rect 11868 14170 11892 14172
rect 11948 14170 11972 14172
rect 12028 14170 12052 14172
rect 12108 14170 12114 14172
rect 11868 14118 11870 14170
rect 12050 14118 12052 14170
rect 11806 14116 11812 14118
rect 11868 14116 11892 14118
rect 11948 14116 11972 14118
rect 12028 14116 12052 14118
rect 12108 14116 12114 14118
rect 11806 14107 12114 14116
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 11624 12986 11652 13262
rect 11806 13084 12114 13093
rect 11806 13082 11812 13084
rect 11868 13082 11892 13084
rect 11948 13082 11972 13084
rect 12028 13082 12052 13084
rect 12108 13082 12114 13084
rect 11868 13030 11870 13082
rect 12050 13030 12052 13082
rect 11806 13028 11812 13030
rect 11868 13028 11892 13030
rect 11948 13028 11972 13030
rect 12028 13028 12052 13030
rect 12108 13028 12114 13030
rect 11806 13019 12114 13028
rect 12452 12986 12480 13262
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 11624 12102 11652 12786
rect 12360 12102 12388 12786
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 11256 8498 11284 10406
rect 11716 9450 11744 12038
rect 11806 11996 12114 12005
rect 11806 11994 11812 11996
rect 11868 11994 11892 11996
rect 11948 11994 11972 11996
rect 12028 11994 12052 11996
rect 12108 11994 12114 11996
rect 11868 11942 11870 11994
rect 12050 11942 12052 11994
rect 11806 11940 11812 11942
rect 11868 11940 11892 11942
rect 11948 11940 11972 11942
rect 12028 11940 12052 11942
rect 12108 11940 12114 11942
rect 11806 11931 12114 11940
rect 11806 10908 12114 10917
rect 11806 10906 11812 10908
rect 11868 10906 11892 10908
rect 11948 10906 11972 10908
rect 12028 10906 12052 10908
rect 12108 10906 12114 10908
rect 11868 10854 11870 10906
rect 12050 10854 12052 10906
rect 11806 10852 11812 10854
rect 11868 10852 11892 10854
rect 11948 10852 11972 10854
rect 12028 10852 12052 10854
rect 12108 10852 12114 10854
rect 11806 10843 12114 10852
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 11806 9820 12114 9829
rect 11806 9818 11812 9820
rect 11868 9818 11892 9820
rect 11948 9818 11972 9820
rect 12028 9818 12052 9820
rect 12108 9818 12114 9820
rect 11868 9766 11870 9818
rect 12050 9766 12052 9818
rect 11806 9764 11812 9766
rect 11868 9764 11892 9766
rect 11948 9764 11972 9766
rect 12028 9764 12052 9766
rect 12108 9764 12114 9766
rect 11806 9755 12114 9764
rect 12176 9722 12204 10610
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12360 9994 12388 10542
rect 12348 9988 12400 9994
rect 12348 9930 12400 9936
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 11704 9444 11756 9450
rect 11704 9386 11756 9392
rect 11806 8732 12114 8741
rect 11806 8730 11812 8732
rect 11868 8730 11892 8732
rect 11948 8730 11972 8732
rect 12028 8730 12052 8732
rect 12108 8730 12114 8732
rect 11868 8678 11870 8730
rect 12050 8678 12052 8730
rect 11806 8676 11812 8678
rect 11868 8676 11892 8678
rect 11948 8676 11972 8678
rect 12028 8676 12052 8678
rect 12108 8676 12114 8678
rect 11806 8667 12114 8676
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 11806 7644 12114 7653
rect 11806 7642 11812 7644
rect 11868 7642 11892 7644
rect 11948 7642 11972 7644
rect 12028 7642 12052 7644
rect 12108 7642 12114 7644
rect 11868 7590 11870 7642
rect 12050 7590 12052 7642
rect 11806 7588 11812 7590
rect 11868 7588 11892 7590
rect 11948 7588 11972 7590
rect 12028 7588 12052 7590
rect 12108 7588 12114 7590
rect 11806 7579 12114 7588
rect 11704 7472 11756 7478
rect 11704 7414 11756 7420
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 11716 6322 11744 7414
rect 11806 6556 12114 6565
rect 11806 6554 11812 6556
rect 11868 6554 11892 6556
rect 11948 6554 11972 6556
rect 12028 6554 12052 6556
rect 12108 6554 12114 6556
rect 11868 6502 11870 6554
rect 12050 6502 12052 6554
rect 11806 6500 11812 6502
rect 11868 6500 11892 6502
rect 11948 6500 11972 6502
rect 12028 6500 12052 6502
rect 12108 6500 12114 6502
rect 11806 6491 12114 6500
rect 9312 6316 9364 6322
rect 11704 6316 11756 6322
rect 9364 6276 9536 6304
rect 9312 6258 9364 6264
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 6378 4380 6686 4389
rect 6378 4378 6384 4380
rect 6440 4378 6464 4380
rect 6520 4378 6544 4380
rect 6600 4378 6624 4380
rect 6680 4378 6686 4380
rect 6440 4326 6442 4378
rect 6622 4326 6624 4378
rect 6378 4324 6384 4326
rect 6440 4324 6464 4326
rect 6520 4324 6544 4326
rect 6600 4324 6624 4326
rect 6680 4324 6686 4326
rect 6378 4315 6686 4324
rect 7024 4214 7052 4558
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7656 4548 7708 4554
rect 7656 4490 7708 4496
rect 7012 4208 7064 4214
rect 7012 4150 7064 4156
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5552 3738 5672 3754
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 5540 3732 5672 3738
rect 5592 3726 5672 3732
rect 5540 3674 5592 3680
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 5092 2514 5120 3470
rect 5552 3058 5580 3674
rect 5920 3534 5948 3878
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 4344 2508 4396 2514
rect 4344 2450 4396 2456
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 5276 2446 5304 2790
rect 5736 2650 5764 3402
rect 5920 2990 5948 3470
rect 6378 3292 6686 3301
rect 6378 3290 6384 3292
rect 6440 3290 6464 3292
rect 6520 3290 6544 3292
rect 6600 3290 6624 3292
rect 6680 3290 6686 3292
rect 6440 3238 6442 3290
rect 6622 3238 6624 3290
rect 6378 3236 6384 3238
rect 6440 3236 6464 3238
rect 6520 3236 6544 3238
rect 6600 3236 6624 3238
rect 6680 3236 6686 3238
rect 6378 3227 6686 3236
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 7116 2650 7144 4490
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7576 2446 7604 4422
rect 7668 3194 7696 4490
rect 8036 3194 8064 4762
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8220 3466 8248 3674
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8220 2990 8248 3402
rect 8496 2990 8524 3878
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8220 2514 8248 2926
rect 8772 2514 8800 6054
rect 9092 6012 9400 6021
rect 9092 6010 9098 6012
rect 9154 6010 9178 6012
rect 9234 6010 9258 6012
rect 9314 6010 9338 6012
rect 9394 6010 9400 6012
rect 9154 5958 9156 6010
rect 9336 5958 9338 6010
rect 9092 5956 9098 5958
rect 9154 5956 9178 5958
rect 9234 5956 9258 5958
rect 9314 5956 9338 5958
rect 9394 5956 9400 5958
rect 9092 5947 9400 5956
rect 9508 5710 9536 6276
rect 11704 6258 11756 6264
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9508 5302 9536 5646
rect 11806 5468 12114 5477
rect 11806 5466 11812 5468
rect 11868 5466 11892 5468
rect 11948 5466 11972 5468
rect 12028 5466 12052 5468
rect 12108 5466 12114 5468
rect 11868 5414 11870 5466
rect 12050 5414 12052 5466
rect 11806 5412 11812 5414
rect 11868 5412 11892 5414
rect 11948 5412 11972 5414
rect 12028 5412 12052 5414
rect 12108 5412 12114 5414
rect 11806 5403 12114 5412
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 9092 4924 9400 4933
rect 9092 4922 9098 4924
rect 9154 4922 9178 4924
rect 9234 4922 9258 4924
rect 9314 4922 9338 4924
rect 9394 4922 9400 4924
rect 9154 4870 9156 4922
rect 9336 4870 9338 4922
rect 9092 4868 9098 4870
rect 9154 4868 9178 4870
rect 9234 4868 9258 4870
rect 9314 4868 9338 4870
rect 9394 4868 9400 4870
rect 9092 4859 9400 4868
rect 9508 4690 9536 5238
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9508 4146 9536 4626
rect 11806 4380 12114 4389
rect 11806 4378 11812 4380
rect 11868 4378 11892 4380
rect 11948 4378 11972 4380
rect 12028 4378 12052 4380
rect 12108 4378 12114 4380
rect 11868 4326 11870 4378
rect 12050 4326 12052 4378
rect 11806 4324 11812 4326
rect 11868 4324 11892 4326
rect 11948 4324 11972 4326
rect 12028 4324 12052 4326
rect 12108 4324 12114 4326
rect 11806 4315 12114 4324
rect 12176 4214 12204 7822
rect 12268 6390 12296 8434
rect 12360 7818 12388 9930
rect 12636 8022 12664 12786
rect 13096 12442 13124 13874
rect 13280 13530 13308 13874
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13464 13326 13492 13874
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 13188 11098 13216 12378
rect 13280 12084 13308 13194
rect 13464 13002 13492 13262
rect 13372 12974 13492 13002
rect 13372 12238 13400 12974
rect 13556 12442 13584 13806
rect 13648 12442 13676 13806
rect 14384 13530 14412 16186
rect 14520 15804 14828 15813
rect 14520 15802 14526 15804
rect 14582 15802 14606 15804
rect 14662 15802 14686 15804
rect 14742 15802 14766 15804
rect 14822 15802 14828 15804
rect 14582 15750 14584 15802
rect 14764 15750 14766 15802
rect 14520 15748 14526 15750
rect 14582 15748 14606 15750
rect 14662 15748 14686 15750
rect 14742 15748 14766 15750
rect 14822 15748 14828 15750
rect 14520 15739 14828 15748
rect 19948 15804 20256 15813
rect 19948 15802 19954 15804
rect 20010 15802 20034 15804
rect 20090 15802 20114 15804
rect 20170 15802 20194 15804
rect 20250 15802 20256 15804
rect 20010 15750 20012 15802
rect 20192 15750 20194 15802
rect 19948 15748 19954 15750
rect 20010 15748 20034 15750
rect 20090 15748 20114 15750
rect 20170 15748 20194 15750
rect 20250 15748 20256 15750
rect 19948 15739 20256 15748
rect 17234 15260 17542 15269
rect 17234 15258 17240 15260
rect 17296 15258 17320 15260
rect 17376 15258 17400 15260
rect 17456 15258 17480 15260
rect 17536 15258 17542 15260
rect 17296 15206 17298 15258
rect 17478 15206 17480 15258
rect 17234 15204 17240 15206
rect 17296 15204 17320 15206
rect 17376 15204 17400 15206
rect 17456 15204 17480 15206
rect 17536 15204 17542 15206
rect 17234 15195 17542 15204
rect 22662 15260 22970 15269
rect 22662 15258 22668 15260
rect 22724 15258 22748 15260
rect 22804 15258 22828 15260
rect 22884 15258 22908 15260
rect 22964 15258 22970 15260
rect 22724 15206 22726 15258
rect 22906 15206 22908 15258
rect 22662 15204 22668 15206
rect 22724 15204 22748 15206
rect 22804 15204 22828 15206
rect 22884 15204 22908 15206
rect 22964 15204 22970 15206
rect 22662 15195 22970 15204
rect 14520 14716 14828 14725
rect 14520 14714 14526 14716
rect 14582 14714 14606 14716
rect 14662 14714 14686 14716
rect 14742 14714 14766 14716
rect 14822 14714 14828 14716
rect 14582 14662 14584 14714
rect 14764 14662 14766 14714
rect 14520 14660 14526 14662
rect 14582 14660 14606 14662
rect 14662 14660 14686 14662
rect 14742 14660 14766 14662
rect 14822 14660 14828 14662
rect 14520 14651 14828 14660
rect 19948 14716 20256 14725
rect 19948 14714 19954 14716
rect 20010 14714 20034 14716
rect 20090 14714 20114 14716
rect 20170 14714 20194 14716
rect 20250 14714 20256 14716
rect 20010 14662 20012 14714
rect 20192 14662 20194 14714
rect 19948 14660 19954 14662
rect 20010 14660 20034 14662
rect 20090 14660 20114 14662
rect 20170 14660 20194 14662
rect 20250 14660 20256 14662
rect 19948 14651 20256 14660
rect 17234 14172 17542 14181
rect 17234 14170 17240 14172
rect 17296 14170 17320 14172
rect 17376 14170 17400 14172
rect 17456 14170 17480 14172
rect 17536 14170 17542 14172
rect 17296 14118 17298 14170
rect 17478 14118 17480 14170
rect 17234 14116 17240 14118
rect 17296 14116 17320 14118
rect 17376 14116 17400 14118
rect 17456 14116 17480 14118
rect 17536 14116 17542 14118
rect 17234 14107 17542 14116
rect 22662 14172 22970 14181
rect 22662 14170 22668 14172
rect 22724 14170 22748 14172
rect 22804 14170 22828 14172
rect 22884 14170 22908 14172
rect 22964 14170 22970 14172
rect 22724 14118 22726 14170
rect 22906 14118 22908 14170
rect 22662 14116 22668 14118
rect 22724 14116 22748 14118
rect 22804 14116 22828 14118
rect 22884 14116 22908 14118
rect 22964 14116 22970 14118
rect 22662 14107 22970 14116
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 14520 13628 14828 13637
rect 14520 13626 14526 13628
rect 14582 13626 14606 13628
rect 14662 13626 14686 13628
rect 14742 13626 14766 13628
rect 14822 13626 14828 13628
rect 14582 13574 14584 13626
rect 14764 13574 14766 13626
rect 14520 13572 14526 13574
rect 14582 13572 14606 13574
rect 14662 13572 14686 13574
rect 14742 13572 14766 13574
rect 14822 13572 14828 13574
rect 14520 13563 14828 13572
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13740 12646 13768 13262
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13464 12084 13492 12174
rect 13280 12056 13492 12084
rect 13004 11070 13216 11098
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12912 10266 12940 10542
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12348 7812 12400 7818
rect 12348 7754 12400 7760
rect 12360 7410 12388 7754
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12452 6662 12480 7482
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12256 6384 12308 6390
rect 12256 6326 12308 6332
rect 12544 6254 12572 7142
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12636 6254 12664 6734
rect 12728 6730 12756 9862
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12820 8634 12848 8978
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12820 7818 12848 8570
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12912 7410 12940 7686
rect 13004 7562 13032 11070
rect 13176 11008 13228 11014
rect 13176 10950 13228 10956
rect 13188 10742 13216 10950
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 13096 10062 13124 10474
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 13096 9178 13124 9862
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 13280 8906 13308 10406
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13280 7886 13308 8842
rect 13372 8634 13400 8910
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13464 8090 13492 12056
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13556 8906 13584 12038
rect 13648 10266 13676 12378
rect 13740 12306 13768 12582
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13740 10810 13768 11086
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13544 8900 13596 8906
rect 13544 8842 13596 8848
rect 13556 8430 13584 8842
rect 13740 8498 13768 10746
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13360 8016 13412 8022
rect 13556 7970 13584 8366
rect 13360 7958 13412 7964
rect 13372 7886 13400 7958
rect 13464 7942 13584 7970
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13004 7534 13124 7562
rect 12990 7440 13046 7449
rect 12900 7404 12952 7410
rect 12990 7375 12992 7384
rect 12900 7346 12952 7352
rect 13044 7375 13046 7384
rect 12992 7346 13044 7352
rect 13096 6866 13124 7534
rect 13280 6934 13308 7822
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 13372 6882 13400 7822
rect 13464 7750 13492 7942
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13464 7546 13492 7686
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13452 6928 13504 6934
rect 13372 6876 13452 6882
rect 13372 6870 13504 6876
rect 13084 6860 13136 6866
rect 13372 6854 13492 6870
rect 13084 6802 13136 6808
rect 13096 6746 13124 6802
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 13004 6718 13124 6746
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12820 5914 12848 6258
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 13004 5710 13032 6718
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12256 4548 12308 4554
rect 12256 4490 12308 4496
rect 12268 4282 12296 4490
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12624 4480 12676 4486
rect 12624 4422 12676 4428
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 12164 4208 12216 4214
rect 12164 4150 12216 4156
rect 12544 4146 12572 4422
rect 12636 4282 12664 4422
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 8956 2922 8984 4082
rect 9092 3836 9400 3845
rect 9092 3834 9098 3836
rect 9154 3834 9178 3836
rect 9234 3834 9258 3836
rect 9314 3834 9338 3836
rect 9394 3834 9400 3836
rect 9154 3782 9156 3834
rect 9336 3782 9338 3834
rect 9092 3780 9098 3782
rect 9154 3780 9178 3782
rect 9234 3780 9258 3782
rect 9314 3780 9338 3782
rect 9394 3780 9400 3782
rect 9092 3771 9400 3780
rect 9508 3534 9536 4082
rect 9588 4004 9640 4010
rect 9588 3946 9640 3952
rect 9600 3602 9628 3946
rect 9864 3664 9916 3670
rect 10876 3664 10928 3670
rect 9916 3612 10876 3618
rect 9864 3606 10928 3612
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 9588 3596 9640 3602
rect 9876 3590 10916 3606
rect 9588 3538 9640 3544
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 8944 2916 8996 2922
rect 8944 2858 8996 2864
rect 8852 2848 8904 2854
rect 8852 2790 8904 2796
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 8864 2446 8892 2790
rect 9092 2748 9400 2757
rect 9092 2746 9098 2748
rect 9154 2746 9178 2748
rect 9234 2746 9258 2748
rect 9314 2746 9338 2748
rect 9394 2746 9400 2748
rect 9154 2694 9156 2746
rect 9336 2694 9338 2746
rect 9092 2692 9098 2694
rect 9154 2692 9178 2694
rect 9234 2692 9258 2694
rect 9314 2692 9338 2694
rect 9394 2692 9400 2694
rect 9092 2683 9400 2692
rect 9508 2650 9536 2994
rect 9600 2854 9628 3538
rect 11336 3528 11388 3534
rect 10966 3496 11022 3505
rect 10232 3460 10284 3466
rect 11336 3470 11388 3476
rect 10966 3431 10968 3440
rect 10232 3402 10284 3408
rect 11020 3431 11022 3440
rect 10968 3402 11020 3408
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10152 2990 10180 3334
rect 10244 2990 10272 3402
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10888 3058 10916 3334
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 10600 2984 10652 2990
rect 10600 2926 10652 2932
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9600 2446 9628 2790
rect 10152 2446 10180 2926
rect 10244 2854 10272 2926
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 10612 2514 10640 2926
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 8852 2440 8904 2446
rect 8852 2382 8904 2388
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 11348 2378 11376 3470
rect 11624 3126 11652 3606
rect 12728 3534 12756 4558
rect 12820 4078 12848 5510
rect 13004 5166 13032 5646
rect 13096 5370 13124 6258
rect 13280 5778 13308 6598
rect 13372 5914 13400 6734
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13464 5846 13492 6854
rect 13832 6322 13860 13330
rect 13924 12238 13952 13330
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 14016 12434 14044 13262
rect 14016 12406 14136 12434
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 14004 11076 14056 11082
rect 14004 11018 14056 11024
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13924 10674 13952 10950
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 14016 10606 14044 11018
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 13912 8424 13964 8430
rect 13910 8392 13912 8401
rect 13964 8392 13966 8401
rect 13910 8327 13966 8336
rect 13924 6866 13952 8327
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 14108 6322 14136 12406
rect 14188 11280 14240 11286
rect 14188 11222 14240 11228
rect 14278 11248 14334 11257
rect 14200 11082 14228 11222
rect 14278 11183 14280 11192
rect 14332 11183 14334 11192
rect 14280 11154 14332 11160
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 14200 10538 14228 11018
rect 14188 10532 14240 10538
rect 14188 10474 14240 10480
rect 14200 9722 14228 10474
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 14200 8430 14228 9658
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13452 5840 13504 5846
rect 13452 5782 13504 5788
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 13832 5710 13860 6122
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 12992 5160 13044 5166
rect 13096 5137 13124 5306
rect 13740 5250 13768 5306
rect 13556 5234 13768 5250
rect 13544 5228 13768 5234
rect 13596 5222 13768 5228
rect 13544 5170 13596 5176
rect 12992 5102 13044 5108
rect 13082 5128 13138 5137
rect 13832 5098 13860 5646
rect 14108 5370 14136 6258
rect 14292 5574 14320 7142
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 13082 5063 13138 5072
rect 13820 5092 13872 5098
rect 13096 4706 13124 5063
rect 13820 5034 13872 5040
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 13004 4678 13124 4706
rect 13004 4622 13032 4678
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12820 3738 12848 4014
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12716 3528 12768 3534
rect 12636 3476 12716 3482
rect 12636 3470 12768 3476
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12636 3454 12756 3470
rect 11806 3292 12114 3301
rect 11806 3290 11812 3292
rect 11868 3290 11892 3292
rect 11948 3290 11972 3292
rect 12028 3290 12052 3292
rect 12108 3290 12114 3292
rect 11868 3238 11870 3290
rect 12050 3238 12052 3290
rect 11806 3236 11812 3238
rect 11868 3236 11892 3238
rect 11948 3236 11972 3238
rect 12028 3236 12052 3238
rect 12108 3236 12114 3238
rect 11806 3227 12114 3236
rect 11612 3120 11664 3126
rect 11612 3062 11664 3068
rect 12452 2582 12480 3402
rect 12636 2854 12664 3454
rect 12820 2922 12848 3674
rect 12808 2916 12860 2922
rect 12808 2858 12860 2864
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 12452 2446 12480 2518
rect 12636 2446 12664 2790
rect 13096 2446 13124 4558
rect 13188 3602 13216 4558
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13176 3596 13228 3602
rect 13176 3538 13228 3544
rect 13280 3074 13308 4082
rect 13360 3460 13412 3466
rect 13360 3402 13412 3408
rect 13372 3194 13400 3402
rect 13452 3392 13504 3398
rect 13452 3334 13504 3340
rect 13464 3194 13492 3334
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13280 3058 13400 3074
rect 13176 3052 13228 3058
rect 13280 3052 13412 3058
rect 13280 3046 13360 3052
rect 13176 2994 13228 3000
rect 13360 2994 13412 3000
rect 13188 2650 13216 2994
rect 13372 2650 13400 2994
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13924 2378 13952 4966
rect 14108 4758 14136 5306
rect 14096 4752 14148 4758
rect 14096 4694 14148 4700
rect 14384 3534 14412 13466
rect 15212 13258 15240 13806
rect 16764 13796 16816 13802
rect 16764 13738 16816 13744
rect 15844 13456 15896 13462
rect 15844 13398 15896 13404
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 15856 13190 15884 13398
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 16040 12986 16068 13262
rect 16500 13190 16528 13262
rect 16488 13184 16540 13190
rect 16488 13126 16540 13132
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 15120 12628 15148 12786
rect 15396 12782 15424 12922
rect 16776 12918 16804 13738
rect 19948 13628 20256 13637
rect 19948 13626 19954 13628
rect 20010 13626 20034 13628
rect 20090 13626 20114 13628
rect 20170 13626 20194 13628
rect 20250 13626 20256 13628
rect 20010 13574 20012 13626
rect 20192 13574 20194 13626
rect 19948 13572 19954 13574
rect 20010 13572 20034 13574
rect 20090 13572 20114 13574
rect 20170 13572 20194 13574
rect 20250 13572 20256 13574
rect 19948 13563 20256 13572
rect 19800 13524 19852 13530
rect 19800 13466 19852 13472
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 17776 13456 17828 13462
rect 17776 13398 17828 13404
rect 18236 13456 18288 13462
rect 18236 13398 18288 13404
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 16856 13184 16908 13190
rect 16856 13126 16908 13132
rect 16764 12912 16816 12918
rect 16764 12854 16816 12860
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15488 12628 15516 12786
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15120 12600 15516 12628
rect 14520 12540 14828 12549
rect 14520 12538 14526 12540
rect 14582 12538 14606 12540
rect 14662 12538 14686 12540
rect 14742 12538 14766 12540
rect 14822 12538 14828 12540
rect 14582 12486 14584 12538
rect 14764 12486 14766 12538
rect 14520 12484 14526 12486
rect 14582 12484 14606 12486
rect 14662 12484 14686 12486
rect 14742 12484 14766 12486
rect 14822 12484 14828 12486
rect 14520 12475 14828 12484
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 14936 11558 14964 12174
rect 15396 11898 15424 12174
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 14924 11552 14976 11558
rect 14924 11494 14976 11500
rect 14520 11452 14828 11461
rect 14520 11450 14526 11452
rect 14582 11450 14606 11452
rect 14662 11450 14686 11452
rect 14742 11450 14766 11452
rect 14822 11450 14828 11452
rect 14582 11398 14584 11450
rect 14764 11398 14766 11450
rect 14520 11396 14526 11398
rect 14582 11396 14606 11398
rect 14662 11396 14686 11398
rect 14742 11396 14766 11398
rect 14822 11396 14828 11398
rect 14520 11387 14828 11396
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14568 11150 14596 11290
rect 14936 11150 14964 11494
rect 15396 11354 15424 11834
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15488 11234 15516 12600
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15212 11206 15516 11234
rect 15660 11212 15712 11218
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14924 11144 14976 11150
rect 14924 11086 14976 11092
rect 14476 10810 14504 11086
rect 14464 10804 14516 10810
rect 14464 10746 14516 10752
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 14520 10364 14828 10373
rect 14520 10362 14526 10364
rect 14582 10362 14606 10364
rect 14662 10362 14686 10364
rect 14742 10362 14766 10364
rect 14822 10362 14828 10364
rect 14582 10310 14584 10362
rect 14764 10310 14766 10362
rect 14520 10308 14526 10310
rect 14582 10308 14606 10310
rect 14662 10308 14686 10310
rect 14742 10308 14766 10310
rect 14822 10308 14828 10310
rect 14520 10299 14828 10308
rect 15028 9722 15056 10542
rect 15120 9994 15148 10542
rect 15108 9988 15160 9994
rect 15108 9930 15160 9936
rect 15016 9716 15068 9722
rect 15016 9658 15068 9664
rect 14520 9276 14828 9285
rect 14520 9274 14526 9276
rect 14582 9274 14606 9276
rect 14662 9274 14686 9276
rect 14742 9274 14766 9276
rect 14822 9274 14828 9276
rect 14582 9222 14584 9274
rect 14764 9222 14766 9274
rect 14520 9220 14526 9222
rect 14582 9220 14606 9222
rect 14662 9220 14686 9222
rect 14742 9220 14766 9222
rect 14822 9220 14828 9222
rect 14520 9211 14828 9220
rect 15120 9178 15148 9930
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14936 8294 14964 8910
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14520 8188 14828 8197
rect 14520 8186 14526 8188
rect 14582 8186 14606 8188
rect 14662 8186 14686 8188
rect 14742 8186 14766 8188
rect 14822 8186 14828 8188
rect 14582 8134 14584 8186
rect 14764 8134 14766 8186
rect 14520 8132 14526 8134
rect 14582 8132 14606 8134
rect 14662 8132 14686 8134
rect 14742 8132 14766 8134
rect 14822 8132 14828 8134
rect 14520 8123 14828 8132
rect 14936 7954 14964 8230
rect 14924 7948 14976 7954
rect 14924 7890 14976 7896
rect 15028 7342 15056 8774
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 15120 8090 15148 8366
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15108 7744 15160 7750
rect 15108 7686 15160 7692
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 15120 7206 15148 7686
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 14520 7100 14828 7109
rect 14520 7098 14526 7100
rect 14582 7098 14606 7100
rect 14662 7098 14686 7100
rect 14742 7098 14766 7100
rect 14822 7098 14828 7100
rect 14582 7046 14584 7098
rect 14764 7046 14766 7098
rect 14520 7044 14526 7046
rect 14582 7044 14606 7046
rect 14662 7044 14686 7046
rect 14742 7044 14766 7046
rect 14822 7044 14828 7046
rect 14520 7035 14828 7044
rect 15212 6866 15240 11206
rect 15660 11154 15712 11160
rect 15476 11144 15528 11150
rect 15290 11112 15346 11121
rect 15476 11086 15528 11092
rect 15290 11047 15292 11056
rect 15344 11047 15346 11056
rect 15292 11018 15344 11024
rect 15488 10810 15516 11086
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15672 10266 15700 11154
rect 15764 11150 15792 12038
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15292 8628 15344 8634
rect 15344 8588 15608 8616
rect 15292 8570 15344 8576
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15212 6322 15240 6802
rect 15304 6798 15332 7890
rect 15396 7478 15424 8434
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15488 8090 15516 8366
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 15384 7472 15436 7478
rect 15384 7414 15436 7420
rect 15580 7410 15608 8588
rect 15752 8560 15804 8566
rect 15750 8528 15752 8537
rect 15804 8528 15806 8537
rect 15856 8498 15884 12718
rect 16028 12640 16080 12646
rect 16028 12582 16080 12588
rect 15936 11620 15988 11626
rect 15936 11562 15988 11568
rect 15948 10674 15976 11562
rect 16040 10810 16068 12582
rect 16764 12368 16816 12374
rect 16764 12310 16816 12316
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16500 11694 16528 12174
rect 16592 11898 16620 12174
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16396 11280 16448 11286
rect 16394 11248 16396 11257
rect 16448 11248 16450 11257
rect 16394 11183 16450 11192
rect 16500 11082 16528 11630
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15750 8463 15806 8472
rect 15844 8492 15896 8498
rect 15764 8294 15792 8463
rect 15844 8434 15896 8440
rect 15752 8288 15804 8294
rect 15752 8230 15804 8236
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15764 6934 15792 8026
rect 15856 7954 15884 8434
rect 15948 8294 15976 10610
rect 16040 9926 16068 10746
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16224 10266 16252 10610
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16316 10146 16344 10542
rect 16224 10118 16344 10146
rect 16224 9926 16252 10118
rect 16028 9920 16080 9926
rect 16028 9862 16080 9868
rect 16212 9920 16264 9926
rect 16212 9862 16264 9868
rect 15936 8288 15988 8294
rect 15936 8230 15988 8236
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15752 6928 15804 6934
rect 15752 6870 15804 6876
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15304 6390 15332 6734
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 14924 6248 14976 6254
rect 14924 6190 14976 6196
rect 14520 6012 14828 6021
rect 14520 6010 14526 6012
rect 14582 6010 14606 6012
rect 14662 6010 14686 6012
rect 14742 6010 14766 6012
rect 14822 6010 14828 6012
rect 14582 5958 14584 6010
rect 14764 5958 14766 6010
rect 14520 5956 14526 5958
rect 14582 5956 14606 5958
rect 14662 5956 14686 5958
rect 14742 5956 14766 5958
rect 14822 5956 14828 5958
rect 14520 5947 14828 5956
rect 14936 5794 14964 6190
rect 14844 5766 15056 5794
rect 15120 5778 15148 6258
rect 15200 5840 15252 5846
rect 15200 5782 15252 5788
rect 14844 5710 14872 5766
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14738 5128 14794 5137
rect 14738 5063 14740 5072
rect 14792 5063 14794 5072
rect 14740 5034 14792 5040
rect 14520 4924 14828 4933
rect 14520 4922 14526 4924
rect 14582 4922 14606 4924
rect 14662 4922 14686 4924
rect 14742 4922 14766 4924
rect 14822 4922 14828 4924
rect 14582 4870 14584 4922
rect 14764 4870 14766 4922
rect 14520 4868 14526 4870
rect 14582 4868 14606 4870
rect 14662 4868 14686 4870
rect 14742 4868 14766 4870
rect 14822 4868 14828 4870
rect 14520 4859 14828 4868
rect 14832 4752 14884 4758
rect 14832 4694 14884 4700
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14476 4146 14504 4558
rect 14752 4282 14780 4626
rect 14740 4276 14792 4282
rect 14740 4218 14792 4224
rect 14844 4146 14872 4694
rect 14936 4622 14964 5170
rect 15028 4690 15056 5766
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15108 5636 15160 5642
rect 15108 5578 15160 5584
rect 15120 5302 15148 5578
rect 15108 5296 15160 5302
rect 15108 5238 15160 5244
rect 15016 4684 15068 4690
rect 15016 4626 15068 4632
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 14520 3836 14828 3845
rect 14520 3834 14526 3836
rect 14582 3834 14606 3836
rect 14662 3834 14686 3836
rect 14742 3834 14766 3836
rect 14822 3834 14828 3836
rect 14582 3782 14584 3834
rect 14764 3782 14766 3834
rect 14520 3780 14526 3782
rect 14582 3780 14606 3782
rect 14662 3780 14686 3782
rect 14742 3780 14766 3782
rect 14822 3780 14828 3782
rect 14520 3771 14828 3780
rect 14936 3738 14964 4558
rect 15016 4548 15068 4554
rect 15016 4490 15068 4496
rect 15028 3942 15056 4490
rect 15120 4146 15148 5238
rect 15212 4146 15240 5782
rect 15672 5574 15700 6258
rect 15764 6254 15792 6870
rect 16040 6662 16068 9862
rect 16224 8838 16252 9862
rect 16500 9722 16528 11018
rect 16488 9716 16540 9722
rect 16488 9658 16540 9664
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 16500 8974 16528 9522
rect 16592 9110 16620 11834
rect 16684 11150 16712 12174
rect 16776 11762 16804 12310
rect 16868 12306 16896 13126
rect 16948 12912 17000 12918
rect 16948 12854 17000 12860
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16672 11008 16724 11014
rect 16672 10950 16724 10956
rect 16684 10742 16712 10950
rect 16672 10736 16724 10742
rect 16672 10678 16724 10684
rect 16776 10470 16804 11086
rect 16868 11082 16896 11698
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16764 10464 16816 10470
rect 16764 10406 16816 10412
rect 16868 10282 16896 11018
rect 16960 10674 16988 12854
rect 17052 12850 17080 13330
rect 17234 13084 17542 13093
rect 17234 13082 17240 13084
rect 17296 13082 17320 13084
rect 17376 13082 17400 13084
rect 17456 13082 17480 13084
rect 17536 13082 17542 13084
rect 17296 13030 17298 13082
rect 17478 13030 17480 13082
rect 17234 13028 17240 13030
rect 17296 13028 17320 13030
rect 17376 13028 17400 13030
rect 17456 13028 17480 13030
rect 17536 13028 17542 13030
rect 17234 13019 17542 13028
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17236 12238 17264 12582
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17328 12084 17356 12174
rect 17144 12056 17356 12084
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16948 10532 17000 10538
rect 16948 10474 17000 10480
rect 16684 10254 16896 10282
rect 16684 10062 16712 10254
rect 16960 10130 16988 10474
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16580 9104 16632 9110
rect 16580 9046 16632 9052
rect 16776 9042 16804 9998
rect 16960 9722 16988 10066
rect 17144 9722 17172 12056
rect 17234 11996 17542 12005
rect 17234 11994 17240 11996
rect 17296 11994 17320 11996
rect 17376 11994 17400 11996
rect 17456 11994 17480 11996
rect 17536 11994 17542 11996
rect 17296 11942 17298 11994
rect 17478 11942 17480 11994
rect 17234 11940 17240 11942
rect 17296 11940 17320 11942
rect 17376 11940 17400 11942
rect 17456 11940 17480 11942
rect 17536 11940 17542 11942
rect 17234 11931 17542 11940
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17420 11354 17448 11698
rect 17408 11348 17460 11354
rect 17408 11290 17460 11296
rect 17512 11014 17540 11834
rect 17500 11008 17552 11014
rect 17500 10950 17552 10956
rect 17234 10908 17542 10917
rect 17234 10906 17240 10908
rect 17296 10906 17320 10908
rect 17376 10906 17400 10908
rect 17456 10906 17480 10908
rect 17536 10906 17542 10908
rect 17296 10854 17298 10906
rect 17478 10854 17480 10906
rect 17234 10852 17240 10854
rect 17296 10852 17320 10854
rect 17376 10852 17400 10854
rect 17456 10852 17480 10854
rect 17536 10852 17542 10854
rect 17234 10843 17542 10852
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17420 10470 17448 10610
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17512 10198 17540 10406
rect 17500 10192 17552 10198
rect 17500 10134 17552 10140
rect 17604 10062 17632 13398
rect 17684 13252 17736 13258
rect 17684 13194 17736 13200
rect 17696 12714 17724 13194
rect 17684 12708 17736 12714
rect 17684 12650 17736 12656
rect 17696 12238 17724 12650
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17696 11762 17724 12038
rect 17788 11898 17816 13398
rect 18248 12850 18276 13398
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19524 13320 19576 13326
rect 19524 13262 19576 13268
rect 18512 13252 18564 13258
rect 18512 13194 18564 13200
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 18340 12850 18368 13126
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 17880 12442 17908 12786
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17880 11642 17908 12378
rect 17788 11614 17908 11642
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17696 10169 17724 11154
rect 17788 11150 17816 11614
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 17880 11218 17908 11494
rect 18156 11218 18184 12582
rect 18236 11620 18288 11626
rect 18236 11562 18288 11568
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 18144 11212 18196 11218
rect 18144 11154 18196 11160
rect 18248 11150 18276 11562
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17682 10160 17738 10169
rect 17682 10095 17738 10104
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17234 9820 17542 9829
rect 17234 9818 17240 9820
rect 17296 9818 17320 9820
rect 17376 9818 17400 9820
rect 17456 9818 17480 9820
rect 17536 9818 17542 9820
rect 17296 9766 17298 9818
rect 17478 9766 17480 9818
rect 17234 9764 17240 9766
rect 17296 9764 17320 9766
rect 17376 9764 17400 9766
rect 17456 9764 17480 9766
rect 17536 9764 17542 9766
rect 17234 9755 17542 9764
rect 16948 9716 17000 9722
rect 16948 9658 17000 9664
rect 17132 9716 17184 9722
rect 17132 9658 17184 9664
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16764 9036 16816 9042
rect 16764 8978 16816 8984
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16868 8922 16896 9522
rect 16960 9042 16988 9658
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16224 8022 16252 8774
rect 16500 8566 16528 8910
rect 16868 8906 16988 8922
rect 16868 8900 17000 8906
rect 16868 8894 16948 8900
rect 16948 8842 17000 8848
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16488 8560 16540 8566
rect 16488 8502 16540 8508
rect 16212 8016 16264 8022
rect 16212 7958 16264 7964
rect 16500 6866 16528 8502
rect 16868 8498 16896 8774
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16960 8430 16988 8842
rect 17144 8548 17172 9658
rect 17604 9654 17632 9998
rect 17684 9716 17736 9722
rect 17684 9658 17736 9664
rect 17592 9648 17644 9654
rect 17592 9590 17644 9596
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 17236 8838 17264 9522
rect 17696 9450 17724 9658
rect 17788 9586 17816 10950
rect 17880 10606 17908 11018
rect 17972 10742 18000 11086
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17880 9722 17908 10406
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 17684 9444 17736 9450
rect 17684 9386 17736 9392
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17604 8838 17632 8910
rect 17684 8900 17736 8906
rect 17684 8842 17736 8848
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17234 8732 17542 8741
rect 17234 8730 17240 8732
rect 17296 8730 17320 8732
rect 17376 8730 17400 8732
rect 17456 8730 17480 8732
rect 17536 8730 17542 8732
rect 17296 8678 17298 8730
rect 17478 8678 17480 8730
rect 17234 8676 17240 8678
rect 17296 8676 17320 8678
rect 17376 8676 17400 8678
rect 17456 8676 17480 8678
rect 17536 8676 17542 8678
rect 17234 8667 17542 8676
rect 17604 8634 17632 8774
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17144 8520 17264 8548
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 17236 8276 17264 8520
rect 17696 8498 17724 8842
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17408 8424 17460 8430
rect 17144 8248 17264 8276
rect 17328 8372 17408 8378
rect 17512 8401 17540 8434
rect 17328 8366 17460 8372
rect 17498 8392 17554 8401
rect 17328 8350 17448 8366
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16960 7342 16988 7890
rect 17144 7410 17172 8248
rect 17328 8090 17356 8350
rect 17498 8327 17554 8336
rect 17592 8288 17644 8294
rect 17420 8236 17592 8242
rect 17420 8230 17644 8236
rect 17420 8214 17632 8230
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17420 7954 17448 8214
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17234 7644 17542 7653
rect 17234 7642 17240 7644
rect 17296 7642 17320 7644
rect 17376 7642 17400 7644
rect 17456 7642 17480 7644
rect 17536 7642 17542 7644
rect 17296 7590 17298 7642
rect 17478 7590 17480 7642
rect 17234 7588 17240 7590
rect 17296 7588 17320 7590
rect 17376 7588 17400 7590
rect 17456 7588 17480 7590
rect 17536 7588 17542 7590
rect 17234 7579 17542 7588
rect 17604 7546 17632 8026
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 16776 6322 16804 6666
rect 16960 6458 16988 7278
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 16764 6316 16816 6322
rect 16764 6258 16816 6264
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15764 5642 15792 6190
rect 15948 5914 15976 6258
rect 17052 6186 17080 6734
rect 17144 6458 17172 7346
rect 17592 7336 17644 7342
rect 17592 7278 17644 7284
rect 17604 6866 17632 7278
rect 17696 6866 17724 8434
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17684 6860 17736 6866
rect 17684 6802 17736 6808
rect 17512 6746 17540 6802
rect 17512 6718 17632 6746
rect 17234 6556 17542 6565
rect 17234 6554 17240 6556
rect 17296 6554 17320 6556
rect 17376 6554 17400 6556
rect 17456 6554 17480 6556
rect 17536 6554 17542 6556
rect 17296 6502 17298 6554
rect 17478 6502 17480 6554
rect 17234 6500 17240 6502
rect 17296 6500 17320 6502
rect 17376 6500 17400 6502
rect 17456 6500 17480 6502
rect 17536 6500 17542 6502
rect 17234 6491 17542 6500
rect 17132 6452 17184 6458
rect 17132 6394 17184 6400
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 17040 6180 17092 6186
rect 17040 6122 17092 6128
rect 17052 5914 17080 6122
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 15752 5636 15804 5642
rect 15752 5578 15804 5584
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15672 5302 15700 5510
rect 15660 5296 15712 5302
rect 15660 5238 15712 5244
rect 17144 5250 17172 6258
rect 17234 5468 17542 5477
rect 17234 5466 17240 5468
rect 17296 5466 17320 5468
rect 17376 5466 17400 5468
rect 17456 5466 17480 5468
rect 17536 5466 17542 5468
rect 17296 5414 17298 5466
rect 17478 5414 17480 5466
rect 17234 5412 17240 5414
rect 17296 5412 17320 5414
rect 17376 5412 17400 5414
rect 17456 5412 17480 5414
rect 17536 5412 17542 5414
rect 17234 5403 17542 5412
rect 15672 4826 15700 5238
rect 17144 5234 17264 5250
rect 17144 5228 17276 5234
rect 17144 5222 17224 5228
rect 17224 5170 17276 5176
rect 17132 5160 17184 5166
rect 17132 5102 17184 5108
rect 15660 4820 15712 4826
rect 15660 4762 15712 4768
rect 17144 4758 17172 5102
rect 17604 4826 17632 6718
rect 17788 6322 17816 9318
rect 17880 8480 17908 9522
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18064 8634 18092 9454
rect 18248 9042 18276 11086
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18432 9518 18460 10542
rect 18420 9512 18472 9518
rect 18420 9454 18472 9460
rect 18524 9450 18552 13194
rect 19352 12850 19380 13194
rect 19444 12986 19472 13262
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19444 12850 19472 12922
rect 19536 12918 19564 13262
rect 19524 12912 19576 12918
rect 19524 12854 19576 12860
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 18616 12442 18644 12718
rect 18604 12436 18656 12442
rect 18604 12378 18656 12384
rect 19352 12238 19380 12786
rect 19536 12730 19564 12854
rect 19444 12702 19564 12730
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18708 11150 18736 12038
rect 19340 11620 19392 11626
rect 19340 11562 19392 11568
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 18892 10606 18920 11086
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 19260 10690 19288 10950
rect 19352 10810 19380 11562
rect 19444 10810 19472 12702
rect 19524 12640 19576 12646
rect 19524 12582 19576 12588
rect 19536 11830 19564 12582
rect 19812 12374 19840 13466
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 20536 12980 20588 12986
rect 20536 12922 20588 12928
rect 20352 12912 20404 12918
rect 20352 12854 20404 12860
rect 19948 12540 20256 12549
rect 19948 12538 19954 12540
rect 20010 12538 20034 12540
rect 20090 12538 20114 12540
rect 20170 12538 20194 12540
rect 20250 12538 20256 12540
rect 20010 12486 20012 12538
rect 20192 12486 20194 12538
rect 19948 12484 19954 12486
rect 20010 12484 20034 12486
rect 20090 12484 20114 12486
rect 20170 12484 20194 12486
rect 20250 12484 20256 12486
rect 19948 12475 20256 12484
rect 19708 12368 19760 12374
rect 19708 12310 19760 12316
rect 19800 12368 19852 12374
rect 19800 12310 19852 12316
rect 19524 11824 19576 11830
rect 19524 11766 19576 11772
rect 19524 11688 19576 11694
rect 19524 11630 19576 11636
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19260 10662 19380 10690
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 19248 9716 19300 9722
rect 19248 9658 19300 9664
rect 18788 9580 18840 9586
rect 18788 9522 18840 9528
rect 18512 9444 18564 9450
rect 18512 9386 18564 9392
rect 18236 9036 18288 9042
rect 18236 8978 18288 8984
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 17880 8452 18000 8480
rect 17866 8392 17922 8401
rect 17972 8362 18000 8452
rect 17866 8327 17922 8336
rect 17960 8356 18012 8362
rect 17880 7478 17908 8327
rect 17960 8298 18012 8304
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 17868 7472 17920 7478
rect 17868 7414 17920 7420
rect 17880 7002 17908 7414
rect 17868 6996 17920 7002
rect 17868 6938 17920 6944
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 18156 6118 18184 7686
rect 18248 6322 18276 8978
rect 18800 8906 18828 9522
rect 19260 8974 19288 9658
rect 19352 9178 19380 10662
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 18788 8900 18840 8906
rect 18788 8842 18840 8848
rect 19154 8528 19210 8537
rect 19154 8463 19156 8472
rect 19208 8463 19210 8472
rect 19156 8434 19208 8440
rect 19260 7546 19288 8910
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19352 8498 19380 8774
rect 19340 8492 19392 8498
rect 19340 8434 19392 8440
rect 19352 7546 19380 8434
rect 19444 8090 19472 10610
rect 19536 8634 19564 11630
rect 19616 11552 19668 11558
rect 19616 11494 19668 11500
rect 19628 11150 19656 11494
rect 19720 11150 19748 12310
rect 19812 11218 19840 12310
rect 20168 12300 20220 12306
rect 20168 12242 20220 12248
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 20088 11830 20116 12038
rect 20180 11914 20208 12242
rect 20364 12238 20392 12854
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20456 12306 20484 12718
rect 20444 12300 20496 12306
rect 20444 12242 20496 12248
rect 20352 12232 20404 12238
rect 20352 12174 20404 12180
rect 20548 11914 20576 12922
rect 20640 12850 20668 13126
rect 22662 13084 22970 13093
rect 22662 13082 22668 13084
rect 22724 13082 22748 13084
rect 22804 13082 22828 13084
rect 22884 13082 22908 13084
rect 22964 13082 22970 13084
rect 22724 13030 22726 13082
rect 22906 13030 22908 13082
rect 22662 13028 22668 13030
rect 22724 13028 22748 13030
rect 22804 13028 22828 13030
rect 22884 13028 22908 13030
rect 22964 13028 22970 13030
rect 22662 13019 22970 13028
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 20180 11886 20576 11914
rect 20076 11824 20128 11830
rect 20076 11766 20128 11772
rect 19948 11452 20256 11461
rect 19948 11450 19954 11452
rect 20010 11450 20034 11452
rect 20090 11450 20114 11452
rect 20170 11450 20194 11452
rect 20250 11450 20256 11452
rect 20010 11398 20012 11450
rect 20192 11398 20194 11450
rect 19948 11396 19954 11398
rect 20010 11396 20034 11398
rect 20090 11396 20114 11398
rect 20170 11396 20194 11398
rect 20250 11396 20256 11398
rect 19948 11387 20256 11396
rect 19800 11212 19852 11218
rect 19800 11154 19852 11160
rect 19616 11144 19668 11150
rect 19616 11086 19668 11092
rect 19708 11144 19760 11150
rect 19708 11086 19760 11092
rect 19800 11076 19852 11082
rect 19800 11018 19852 11024
rect 19616 10804 19668 10810
rect 19616 10746 19668 10752
rect 19628 10606 19656 10746
rect 19708 10668 19760 10674
rect 19708 10610 19760 10616
rect 19616 10600 19668 10606
rect 19616 10542 19668 10548
rect 19628 10266 19656 10542
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19524 8628 19576 8634
rect 19524 8570 19576 8576
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19260 7410 19288 7482
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 18604 6724 18656 6730
rect 18604 6666 18656 6672
rect 18616 6458 18644 6666
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 19352 6322 19380 7482
rect 19628 6934 19656 10202
rect 19720 10130 19748 10610
rect 19812 10266 19840 11018
rect 19948 10364 20256 10373
rect 19948 10362 19954 10364
rect 20010 10362 20034 10364
rect 20090 10362 20114 10364
rect 20170 10362 20194 10364
rect 20250 10362 20256 10364
rect 20010 10310 20012 10362
rect 20192 10310 20194 10362
rect 19948 10308 19954 10310
rect 20010 10308 20034 10310
rect 20090 10308 20114 10310
rect 20170 10308 20194 10310
rect 20250 10308 20256 10310
rect 19948 10299 20256 10308
rect 19800 10260 19852 10266
rect 19800 10202 19852 10208
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 20364 10062 20392 11886
rect 20444 11076 20496 11082
rect 20444 11018 20496 11024
rect 19800 10056 19852 10062
rect 19800 9998 19852 10004
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 19708 8424 19760 8430
rect 19708 8366 19760 8372
rect 19720 7750 19748 8366
rect 19708 7744 19760 7750
rect 19708 7686 19760 7692
rect 19616 6928 19668 6934
rect 19616 6870 19668 6876
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 17592 4820 17644 4826
rect 17592 4762 17644 4768
rect 17132 4752 17184 4758
rect 17132 4694 17184 4700
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14384 3058 14412 3470
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 2688 2372 2740 2378
rect 2688 2314 2740 2320
rect 11336 2372 11388 2378
rect 11336 2314 11388 2320
rect 13912 2372 13964 2378
rect 13912 2314 13964 2320
rect 14292 2310 14320 2926
rect 15028 2922 15056 3878
rect 15120 3194 15148 4082
rect 15212 3738 15240 4082
rect 17144 4010 17172 4694
rect 17234 4380 17542 4389
rect 17234 4378 17240 4380
rect 17296 4378 17320 4380
rect 17376 4378 17400 4380
rect 17456 4378 17480 4380
rect 17536 4378 17542 4380
rect 17296 4326 17298 4378
rect 17478 4326 17480 4378
rect 17234 4324 17240 4326
rect 17296 4324 17320 4326
rect 17376 4324 17400 4326
rect 17456 4324 17480 4326
rect 17536 4324 17542 4326
rect 17234 4315 17542 4324
rect 17132 4004 17184 4010
rect 17132 3946 17184 3952
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 19444 3505 19472 6598
rect 19628 6458 19656 6734
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19720 6322 19748 7686
rect 19812 7002 19840 9998
rect 20260 9920 20312 9926
rect 20456 9874 20484 11018
rect 20640 10674 20668 12786
rect 21732 12776 21784 12782
rect 21732 12718 21784 12724
rect 21088 12436 21140 12442
rect 21088 12378 21140 12384
rect 20720 12368 20772 12374
rect 20720 12310 20772 12316
rect 20732 12238 20760 12310
rect 20996 12300 21048 12306
rect 20996 12242 21048 12248
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 20824 11898 20852 12174
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20628 10668 20680 10674
rect 20628 10610 20680 10616
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20260 9862 20312 9868
rect 20272 9450 20300 9862
rect 20364 9846 20484 9874
rect 20260 9444 20312 9450
rect 20260 9386 20312 9392
rect 19948 9276 20256 9285
rect 19948 9274 19954 9276
rect 20010 9274 20034 9276
rect 20090 9274 20114 9276
rect 20170 9274 20194 9276
rect 20250 9274 20256 9276
rect 20010 9222 20012 9274
rect 20192 9222 20194 9274
rect 19948 9220 19954 9222
rect 20010 9220 20034 9222
rect 20090 9220 20114 9222
rect 20170 9220 20194 9222
rect 20250 9220 20256 9222
rect 19948 9211 20256 9220
rect 19948 8188 20256 8197
rect 19948 8186 19954 8188
rect 20010 8186 20034 8188
rect 20090 8186 20114 8188
rect 20170 8186 20194 8188
rect 20250 8186 20256 8188
rect 20010 8134 20012 8186
rect 20192 8134 20194 8186
rect 19948 8132 19954 8134
rect 20010 8132 20034 8134
rect 20090 8132 20114 8134
rect 20170 8132 20194 8134
rect 20250 8132 20256 8134
rect 19948 8123 20256 8132
rect 20364 7970 20392 9846
rect 20444 9104 20496 9110
rect 20444 9046 20496 9052
rect 20456 8634 20484 9046
rect 20444 8628 20496 8634
rect 20444 8570 20496 8576
rect 20272 7942 20392 7970
rect 20272 7426 20300 7942
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 20364 7546 20392 7822
rect 20456 7818 20484 8570
rect 20548 8430 20576 10202
rect 20640 9722 20668 10610
rect 20732 9926 20760 11630
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20628 9716 20680 9722
rect 20628 9658 20680 9664
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20628 9444 20680 9450
rect 20628 9386 20680 9392
rect 20640 8922 20668 9386
rect 20732 9382 20760 9522
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20640 8894 20760 8922
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 20548 8294 20576 8366
rect 20536 8288 20588 8294
rect 20536 8230 20588 8236
rect 20444 7812 20496 7818
rect 20444 7754 20496 7760
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20272 7398 20484 7426
rect 20548 7410 20576 8230
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 19948 7100 20256 7109
rect 19948 7098 19954 7100
rect 20010 7098 20034 7100
rect 20090 7098 20114 7100
rect 20170 7098 20194 7100
rect 20250 7098 20256 7100
rect 20010 7046 20012 7098
rect 20192 7046 20194 7098
rect 19948 7044 19954 7046
rect 20010 7044 20034 7046
rect 20090 7044 20114 7046
rect 20170 7044 20194 7046
rect 20250 7044 20256 7046
rect 19948 7035 20256 7044
rect 19800 6996 19852 7002
rect 19800 6938 19852 6944
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 19720 5370 19748 6258
rect 20364 6254 20392 7142
rect 20456 6322 20484 7398
rect 20536 7404 20588 7410
rect 20536 7346 20588 7352
rect 20640 6866 20668 8774
rect 20732 8566 20760 8894
rect 20824 8566 20852 11834
rect 21008 11762 21036 12242
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 21008 10810 21036 11698
rect 21100 11150 21128 12378
rect 21744 12238 21772 12718
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 21272 12096 21324 12102
rect 21272 12038 21324 12044
rect 21180 11552 21232 11558
rect 21180 11494 21232 11500
rect 21192 11286 21220 11494
rect 21284 11354 21312 12038
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21180 11280 21232 11286
rect 21180 11222 21232 11228
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 21180 11144 21232 11150
rect 21180 11086 21232 11092
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 20996 9648 21048 9654
rect 20996 9590 21048 9596
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 20812 8560 20864 8566
rect 20812 8502 20864 8508
rect 20732 7478 20760 8502
rect 21008 8022 21036 9590
rect 21100 9382 21128 11086
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 21192 8974 21220 11086
rect 21272 10600 21324 10606
rect 21272 10542 21324 10548
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 21284 9994 21312 10542
rect 21272 9988 21324 9994
rect 21272 9930 21324 9936
rect 21284 9586 21312 9930
rect 21560 9654 21588 10542
rect 22020 10470 22048 11086
rect 22204 10674 22232 12786
rect 22662 11996 22970 12005
rect 22662 11994 22668 11996
rect 22724 11994 22748 11996
rect 22804 11994 22828 11996
rect 22884 11994 22908 11996
rect 22964 11994 22970 11996
rect 22724 11942 22726 11994
rect 22906 11942 22908 11994
rect 22662 11940 22668 11942
rect 22724 11940 22748 11942
rect 22804 11940 22828 11942
rect 22884 11940 22908 11942
rect 22964 11940 22970 11942
rect 22662 11931 22970 11940
rect 22662 10908 22970 10917
rect 22662 10906 22668 10908
rect 22724 10906 22748 10908
rect 22804 10906 22828 10908
rect 22884 10906 22908 10908
rect 22964 10906 22970 10908
rect 22724 10854 22726 10906
rect 22906 10854 22908 10906
rect 22662 10852 22668 10854
rect 22724 10852 22748 10854
rect 22804 10852 22828 10854
rect 22884 10852 22908 10854
rect 22964 10852 22970 10854
rect 22662 10843 22970 10852
rect 22192 10668 22244 10674
rect 22192 10610 22244 10616
rect 22008 10464 22060 10470
rect 22008 10406 22060 10412
rect 21548 9648 21600 9654
rect 21548 9590 21600 9596
rect 21272 9580 21324 9586
rect 22020 9568 22048 10406
rect 22662 9820 22970 9829
rect 22662 9818 22668 9820
rect 22724 9818 22748 9820
rect 22804 9818 22828 9820
rect 22884 9818 22908 9820
rect 22964 9818 22970 9820
rect 22724 9766 22726 9818
rect 22906 9766 22908 9818
rect 22662 9764 22668 9766
rect 22724 9764 22748 9766
rect 22804 9764 22828 9766
rect 22884 9764 22908 9766
rect 22964 9764 22970 9766
rect 22662 9755 22970 9764
rect 22100 9580 22152 9586
rect 22020 9540 22100 9568
rect 21272 9522 21324 9528
rect 22100 9522 22152 9528
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 22008 9376 22060 9382
rect 22008 9318 22060 9324
rect 21284 8974 21312 9318
rect 22020 9042 22048 9318
rect 22008 9036 22060 9042
rect 22008 8978 22060 8984
rect 21180 8968 21232 8974
rect 21180 8910 21232 8916
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 22662 8732 22970 8741
rect 22662 8730 22668 8732
rect 22724 8730 22748 8732
rect 22804 8730 22828 8732
rect 22884 8730 22908 8732
rect 22964 8730 22970 8732
rect 22724 8678 22726 8730
rect 22906 8678 22908 8730
rect 22662 8676 22668 8678
rect 22724 8676 22748 8678
rect 22804 8676 22828 8678
rect 22884 8676 22908 8678
rect 22964 8676 22970 8678
rect 22662 8667 22970 8676
rect 20996 8016 21048 8022
rect 20996 7958 21048 7964
rect 22662 7644 22970 7653
rect 22662 7642 22668 7644
rect 22724 7642 22748 7644
rect 22804 7642 22828 7644
rect 22884 7642 22908 7644
rect 22964 7642 22970 7644
rect 22724 7590 22726 7642
rect 22906 7590 22908 7642
rect 22662 7588 22668 7590
rect 22724 7588 22748 7590
rect 22804 7588 22828 7590
rect 22884 7588 22908 7590
rect 22964 7588 22970 7590
rect 22662 7579 22970 7588
rect 20720 7472 20772 7478
rect 20720 7414 20772 7420
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 22662 6556 22970 6565
rect 22662 6554 22668 6556
rect 22724 6554 22748 6556
rect 22804 6554 22828 6556
rect 22884 6554 22908 6556
rect 22964 6554 22970 6556
rect 22724 6502 22726 6554
rect 22906 6502 22908 6554
rect 22662 6500 22668 6502
rect 22724 6500 22748 6502
rect 22804 6500 22828 6502
rect 22884 6500 22908 6502
rect 22964 6500 22970 6502
rect 22662 6491 22970 6500
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20352 6248 20404 6254
rect 20352 6190 20404 6196
rect 19948 6012 20256 6021
rect 19948 6010 19954 6012
rect 20010 6010 20034 6012
rect 20090 6010 20114 6012
rect 20170 6010 20194 6012
rect 20250 6010 20256 6012
rect 20010 5958 20012 6010
rect 20192 5958 20194 6010
rect 19948 5956 19954 5958
rect 20010 5956 20034 5958
rect 20090 5956 20114 5958
rect 20170 5956 20194 5958
rect 20250 5956 20256 5958
rect 19948 5947 20256 5956
rect 22662 5468 22970 5477
rect 22662 5466 22668 5468
rect 22724 5466 22748 5468
rect 22804 5466 22828 5468
rect 22884 5466 22908 5468
rect 22964 5466 22970 5468
rect 22724 5414 22726 5466
rect 22906 5414 22908 5466
rect 22662 5412 22668 5414
rect 22724 5412 22748 5414
rect 22804 5412 22828 5414
rect 22884 5412 22908 5414
rect 22964 5412 22970 5414
rect 22662 5403 22970 5412
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19948 4924 20256 4933
rect 19948 4922 19954 4924
rect 20010 4922 20034 4924
rect 20090 4922 20114 4924
rect 20170 4922 20194 4924
rect 20250 4922 20256 4924
rect 20010 4870 20012 4922
rect 20192 4870 20194 4922
rect 19948 4868 19954 4870
rect 20010 4868 20034 4870
rect 20090 4868 20114 4870
rect 20170 4868 20194 4870
rect 20250 4868 20256 4870
rect 19948 4859 20256 4868
rect 22662 4380 22970 4389
rect 22662 4378 22668 4380
rect 22724 4378 22748 4380
rect 22804 4378 22828 4380
rect 22884 4378 22908 4380
rect 22964 4378 22970 4380
rect 22724 4326 22726 4378
rect 22906 4326 22908 4378
rect 22662 4324 22668 4326
rect 22724 4324 22748 4326
rect 22804 4324 22828 4326
rect 22884 4324 22908 4326
rect 22964 4324 22970 4326
rect 22662 4315 22970 4324
rect 19948 3836 20256 3845
rect 19948 3834 19954 3836
rect 20010 3834 20034 3836
rect 20090 3834 20114 3836
rect 20170 3834 20194 3836
rect 20250 3834 20256 3836
rect 20010 3782 20012 3834
rect 20192 3782 20194 3834
rect 19948 3780 19954 3782
rect 20010 3780 20034 3782
rect 20090 3780 20114 3782
rect 20170 3780 20194 3782
rect 20250 3780 20256 3782
rect 19948 3771 20256 3780
rect 19430 3496 19486 3505
rect 19430 3431 19486 3440
rect 17234 3292 17542 3301
rect 17234 3290 17240 3292
rect 17296 3290 17320 3292
rect 17376 3290 17400 3292
rect 17456 3290 17480 3292
rect 17536 3290 17542 3292
rect 17296 3238 17298 3290
rect 17478 3238 17480 3290
rect 17234 3236 17240 3238
rect 17296 3236 17320 3238
rect 17376 3236 17400 3238
rect 17456 3236 17480 3238
rect 17536 3236 17542 3238
rect 17234 3227 17542 3236
rect 22662 3292 22970 3301
rect 22662 3290 22668 3292
rect 22724 3290 22748 3292
rect 22804 3290 22828 3292
rect 22884 3290 22908 3292
rect 22964 3290 22970 3292
rect 22724 3238 22726 3290
rect 22906 3238 22908 3290
rect 22662 3236 22668 3238
rect 22724 3236 22748 3238
rect 22804 3236 22828 3238
rect 22884 3236 22908 3238
rect 22964 3236 22970 3238
rect 22662 3227 22970 3236
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15016 2916 15068 2922
rect 15016 2858 15068 2864
rect 14520 2748 14828 2757
rect 14520 2746 14526 2748
rect 14582 2746 14606 2748
rect 14662 2746 14686 2748
rect 14742 2746 14766 2748
rect 14822 2746 14828 2748
rect 14582 2694 14584 2746
rect 14764 2694 14766 2746
rect 14520 2692 14526 2694
rect 14582 2692 14606 2694
rect 14662 2692 14686 2694
rect 14742 2692 14766 2694
rect 14822 2692 14828 2694
rect 14520 2683 14828 2692
rect 19948 2748 20256 2757
rect 19948 2746 19954 2748
rect 20010 2746 20034 2748
rect 20090 2746 20114 2748
rect 20170 2746 20194 2748
rect 20250 2746 20256 2748
rect 20010 2694 20012 2746
rect 20192 2694 20194 2746
rect 19948 2692 19954 2694
rect 20010 2692 20034 2694
rect 20090 2692 20114 2694
rect 20170 2692 20194 2694
rect 20250 2692 20256 2694
rect 19948 2683 20256 2692
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 6378 2204 6686 2213
rect 6378 2202 6384 2204
rect 6440 2202 6464 2204
rect 6520 2202 6544 2204
rect 6600 2202 6624 2204
rect 6680 2202 6686 2204
rect 6440 2150 6442 2202
rect 6622 2150 6624 2202
rect 6378 2148 6384 2150
rect 6440 2148 6464 2150
rect 6520 2148 6544 2150
rect 6600 2148 6624 2150
rect 6680 2148 6686 2150
rect 6378 2139 6686 2148
rect 11806 2204 12114 2213
rect 11806 2202 11812 2204
rect 11868 2202 11892 2204
rect 11948 2202 11972 2204
rect 12028 2202 12052 2204
rect 12108 2202 12114 2204
rect 11868 2150 11870 2202
rect 12050 2150 12052 2202
rect 11806 2148 11812 2150
rect 11868 2148 11892 2150
rect 11948 2148 11972 2150
rect 12028 2148 12052 2150
rect 12108 2148 12114 2150
rect 11806 2139 12114 2148
rect 17234 2204 17542 2213
rect 17234 2202 17240 2204
rect 17296 2202 17320 2204
rect 17376 2202 17400 2204
rect 17456 2202 17480 2204
rect 17536 2202 17542 2204
rect 17296 2150 17298 2202
rect 17478 2150 17480 2202
rect 17234 2148 17240 2150
rect 17296 2148 17320 2150
rect 17376 2148 17400 2150
rect 17456 2148 17480 2150
rect 17536 2148 17542 2150
rect 17234 2139 17542 2148
rect 22662 2204 22970 2213
rect 22662 2202 22668 2204
rect 22724 2202 22748 2204
rect 22804 2202 22828 2204
rect 22884 2202 22908 2204
rect 22964 2202 22970 2204
rect 22724 2150 22726 2202
rect 22906 2150 22908 2202
rect 22662 2148 22668 2150
rect 22724 2148 22748 2150
rect 22804 2148 22828 2150
rect 22884 2148 22908 2150
rect 22964 2148 22970 2150
rect 22662 2139 22970 2148
<< via2 >>
rect 6384 21786 6440 21788
rect 6464 21786 6520 21788
rect 6544 21786 6600 21788
rect 6624 21786 6680 21788
rect 6384 21734 6430 21786
rect 6430 21734 6440 21786
rect 6464 21734 6494 21786
rect 6494 21734 6506 21786
rect 6506 21734 6520 21786
rect 6544 21734 6558 21786
rect 6558 21734 6570 21786
rect 6570 21734 6600 21786
rect 6624 21734 6634 21786
rect 6634 21734 6680 21786
rect 6384 21732 6440 21734
rect 6464 21732 6520 21734
rect 6544 21732 6600 21734
rect 6624 21732 6680 21734
rect 11812 21786 11868 21788
rect 11892 21786 11948 21788
rect 11972 21786 12028 21788
rect 12052 21786 12108 21788
rect 11812 21734 11858 21786
rect 11858 21734 11868 21786
rect 11892 21734 11922 21786
rect 11922 21734 11934 21786
rect 11934 21734 11948 21786
rect 11972 21734 11986 21786
rect 11986 21734 11998 21786
rect 11998 21734 12028 21786
rect 12052 21734 12062 21786
rect 12062 21734 12108 21786
rect 11812 21732 11868 21734
rect 11892 21732 11948 21734
rect 11972 21732 12028 21734
rect 12052 21732 12108 21734
rect 17240 21786 17296 21788
rect 17320 21786 17376 21788
rect 17400 21786 17456 21788
rect 17480 21786 17536 21788
rect 17240 21734 17286 21786
rect 17286 21734 17296 21786
rect 17320 21734 17350 21786
rect 17350 21734 17362 21786
rect 17362 21734 17376 21786
rect 17400 21734 17414 21786
rect 17414 21734 17426 21786
rect 17426 21734 17456 21786
rect 17480 21734 17490 21786
rect 17490 21734 17536 21786
rect 17240 21732 17296 21734
rect 17320 21732 17376 21734
rect 17400 21732 17456 21734
rect 17480 21732 17536 21734
rect 22668 21786 22724 21788
rect 22748 21786 22804 21788
rect 22828 21786 22884 21788
rect 22908 21786 22964 21788
rect 22668 21734 22714 21786
rect 22714 21734 22724 21786
rect 22748 21734 22778 21786
rect 22778 21734 22790 21786
rect 22790 21734 22804 21786
rect 22828 21734 22842 21786
rect 22842 21734 22854 21786
rect 22854 21734 22884 21786
rect 22908 21734 22918 21786
rect 22918 21734 22964 21786
rect 22668 21732 22724 21734
rect 22748 21732 22804 21734
rect 22828 21732 22884 21734
rect 22908 21732 22964 21734
rect 3670 21242 3726 21244
rect 3750 21242 3806 21244
rect 3830 21242 3886 21244
rect 3910 21242 3966 21244
rect 3670 21190 3716 21242
rect 3716 21190 3726 21242
rect 3750 21190 3780 21242
rect 3780 21190 3792 21242
rect 3792 21190 3806 21242
rect 3830 21190 3844 21242
rect 3844 21190 3856 21242
rect 3856 21190 3886 21242
rect 3910 21190 3920 21242
rect 3920 21190 3966 21242
rect 3670 21188 3726 21190
rect 3750 21188 3806 21190
rect 3830 21188 3886 21190
rect 3910 21188 3966 21190
rect 9098 21242 9154 21244
rect 9178 21242 9234 21244
rect 9258 21242 9314 21244
rect 9338 21242 9394 21244
rect 9098 21190 9144 21242
rect 9144 21190 9154 21242
rect 9178 21190 9208 21242
rect 9208 21190 9220 21242
rect 9220 21190 9234 21242
rect 9258 21190 9272 21242
rect 9272 21190 9284 21242
rect 9284 21190 9314 21242
rect 9338 21190 9348 21242
rect 9348 21190 9394 21242
rect 9098 21188 9154 21190
rect 9178 21188 9234 21190
rect 9258 21188 9314 21190
rect 9338 21188 9394 21190
rect 14526 21242 14582 21244
rect 14606 21242 14662 21244
rect 14686 21242 14742 21244
rect 14766 21242 14822 21244
rect 14526 21190 14572 21242
rect 14572 21190 14582 21242
rect 14606 21190 14636 21242
rect 14636 21190 14648 21242
rect 14648 21190 14662 21242
rect 14686 21190 14700 21242
rect 14700 21190 14712 21242
rect 14712 21190 14742 21242
rect 14766 21190 14776 21242
rect 14776 21190 14822 21242
rect 14526 21188 14582 21190
rect 14606 21188 14662 21190
rect 14686 21188 14742 21190
rect 14766 21188 14822 21190
rect 19954 21242 20010 21244
rect 20034 21242 20090 21244
rect 20114 21242 20170 21244
rect 20194 21242 20250 21244
rect 19954 21190 20000 21242
rect 20000 21190 20010 21242
rect 20034 21190 20064 21242
rect 20064 21190 20076 21242
rect 20076 21190 20090 21242
rect 20114 21190 20128 21242
rect 20128 21190 20140 21242
rect 20140 21190 20170 21242
rect 20194 21190 20204 21242
rect 20204 21190 20250 21242
rect 19954 21188 20010 21190
rect 20034 21188 20090 21190
rect 20114 21188 20170 21190
rect 20194 21188 20250 21190
rect 6384 20698 6440 20700
rect 6464 20698 6520 20700
rect 6544 20698 6600 20700
rect 6624 20698 6680 20700
rect 6384 20646 6430 20698
rect 6430 20646 6440 20698
rect 6464 20646 6494 20698
rect 6494 20646 6506 20698
rect 6506 20646 6520 20698
rect 6544 20646 6558 20698
rect 6558 20646 6570 20698
rect 6570 20646 6600 20698
rect 6624 20646 6634 20698
rect 6634 20646 6680 20698
rect 6384 20644 6440 20646
rect 6464 20644 6520 20646
rect 6544 20644 6600 20646
rect 6624 20644 6680 20646
rect 11812 20698 11868 20700
rect 11892 20698 11948 20700
rect 11972 20698 12028 20700
rect 12052 20698 12108 20700
rect 11812 20646 11858 20698
rect 11858 20646 11868 20698
rect 11892 20646 11922 20698
rect 11922 20646 11934 20698
rect 11934 20646 11948 20698
rect 11972 20646 11986 20698
rect 11986 20646 11998 20698
rect 11998 20646 12028 20698
rect 12052 20646 12062 20698
rect 12062 20646 12108 20698
rect 11812 20644 11868 20646
rect 11892 20644 11948 20646
rect 11972 20644 12028 20646
rect 12052 20644 12108 20646
rect 17240 20698 17296 20700
rect 17320 20698 17376 20700
rect 17400 20698 17456 20700
rect 17480 20698 17536 20700
rect 17240 20646 17286 20698
rect 17286 20646 17296 20698
rect 17320 20646 17350 20698
rect 17350 20646 17362 20698
rect 17362 20646 17376 20698
rect 17400 20646 17414 20698
rect 17414 20646 17426 20698
rect 17426 20646 17456 20698
rect 17480 20646 17490 20698
rect 17490 20646 17536 20698
rect 17240 20644 17296 20646
rect 17320 20644 17376 20646
rect 17400 20644 17456 20646
rect 17480 20644 17536 20646
rect 22668 20698 22724 20700
rect 22748 20698 22804 20700
rect 22828 20698 22884 20700
rect 22908 20698 22964 20700
rect 22668 20646 22714 20698
rect 22714 20646 22724 20698
rect 22748 20646 22778 20698
rect 22778 20646 22790 20698
rect 22790 20646 22804 20698
rect 22828 20646 22842 20698
rect 22842 20646 22854 20698
rect 22854 20646 22884 20698
rect 22908 20646 22918 20698
rect 22918 20646 22964 20698
rect 22668 20644 22724 20646
rect 22748 20644 22804 20646
rect 22828 20644 22884 20646
rect 22908 20644 22964 20646
rect 3670 20154 3726 20156
rect 3750 20154 3806 20156
rect 3830 20154 3886 20156
rect 3910 20154 3966 20156
rect 3670 20102 3716 20154
rect 3716 20102 3726 20154
rect 3750 20102 3780 20154
rect 3780 20102 3792 20154
rect 3792 20102 3806 20154
rect 3830 20102 3844 20154
rect 3844 20102 3856 20154
rect 3856 20102 3886 20154
rect 3910 20102 3920 20154
rect 3920 20102 3966 20154
rect 3670 20100 3726 20102
rect 3750 20100 3806 20102
rect 3830 20100 3886 20102
rect 3910 20100 3966 20102
rect 9098 20154 9154 20156
rect 9178 20154 9234 20156
rect 9258 20154 9314 20156
rect 9338 20154 9394 20156
rect 9098 20102 9144 20154
rect 9144 20102 9154 20154
rect 9178 20102 9208 20154
rect 9208 20102 9220 20154
rect 9220 20102 9234 20154
rect 9258 20102 9272 20154
rect 9272 20102 9284 20154
rect 9284 20102 9314 20154
rect 9338 20102 9348 20154
rect 9348 20102 9394 20154
rect 9098 20100 9154 20102
rect 9178 20100 9234 20102
rect 9258 20100 9314 20102
rect 9338 20100 9394 20102
rect 14526 20154 14582 20156
rect 14606 20154 14662 20156
rect 14686 20154 14742 20156
rect 14766 20154 14822 20156
rect 14526 20102 14572 20154
rect 14572 20102 14582 20154
rect 14606 20102 14636 20154
rect 14636 20102 14648 20154
rect 14648 20102 14662 20154
rect 14686 20102 14700 20154
rect 14700 20102 14712 20154
rect 14712 20102 14742 20154
rect 14766 20102 14776 20154
rect 14776 20102 14822 20154
rect 14526 20100 14582 20102
rect 14606 20100 14662 20102
rect 14686 20100 14742 20102
rect 14766 20100 14822 20102
rect 19954 20154 20010 20156
rect 20034 20154 20090 20156
rect 20114 20154 20170 20156
rect 20194 20154 20250 20156
rect 19954 20102 20000 20154
rect 20000 20102 20010 20154
rect 20034 20102 20064 20154
rect 20064 20102 20076 20154
rect 20076 20102 20090 20154
rect 20114 20102 20128 20154
rect 20128 20102 20140 20154
rect 20140 20102 20170 20154
rect 20194 20102 20204 20154
rect 20204 20102 20250 20154
rect 19954 20100 20010 20102
rect 20034 20100 20090 20102
rect 20114 20100 20170 20102
rect 20194 20100 20250 20102
rect 938 19796 940 19816
rect 940 19796 992 19816
rect 992 19796 994 19816
rect 938 19760 994 19796
rect 6384 19610 6440 19612
rect 6464 19610 6520 19612
rect 6544 19610 6600 19612
rect 6624 19610 6680 19612
rect 6384 19558 6430 19610
rect 6430 19558 6440 19610
rect 6464 19558 6494 19610
rect 6494 19558 6506 19610
rect 6506 19558 6520 19610
rect 6544 19558 6558 19610
rect 6558 19558 6570 19610
rect 6570 19558 6600 19610
rect 6624 19558 6634 19610
rect 6634 19558 6680 19610
rect 6384 19556 6440 19558
rect 6464 19556 6520 19558
rect 6544 19556 6600 19558
rect 6624 19556 6680 19558
rect 11812 19610 11868 19612
rect 11892 19610 11948 19612
rect 11972 19610 12028 19612
rect 12052 19610 12108 19612
rect 11812 19558 11858 19610
rect 11858 19558 11868 19610
rect 11892 19558 11922 19610
rect 11922 19558 11934 19610
rect 11934 19558 11948 19610
rect 11972 19558 11986 19610
rect 11986 19558 11998 19610
rect 11998 19558 12028 19610
rect 12052 19558 12062 19610
rect 12062 19558 12108 19610
rect 11812 19556 11868 19558
rect 11892 19556 11948 19558
rect 11972 19556 12028 19558
rect 12052 19556 12108 19558
rect 17240 19610 17296 19612
rect 17320 19610 17376 19612
rect 17400 19610 17456 19612
rect 17480 19610 17536 19612
rect 17240 19558 17286 19610
rect 17286 19558 17296 19610
rect 17320 19558 17350 19610
rect 17350 19558 17362 19610
rect 17362 19558 17376 19610
rect 17400 19558 17414 19610
rect 17414 19558 17426 19610
rect 17426 19558 17456 19610
rect 17480 19558 17490 19610
rect 17490 19558 17536 19610
rect 17240 19556 17296 19558
rect 17320 19556 17376 19558
rect 17400 19556 17456 19558
rect 17480 19556 17536 19558
rect 22668 19610 22724 19612
rect 22748 19610 22804 19612
rect 22828 19610 22884 19612
rect 22908 19610 22964 19612
rect 22668 19558 22714 19610
rect 22714 19558 22724 19610
rect 22748 19558 22778 19610
rect 22778 19558 22790 19610
rect 22790 19558 22804 19610
rect 22828 19558 22842 19610
rect 22842 19558 22854 19610
rect 22854 19558 22884 19610
rect 22908 19558 22918 19610
rect 22918 19558 22964 19610
rect 22668 19556 22724 19558
rect 22748 19556 22804 19558
rect 22828 19556 22884 19558
rect 22908 19556 22964 19558
rect 3670 19066 3726 19068
rect 3750 19066 3806 19068
rect 3830 19066 3886 19068
rect 3910 19066 3966 19068
rect 3670 19014 3716 19066
rect 3716 19014 3726 19066
rect 3750 19014 3780 19066
rect 3780 19014 3792 19066
rect 3792 19014 3806 19066
rect 3830 19014 3844 19066
rect 3844 19014 3856 19066
rect 3856 19014 3886 19066
rect 3910 19014 3920 19066
rect 3920 19014 3966 19066
rect 3670 19012 3726 19014
rect 3750 19012 3806 19014
rect 3830 19012 3886 19014
rect 3910 19012 3966 19014
rect 9098 19066 9154 19068
rect 9178 19066 9234 19068
rect 9258 19066 9314 19068
rect 9338 19066 9394 19068
rect 9098 19014 9144 19066
rect 9144 19014 9154 19066
rect 9178 19014 9208 19066
rect 9208 19014 9220 19066
rect 9220 19014 9234 19066
rect 9258 19014 9272 19066
rect 9272 19014 9284 19066
rect 9284 19014 9314 19066
rect 9338 19014 9348 19066
rect 9348 19014 9394 19066
rect 9098 19012 9154 19014
rect 9178 19012 9234 19014
rect 9258 19012 9314 19014
rect 9338 19012 9394 19014
rect 14526 19066 14582 19068
rect 14606 19066 14662 19068
rect 14686 19066 14742 19068
rect 14766 19066 14822 19068
rect 14526 19014 14572 19066
rect 14572 19014 14582 19066
rect 14606 19014 14636 19066
rect 14636 19014 14648 19066
rect 14648 19014 14662 19066
rect 14686 19014 14700 19066
rect 14700 19014 14712 19066
rect 14712 19014 14742 19066
rect 14766 19014 14776 19066
rect 14776 19014 14822 19066
rect 14526 19012 14582 19014
rect 14606 19012 14662 19014
rect 14686 19012 14742 19014
rect 14766 19012 14822 19014
rect 19954 19066 20010 19068
rect 20034 19066 20090 19068
rect 20114 19066 20170 19068
rect 20194 19066 20250 19068
rect 19954 19014 20000 19066
rect 20000 19014 20010 19066
rect 20034 19014 20064 19066
rect 20064 19014 20076 19066
rect 20076 19014 20090 19066
rect 20114 19014 20128 19066
rect 20128 19014 20140 19066
rect 20140 19014 20170 19066
rect 20194 19014 20204 19066
rect 20204 19014 20250 19066
rect 19954 19012 20010 19014
rect 20034 19012 20090 19014
rect 20114 19012 20170 19014
rect 20194 19012 20250 19014
rect 6384 18522 6440 18524
rect 6464 18522 6520 18524
rect 6544 18522 6600 18524
rect 6624 18522 6680 18524
rect 6384 18470 6430 18522
rect 6430 18470 6440 18522
rect 6464 18470 6494 18522
rect 6494 18470 6506 18522
rect 6506 18470 6520 18522
rect 6544 18470 6558 18522
rect 6558 18470 6570 18522
rect 6570 18470 6600 18522
rect 6624 18470 6634 18522
rect 6634 18470 6680 18522
rect 6384 18468 6440 18470
rect 6464 18468 6520 18470
rect 6544 18468 6600 18470
rect 6624 18468 6680 18470
rect 11812 18522 11868 18524
rect 11892 18522 11948 18524
rect 11972 18522 12028 18524
rect 12052 18522 12108 18524
rect 11812 18470 11858 18522
rect 11858 18470 11868 18522
rect 11892 18470 11922 18522
rect 11922 18470 11934 18522
rect 11934 18470 11948 18522
rect 11972 18470 11986 18522
rect 11986 18470 11998 18522
rect 11998 18470 12028 18522
rect 12052 18470 12062 18522
rect 12062 18470 12108 18522
rect 11812 18468 11868 18470
rect 11892 18468 11948 18470
rect 11972 18468 12028 18470
rect 12052 18468 12108 18470
rect 17240 18522 17296 18524
rect 17320 18522 17376 18524
rect 17400 18522 17456 18524
rect 17480 18522 17536 18524
rect 17240 18470 17286 18522
rect 17286 18470 17296 18522
rect 17320 18470 17350 18522
rect 17350 18470 17362 18522
rect 17362 18470 17376 18522
rect 17400 18470 17414 18522
rect 17414 18470 17426 18522
rect 17426 18470 17456 18522
rect 17480 18470 17490 18522
rect 17490 18470 17536 18522
rect 17240 18468 17296 18470
rect 17320 18468 17376 18470
rect 17400 18468 17456 18470
rect 17480 18468 17536 18470
rect 22668 18522 22724 18524
rect 22748 18522 22804 18524
rect 22828 18522 22884 18524
rect 22908 18522 22964 18524
rect 22668 18470 22714 18522
rect 22714 18470 22724 18522
rect 22748 18470 22778 18522
rect 22778 18470 22790 18522
rect 22790 18470 22804 18522
rect 22828 18470 22842 18522
rect 22842 18470 22854 18522
rect 22854 18470 22884 18522
rect 22908 18470 22918 18522
rect 22918 18470 22964 18522
rect 22668 18468 22724 18470
rect 22748 18468 22804 18470
rect 22828 18468 22884 18470
rect 22908 18468 22964 18470
rect 3670 17978 3726 17980
rect 3750 17978 3806 17980
rect 3830 17978 3886 17980
rect 3910 17978 3966 17980
rect 3670 17926 3716 17978
rect 3716 17926 3726 17978
rect 3750 17926 3780 17978
rect 3780 17926 3792 17978
rect 3792 17926 3806 17978
rect 3830 17926 3844 17978
rect 3844 17926 3856 17978
rect 3856 17926 3886 17978
rect 3910 17926 3920 17978
rect 3920 17926 3966 17978
rect 3670 17924 3726 17926
rect 3750 17924 3806 17926
rect 3830 17924 3886 17926
rect 3910 17924 3966 17926
rect 938 11872 994 11928
rect 3670 16890 3726 16892
rect 3750 16890 3806 16892
rect 3830 16890 3886 16892
rect 3910 16890 3966 16892
rect 3670 16838 3716 16890
rect 3716 16838 3726 16890
rect 3750 16838 3780 16890
rect 3780 16838 3792 16890
rect 3792 16838 3806 16890
rect 3830 16838 3844 16890
rect 3844 16838 3856 16890
rect 3856 16838 3886 16890
rect 3910 16838 3920 16890
rect 3920 16838 3966 16890
rect 3670 16836 3726 16838
rect 3750 16836 3806 16838
rect 3830 16836 3886 16838
rect 3910 16836 3966 16838
rect 3670 15802 3726 15804
rect 3750 15802 3806 15804
rect 3830 15802 3886 15804
rect 3910 15802 3966 15804
rect 3670 15750 3716 15802
rect 3716 15750 3726 15802
rect 3750 15750 3780 15802
rect 3780 15750 3792 15802
rect 3792 15750 3806 15802
rect 3830 15750 3844 15802
rect 3844 15750 3856 15802
rect 3856 15750 3886 15802
rect 3910 15750 3920 15802
rect 3920 15750 3966 15802
rect 3670 15748 3726 15750
rect 3750 15748 3806 15750
rect 3830 15748 3886 15750
rect 3910 15748 3966 15750
rect 3670 14714 3726 14716
rect 3750 14714 3806 14716
rect 3830 14714 3886 14716
rect 3910 14714 3966 14716
rect 3670 14662 3716 14714
rect 3716 14662 3726 14714
rect 3750 14662 3780 14714
rect 3780 14662 3792 14714
rect 3792 14662 3806 14714
rect 3830 14662 3844 14714
rect 3844 14662 3856 14714
rect 3856 14662 3886 14714
rect 3910 14662 3920 14714
rect 3920 14662 3966 14714
rect 3670 14660 3726 14662
rect 3750 14660 3806 14662
rect 3830 14660 3886 14662
rect 3910 14660 3966 14662
rect 3670 13626 3726 13628
rect 3750 13626 3806 13628
rect 3830 13626 3886 13628
rect 3910 13626 3966 13628
rect 3670 13574 3716 13626
rect 3716 13574 3726 13626
rect 3750 13574 3780 13626
rect 3780 13574 3792 13626
rect 3792 13574 3806 13626
rect 3830 13574 3844 13626
rect 3844 13574 3856 13626
rect 3856 13574 3886 13626
rect 3910 13574 3920 13626
rect 3920 13574 3966 13626
rect 3670 13572 3726 13574
rect 3750 13572 3806 13574
rect 3830 13572 3886 13574
rect 3910 13572 3966 13574
rect 3670 12538 3726 12540
rect 3750 12538 3806 12540
rect 3830 12538 3886 12540
rect 3910 12538 3966 12540
rect 3670 12486 3716 12538
rect 3716 12486 3726 12538
rect 3750 12486 3780 12538
rect 3780 12486 3792 12538
rect 3792 12486 3806 12538
rect 3830 12486 3844 12538
rect 3844 12486 3856 12538
rect 3856 12486 3886 12538
rect 3910 12486 3920 12538
rect 3920 12486 3966 12538
rect 3670 12484 3726 12486
rect 3750 12484 3806 12486
rect 3830 12484 3886 12486
rect 3910 12484 3966 12486
rect 3670 11450 3726 11452
rect 3750 11450 3806 11452
rect 3830 11450 3886 11452
rect 3910 11450 3966 11452
rect 3670 11398 3716 11450
rect 3716 11398 3726 11450
rect 3750 11398 3780 11450
rect 3780 11398 3792 11450
rect 3792 11398 3806 11450
rect 3830 11398 3844 11450
rect 3844 11398 3856 11450
rect 3856 11398 3886 11450
rect 3910 11398 3920 11450
rect 3920 11398 3966 11450
rect 3670 11396 3726 11398
rect 3750 11396 3806 11398
rect 3830 11396 3886 11398
rect 3910 11396 3966 11398
rect 3670 10362 3726 10364
rect 3750 10362 3806 10364
rect 3830 10362 3886 10364
rect 3910 10362 3966 10364
rect 3670 10310 3716 10362
rect 3716 10310 3726 10362
rect 3750 10310 3780 10362
rect 3780 10310 3792 10362
rect 3792 10310 3806 10362
rect 3830 10310 3844 10362
rect 3844 10310 3856 10362
rect 3856 10310 3886 10362
rect 3910 10310 3920 10362
rect 3920 10310 3966 10362
rect 3670 10308 3726 10310
rect 3750 10308 3806 10310
rect 3830 10308 3886 10310
rect 3910 10308 3966 10310
rect 3670 9274 3726 9276
rect 3750 9274 3806 9276
rect 3830 9274 3886 9276
rect 3910 9274 3966 9276
rect 3670 9222 3716 9274
rect 3716 9222 3726 9274
rect 3750 9222 3780 9274
rect 3780 9222 3792 9274
rect 3792 9222 3806 9274
rect 3830 9222 3844 9274
rect 3844 9222 3856 9274
rect 3856 9222 3886 9274
rect 3910 9222 3920 9274
rect 3920 9222 3966 9274
rect 3670 9220 3726 9222
rect 3750 9220 3806 9222
rect 3830 9220 3886 9222
rect 3910 9220 3966 9222
rect 6384 17434 6440 17436
rect 6464 17434 6520 17436
rect 6544 17434 6600 17436
rect 6624 17434 6680 17436
rect 6384 17382 6430 17434
rect 6430 17382 6440 17434
rect 6464 17382 6494 17434
rect 6494 17382 6506 17434
rect 6506 17382 6520 17434
rect 6544 17382 6558 17434
rect 6558 17382 6570 17434
rect 6570 17382 6600 17434
rect 6624 17382 6634 17434
rect 6634 17382 6680 17434
rect 6384 17380 6440 17382
rect 6464 17380 6520 17382
rect 6544 17380 6600 17382
rect 6624 17380 6680 17382
rect 3670 8186 3726 8188
rect 3750 8186 3806 8188
rect 3830 8186 3886 8188
rect 3910 8186 3966 8188
rect 3670 8134 3716 8186
rect 3716 8134 3726 8186
rect 3750 8134 3780 8186
rect 3780 8134 3792 8186
rect 3792 8134 3806 8186
rect 3830 8134 3844 8186
rect 3844 8134 3856 8186
rect 3856 8134 3886 8186
rect 3910 8134 3920 8186
rect 3920 8134 3966 8186
rect 3670 8132 3726 8134
rect 3750 8132 3806 8134
rect 3830 8132 3886 8134
rect 3910 8132 3966 8134
rect 3670 7098 3726 7100
rect 3750 7098 3806 7100
rect 3830 7098 3886 7100
rect 3910 7098 3966 7100
rect 3670 7046 3716 7098
rect 3716 7046 3726 7098
rect 3750 7046 3780 7098
rect 3780 7046 3792 7098
rect 3792 7046 3806 7098
rect 3830 7046 3844 7098
rect 3844 7046 3856 7098
rect 3856 7046 3886 7098
rect 3910 7046 3920 7098
rect 3920 7046 3966 7098
rect 3670 7044 3726 7046
rect 3750 7044 3806 7046
rect 3830 7044 3886 7046
rect 3910 7044 3966 7046
rect 3670 6010 3726 6012
rect 3750 6010 3806 6012
rect 3830 6010 3886 6012
rect 3910 6010 3966 6012
rect 3670 5958 3716 6010
rect 3716 5958 3726 6010
rect 3750 5958 3780 6010
rect 3780 5958 3792 6010
rect 3792 5958 3806 6010
rect 3830 5958 3844 6010
rect 3844 5958 3856 6010
rect 3856 5958 3886 6010
rect 3910 5958 3920 6010
rect 3920 5958 3966 6010
rect 3670 5956 3726 5958
rect 3750 5956 3806 5958
rect 3830 5956 3886 5958
rect 3910 5956 3966 5958
rect 6384 16346 6440 16348
rect 6464 16346 6520 16348
rect 6544 16346 6600 16348
rect 6624 16346 6680 16348
rect 6384 16294 6430 16346
rect 6430 16294 6440 16346
rect 6464 16294 6494 16346
rect 6494 16294 6506 16346
rect 6506 16294 6520 16346
rect 6544 16294 6558 16346
rect 6558 16294 6570 16346
rect 6570 16294 6600 16346
rect 6624 16294 6634 16346
rect 6634 16294 6680 16346
rect 6384 16292 6440 16294
rect 6464 16292 6520 16294
rect 6544 16292 6600 16294
rect 6624 16292 6680 16294
rect 6384 15258 6440 15260
rect 6464 15258 6520 15260
rect 6544 15258 6600 15260
rect 6624 15258 6680 15260
rect 6384 15206 6430 15258
rect 6430 15206 6440 15258
rect 6464 15206 6494 15258
rect 6494 15206 6506 15258
rect 6506 15206 6520 15258
rect 6544 15206 6558 15258
rect 6558 15206 6570 15258
rect 6570 15206 6600 15258
rect 6624 15206 6634 15258
rect 6634 15206 6680 15258
rect 6384 15204 6440 15206
rect 6464 15204 6520 15206
rect 6544 15204 6600 15206
rect 6624 15204 6680 15206
rect 3670 4922 3726 4924
rect 3750 4922 3806 4924
rect 3830 4922 3886 4924
rect 3910 4922 3966 4924
rect 3670 4870 3716 4922
rect 3716 4870 3726 4922
rect 3750 4870 3780 4922
rect 3780 4870 3792 4922
rect 3792 4870 3806 4922
rect 3830 4870 3844 4922
rect 3844 4870 3856 4922
rect 3856 4870 3886 4922
rect 3910 4870 3920 4922
rect 3920 4870 3966 4922
rect 3670 4868 3726 4870
rect 3750 4868 3806 4870
rect 3830 4868 3886 4870
rect 3910 4868 3966 4870
rect 3146 3984 3202 4040
rect 3670 3834 3726 3836
rect 3750 3834 3806 3836
rect 3830 3834 3886 3836
rect 3910 3834 3966 3836
rect 3670 3782 3716 3834
rect 3716 3782 3726 3834
rect 3750 3782 3780 3834
rect 3780 3782 3792 3834
rect 3792 3782 3806 3834
rect 3830 3782 3844 3834
rect 3844 3782 3856 3834
rect 3856 3782 3886 3834
rect 3910 3782 3920 3834
rect 3920 3782 3966 3834
rect 3670 3780 3726 3782
rect 3750 3780 3806 3782
rect 3830 3780 3886 3782
rect 3910 3780 3966 3782
rect 3670 2746 3726 2748
rect 3750 2746 3806 2748
rect 3830 2746 3886 2748
rect 3910 2746 3966 2748
rect 3670 2694 3716 2746
rect 3716 2694 3726 2746
rect 3750 2694 3780 2746
rect 3780 2694 3792 2746
rect 3792 2694 3806 2746
rect 3830 2694 3844 2746
rect 3844 2694 3856 2746
rect 3856 2694 3886 2746
rect 3910 2694 3920 2746
rect 3920 2694 3966 2746
rect 3670 2692 3726 2694
rect 3750 2692 3806 2694
rect 3830 2692 3886 2694
rect 3910 2692 3966 2694
rect 6384 14170 6440 14172
rect 6464 14170 6520 14172
rect 6544 14170 6600 14172
rect 6624 14170 6680 14172
rect 6384 14118 6430 14170
rect 6430 14118 6440 14170
rect 6464 14118 6494 14170
rect 6494 14118 6506 14170
rect 6506 14118 6520 14170
rect 6544 14118 6558 14170
rect 6558 14118 6570 14170
rect 6570 14118 6600 14170
rect 6624 14118 6634 14170
rect 6634 14118 6680 14170
rect 6384 14116 6440 14118
rect 6464 14116 6520 14118
rect 6544 14116 6600 14118
rect 6624 14116 6680 14118
rect 9098 17978 9154 17980
rect 9178 17978 9234 17980
rect 9258 17978 9314 17980
rect 9338 17978 9394 17980
rect 9098 17926 9144 17978
rect 9144 17926 9154 17978
rect 9178 17926 9208 17978
rect 9208 17926 9220 17978
rect 9220 17926 9234 17978
rect 9258 17926 9272 17978
rect 9272 17926 9284 17978
rect 9284 17926 9314 17978
rect 9338 17926 9348 17978
rect 9348 17926 9394 17978
rect 9098 17924 9154 17926
rect 9178 17924 9234 17926
rect 9258 17924 9314 17926
rect 9338 17924 9394 17926
rect 14526 17978 14582 17980
rect 14606 17978 14662 17980
rect 14686 17978 14742 17980
rect 14766 17978 14822 17980
rect 14526 17926 14572 17978
rect 14572 17926 14582 17978
rect 14606 17926 14636 17978
rect 14636 17926 14648 17978
rect 14648 17926 14662 17978
rect 14686 17926 14700 17978
rect 14700 17926 14712 17978
rect 14712 17926 14742 17978
rect 14766 17926 14776 17978
rect 14776 17926 14822 17978
rect 14526 17924 14582 17926
rect 14606 17924 14662 17926
rect 14686 17924 14742 17926
rect 14766 17924 14822 17926
rect 19954 17978 20010 17980
rect 20034 17978 20090 17980
rect 20114 17978 20170 17980
rect 20194 17978 20250 17980
rect 19954 17926 20000 17978
rect 20000 17926 20010 17978
rect 20034 17926 20064 17978
rect 20064 17926 20076 17978
rect 20076 17926 20090 17978
rect 20114 17926 20128 17978
rect 20128 17926 20140 17978
rect 20140 17926 20170 17978
rect 20194 17926 20204 17978
rect 20204 17926 20250 17978
rect 19954 17924 20010 17926
rect 20034 17924 20090 17926
rect 20114 17924 20170 17926
rect 20194 17924 20250 17926
rect 9098 16890 9154 16892
rect 9178 16890 9234 16892
rect 9258 16890 9314 16892
rect 9338 16890 9394 16892
rect 9098 16838 9144 16890
rect 9144 16838 9154 16890
rect 9178 16838 9208 16890
rect 9208 16838 9220 16890
rect 9220 16838 9234 16890
rect 9258 16838 9272 16890
rect 9272 16838 9284 16890
rect 9284 16838 9314 16890
rect 9338 16838 9348 16890
rect 9348 16838 9394 16890
rect 9098 16836 9154 16838
rect 9178 16836 9234 16838
rect 9258 16836 9314 16838
rect 9338 16836 9394 16838
rect 9098 15802 9154 15804
rect 9178 15802 9234 15804
rect 9258 15802 9314 15804
rect 9338 15802 9394 15804
rect 9098 15750 9144 15802
rect 9144 15750 9154 15802
rect 9178 15750 9208 15802
rect 9208 15750 9220 15802
rect 9220 15750 9234 15802
rect 9258 15750 9272 15802
rect 9272 15750 9284 15802
rect 9284 15750 9314 15802
rect 9338 15750 9348 15802
rect 9348 15750 9394 15802
rect 9098 15748 9154 15750
rect 9178 15748 9234 15750
rect 9258 15748 9314 15750
rect 9338 15748 9394 15750
rect 6384 13082 6440 13084
rect 6464 13082 6520 13084
rect 6544 13082 6600 13084
rect 6624 13082 6680 13084
rect 6384 13030 6430 13082
rect 6430 13030 6440 13082
rect 6464 13030 6494 13082
rect 6494 13030 6506 13082
rect 6506 13030 6520 13082
rect 6544 13030 6558 13082
rect 6558 13030 6570 13082
rect 6570 13030 6600 13082
rect 6624 13030 6634 13082
rect 6634 13030 6680 13082
rect 6384 13028 6440 13030
rect 6464 13028 6520 13030
rect 6544 13028 6600 13030
rect 6624 13028 6680 13030
rect 6384 11994 6440 11996
rect 6464 11994 6520 11996
rect 6544 11994 6600 11996
rect 6624 11994 6680 11996
rect 6384 11942 6430 11994
rect 6430 11942 6440 11994
rect 6464 11942 6494 11994
rect 6494 11942 6506 11994
rect 6506 11942 6520 11994
rect 6544 11942 6558 11994
rect 6558 11942 6570 11994
rect 6570 11942 6600 11994
rect 6624 11942 6634 11994
rect 6634 11942 6680 11994
rect 6384 11940 6440 11942
rect 6464 11940 6520 11942
rect 6544 11940 6600 11942
rect 6624 11940 6680 11942
rect 6384 10906 6440 10908
rect 6464 10906 6520 10908
rect 6544 10906 6600 10908
rect 6624 10906 6680 10908
rect 6384 10854 6430 10906
rect 6430 10854 6440 10906
rect 6464 10854 6494 10906
rect 6494 10854 6506 10906
rect 6506 10854 6520 10906
rect 6544 10854 6558 10906
rect 6558 10854 6570 10906
rect 6570 10854 6600 10906
rect 6624 10854 6634 10906
rect 6634 10854 6680 10906
rect 6384 10852 6440 10854
rect 6464 10852 6520 10854
rect 6544 10852 6600 10854
rect 6624 10852 6680 10854
rect 6384 9818 6440 9820
rect 6464 9818 6520 9820
rect 6544 9818 6600 9820
rect 6624 9818 6680 9820
rect 6384 9766 6430 9818
rect 6430 9766 6440 9818
rect 6464 9766 6494 9818
rect 6494 9766 6506 9818
rect 6506 9766 6520 9818
rect 6544 9766 6558 9818
rect 6558 9766 6570 9818
rect 6570 9766 6600 9818
rect 6624 9766 6634 9818
rect 6634 9766 6680 9818
rect 6384 9764 6440 9766
rect 6464 9764 6520 9766
rect 6544 9764 6600 9766
rect 6624 9764 6680 9766
rect 6384 8730 6440 8732
rect 6464 8730 6520 8732
rect 6544 8730 6600 8732
rect 6624 8730 6680 8732
rect 6384 8678 6430 8730
rect 6430 8678 6440 8730
rect 6464 8678 6494 8730
rect 6494 8678 6506 8730
rect 6506 8678 6520 8730
rect 6544 8678 6558 8730
rect 6558 8678 6570 8730
rect 6570 8678 6600 8730
rect 6624 8678 6634 8730
rect 6634 8678 6680 8730
rect 6384 8676 6440 8678
rect 6464 8676 6520 8678
rect 6544 8676 6600 8678
rect 6624 8676 6680 8678
rect 11812 17434 11868 17436
rect 11892 17434 11948 17436
rect 11972 17434 12028 17436
rect 12052 17434 12108 17436
rect 11812 17382 11858 17434
rect 11858 17382 11868 17434
rect 11892 17382 11922 17434
rect 11922 17382 11934 17434
rect 11934 17382 11948 17434
rect 11972 17382 11986 17434
rect 11986 17382 11998 17434
rect 11998 17382 12028 17434
rect 12052 17382 12062 17434
rect 12062 17382 12108 17434
rect 11812 17380 11868 17382
rect 11892 17380 11948 17382
rect 11972 17380 12028 17382
rect 12052 17380 12108 17382
rect 17240 17434 17296 17436
rect 17320 17434 17376 17436
rect 17400 17434 17456 17436
rect 17480 17434 17536 17436
rect 17240 17382 17286 17434
rect 17286 17382 17296 17434
rect 17320 17382 17350 17434
rect 17350 17382 17362 17434
rect 17362 17382 17376 17434
rect 17400 17382 17414 17434
rect 17414 17382 17426 17434
rect 17426 17382 17456 17434
rect 17480 17382 17490 17434
rect 17490 17382 17536 17434
rect 17240 17380 17296 17382
rect 17320 17380 17376 17382
rect 17400 17380 17456 17382
rect 17480 17380 17536 17382
rect 22668 17434 22724 17436
rect 22748 17434 22804 17436
rect 22828 17434 22884 17436
rect 22908 17434 22964 17436
rect 22668 17382 22714 17434
rect 22714 17382 22724 17434
rect 22748 17382 22778 17434
rect 22778 17382 22790 17434
rect 22790 17382 22804 17434
rect 22828 17382 22842 17434
rect 22842 17382 22854 17434
rect 22854 17382 22884 17434
rect 22908 17382 22918 17434
rect 22918 17382 22964 17434
rect 22668 17380 22724 17382
rect 22748 17380 22804 17382
rect 22828 17380 22884 17382
rect 22908 17380 22964 17382
rect 6384 7642 6440 7644
rect 6464 7642 6520 7644
rect 6544 7642 6600 7644
rect 6624 7642 6680 7644
rect 6384 7590 6430 7642
rect 6430 7590 6440 7642
rect 6464 7590 6494 7642
rect 6494 7590 6506 7642
rect 6506 7590 6520 7642
rect 6544 7590 6558 7642
rect 6558 7590 6570 7642
rect 6570 7590 6600 7642
rect 6624 7590 6634 7642
rect 6634 7590 6680 7642
rect 6384 7588 6440 7590
rect 6464 7588 6520 7590
rect 6544 7588 6600 7590
rect 6624 7588 6680 7590
rect 6384 6554 6440 6556
rect 6464 6554 6520 6556
rect 6544 6554 6600 6556
rect 6624 6554 6680 6556
rect 6384 6502 6430 6554
rect 6430 6502 6440 6554
rect 6464 6502 6494 6554
rect 6494 6502 6506 6554
rect 6506 6502 6520 6554
rect 6544 6502 6558 6554
rect 6558 6502 6570 6554
rect 6570 6502 6600 6554
rect 6624 6502 6634 6554
rect 6634 6502 6680 6554
rect 6384 6500 6440 6502
rect 6464 6500 6520 6502
rect 6544 6500 6600 6502
rect 6624 6500 6680 6502
rect 6384 5466 6440 5468
rect 6464 5466 6520 5468
rect 6544 5466 6600 5468
rect 6624 5466 6680 5468
rect 6384 5414 6430 5466
rect 6430 5414 6440 5466
rect 6464 5414 6494 5466
rect 6494 5414 6506 5466
rect 6506 5414 6520 5466
rect 6544 5414 6558 5466
rect 6558 5414 6570 5466
rect 6570 5414 6600 5466
rect 6624 5414 6634 5466
rect 6634 5414 6680 5466
rect 6384 5412 6440 5414
rect 6464 5412 6520 5414
rect 6544 5412 6600 5414
rect 6624 5412 6680 5414
rect 9098 14714 9154 14716
rect 9178 14714 9234 14716
rect 9258 14714 9314 14716
rect 9338 14714 9394 14716
rect 9098 14662 9144 14714
rect 9144 14662 9154 14714
rect 9178 14662 9208 14714
rect 9208 14662 9220 14714
rect 9220 14662 9234 14714
rect 9258 14662 9272 14714
rect 9272 14662 9284 14714
rect 9284 14662 9314 14714
rect 9338 14662 9348 14714
rect 9348 14662 9394 14714
rect 9098 14660 9154 14662
rect 9178 14660 9234 14662
rect 9258 14660 9314 14662
rect 9338 14660 9394 14662
rect 14526 16890 14582 16892
rect 14606 16890 14662 16892
rect 14686 16890 14742 16892
rect 14766 16890 14822 16892
rect 14526 16838 14572 16890
rect 14572 16838 14582 16890
rect 14606 16838 14636 16890
rect 14636 16838 14648 16890
rect 14648 16838 14662 16890
rect 14686 16838 14700 16890
rect 14700 16838 14712 16890
rect 14712 16838 14742 16890
rect 14766 16838 14776 16890
rect 14776 16838 14822 16890
rect 14526 16836 14582 16838
rect 14606 16836 14662 16838
rect 14686 16836 14742 16838
rect 14766 16836 14822 16838
rect 19954 16890 20010 16892
rect 20034 16890 20090 16892
rect 20114 16890 20170 16892
rect 20194 16890 20250 16892
rect 19954 16838 20000 16890
rect 20000 16838 20010 16890
rect 20034 16838 20064 16890
rect 20064 16838 20076 16890
rect 20076 16838 20090 16890
rect 20114 16838 20128 16890
rect 20128 16838 20140 16890
rect 20140 16838 20170 16890
rect 20194 16838 20204 16890
rect 20204 16838 20250 16890
rect 19954 16836 20010 16838
rect 20034 16836 20090 16838
rect 20114 16836 20170 16838
rect 20194 16836 20250 16838
rect 11812 16346 11868 16348
rect 11892 16346 11948 16348
rect 11972 16346 12028 16348
rect 12052 16346 12108 16348
rect 11812 16294 11858 16346
rect 11858 16294 11868 16346
rect 11892 16294 11922 16346
rect 11922 16294 11934 16346
rect 11934 16294 11948 16346
rect 11972 16294 11986 16346
rect 11986 16294 11998 16346
rect 11998 16294 12028 16346
rect 12052 16294 12062 16346
rect 12062 16294 12108 16346
rect 11812 16292 11868 16294
rect 11892 16292 11948 16294
rect 11972 16292 12028 16294
rect 12052 16292 12108 16294
rect 17240 16346 17296 16348
rect 17320 16346 17376 16348
rect 17400 16346 17456 16348
rect 17480 16346 17536 16348
rect 17240 16294 17286 16346
rect 17286 16294 17296 16346
rect 17320 16294 17350 16346
rect 17350 16294 17362 16346
rect 17362 16294 17376 16346
rect 17400 16294 17414 16346
rect 17414 16294 17426 16346
rect 17426 16294 17456 16346
rect 17480 16294 17490 16346
rect 17490 16294 17536 16346
rect 17240 16292 17296 16294
rect 17320 16292 17376 16294
rect 17400 16292 17456 16294
rect 17480 16292 17536 16294
rect 22668 16346 22724 16348
rect 22748 16346 22804 16348
rect 22828 16346 22884 16348
rect 22908 16346 22964 16348
rect 22668 16294 22714 16346
rect 22714 16294 22724 16346
rect 22748 16294 22778 16346
rect 22778 16294 22790 16346
rect 22790 16294 22804 16346
rect 22828 16294 22842 16346
rect 22842 16294 22854 16346
rect 22854 16294 22884 16346
rect 22908 16294 22918 16346
rect 22918 16294 22964 16346
rect 22668 16292 22724 16294
rect 22748 16292 22804 16294
rect 22828 16292 22884 16294
rect 22908 16292 22964 16294
rect 9098 13626 9154 13628
rect 9178 13626 9234 13628
rect 9258 13626 9314 13628
rect 9338 13626 9394 13628
rect 9098 13574 9144 13626
rect 9144 13574 9154 13626
rect 9178 13574 9208 13626
rect 9208 13574 9220 13626
rect 9220 13574 9234 13626
rect 9258 13574 9272 13626
rect 9272 13574 9284 13626
rect 9284 13574 9314 13626
rect 9338 13574 9348 13626
rect 9348 13574 9394 13626
rect 9098 13572 9154 13574
rect 9178 13572 9234 13574
rect 9258 13572 9314 13574
rect 9338 13572 9394 13574
rect 9098 12538 9154 12540
rect 9178 12538 9234 12540
rect 9258 12538 9314 12540
rect 9338 12538 9394 12540
rect 9098 12486 9144 12538
rect 9144 12486 9154 12538
rect 9178 12486 9208 12538
rect 9208 12486 9220 12538
rect 9220 12486 9234 12538
rect 9258 12486 9272 12538
rect 9272 12486 9284 12538
rect 9284 12486 9314 12538
rect 9338 12486 9348 12538
rect 9348 12486 9394 12538
rect 9098 12484 9154 12486
rect 9178 12484 9234 12486
rect 9258 12484 9314 12486
rect 9338 12484 9394 12486
rect 9098 11450 9154 11452
rect 9178 11450 9234 11452
rect 9258 11450 9314 11452
rect 9338 11450 9394 11452
rect 9098 11398 9144 11450
rect 9144 11398 9154 11450
rect 9178 11398 9208 11450
rect 9208 11398 9220 11450
rect 9220 11398 9234 11450
rect 9258 11398 9272 11450
rect 9272 11398 9284 11450
rect 9284 11398 9314 11450
rect 9338 11398 9348 11450
rect 9348 11398 9394 11450
rect 9098 11396 9154 11398
rect 9178 11396 9234 11398
rect 9258 11396 9314 11398
rect 9338 11396 9394 11398
rect 9098 10362 9154 10364
rect 9178 10362 9234 10364
rect 9258 10362 9314 10364
rect 9338 10362 9394 10364
rect 9098 10310 9144 10362
rect 9144 10310 9154 10362
rect 9178 10310 9208 10362
rect 9208 10310 9220 10362
rect 9220 10310 9234 10362
rect 9258 10310 9272 10362
rect 9272 10310 9284 10362
rect 9284 10310 9314 10362
rect 9338 10310 9348 10362
rect 9348 10310 9394 10362
rect 9098 10308 9154 10310
rect 9178 10308 9234 10310
rect 9258 10308 9314 10310
rect 9338 10308 9394 10310
rect 11812 15258 11868 15260
rect 11892 15258 11948 15260
rect 11972 15258 12028 15260
rect 12052 15258 12108 15260
rect 11812 15206 11858 15258
rect 11858 15206 11868 15258
rect 11892 15206 11922 15258
rect 11922 15206 11934 15258
rect 11934 15206 11948 15258
rect 11972 15206 11986 15258
rect 11986 15206 11998 15258
rect 11998 15206 12028 15258
rect 12052 15206 12062 15258
rect 12062 15206 12108 15258
rect 11812 15204 11868 15206
rect 11892 15204 11948 15206
rect 11972 15204 12028 15206
rect 12052 15204 12108 15206
rect 9098 9274 9154 9276
rect 9178 9274 9234 9276
rect 9258 9274 9314 9276
rect 9338 9274 9394 9276
rect 9098 9222 9144 9274
rect 9144 9222 9154 9274
rect 9178 9222 9208 9274
rect 9208 9222 9220 9274
rect 9220 9222 9234 9274
rect 9258 9222 9272 9274
rect 9272 9222 9284 9274
rect 9284 9222 9314 9274
rect 9338 9222 9348 9274
rect 9348 9222 9394 9274
rect 9098 9220 9154 9222
rect 9178 9220 9234 9222
rect 9258 9220 9314 9222
rect 9338 9220 9394 9222
rect 9098 8186 9154 8188
rect 9178 8186 9234 8188
rect 9258 8186 9314 8188
rect 9338 8186 9394 8188
rect 9098 8134 9144 8186
rect 9144 8134 9154 8186
rect 9178 8134 9208 8186
rect 9208 8134 9220 8186
rect 9220 8134 9234 8186
rect 9258 8134 9272 8186
rect 9272 8134 9284 8186
rect 9284 8134 9314 8186
rect 9338 8134 9348 8186
rect 9348 8134 9394 8186
rect 9098 8132 9154 8134
rect 9178 8132 9234 8134
rect 9258 8132 9314 8134
rect 9338 8132 9394 8134
rect 9098 7098 9154 7100
rect 9178 7098 9234 7100
rect 9258 7098 9314 7100
rect 9338 7098 9394 7100
rect 9098 7046 9144 7098
rect 9144 7046 9154 7098
rect 9178 7046 9208 7098
rect 9208 7046 9220 7098
rect 9220 7046 9234 7098
rect 9258 7046 9272 7098
rect 9272 7046 9284 7098
rect 9284 7046 9314 7098
rect 9338 7046 9348 7098
rect 9348 7046 9394 7098
rect 9098 7044 9154 7046
rect 9178 7044 9234 7046
rect 9258 7044 9314 7046
rect 9338 7044 9394 7046
rect 10966 10104 11022 10160
rect 11812 14170 11868 14172
rect 11892 14170 11948 14172
rect 11972 14170 12028 14172
rect 12052 14170 12108 14172
rect 11812 14118 11858 14170
rect 11858 14118 11868 14170
rect 11892 14118 11922 14170
rect 11922 14118 11934 14170
rect 11934 14118 11948 14170
rect 11972 14118 11986 14170
rect 11986 14118 11998 14170
rect 11998 14118 12028 14170
rect 12052 14118 12062 14170
rect 12062 14118 12108 14170
rect 11812 14116 11868 14118
rect 11892 14116 11948 14118
rect 11972 14116 12028 14118
rect 12052 14116 12108 14118
rect 11812 13082 11868 13084
rect 11892 13082 11948 13084
rect 11972 13082 12028 13084
rect 12052 13082 12108 13084
rect 11812 13030 11858 13082
rect 11858 13030 11868 13082
rect 11892 13030 11922 13082
rect 11922 13030 11934 13082
rect 11934 13030 11948 13082
rect 11972 13030 11986 13082
rect 11986 13030 11998 13082
rect 11998 13030 12028 13082
rect 12052 13030 12062 13082
rect 12062 13030 12108 13082
rect 11812 13028 11868 13030
rect 11892 13028 11948 13030
rect 11972 13028 12028 13030
rect 12052 13028 12108 13030
rect 11812 11994 11868 11996
rect 11892 11994 11948 11996
rect 11972 11994 12028 11996
rect 12052 11994 12108 11996
rect 11812 11942 11858 11994
rect 11858 11942 11868 11994
rect 11892 11942 11922 11994
rect 11922 11942 11934 11994
rect 11934 11942 11948 11994
rect 11972 11942 11986 11994
rect 11986 11942 11998 11994
rect 11998 11942 12028 11994
rect 12052 11942 12062 11994
rect 12062 11942 12108 11994
rect 11812 11940 11868 11942
rect 11892 11940 11948 11942
rect 11972 11940 12028 11942
rect 12052 11940 12108 11942
rect 11812 10906 11868 10908
rect 11892 10906 11948 10908
rect 11972 10906 12028 10908
rect 12052 10906 12108 10908
rect 11812 10854 11858 10906
rect 11858 10854 11868 10906
rect 11892 10854 11922 10906
rect 11922 10854 11934 10906
rect 11934 10854 11948 10906
rect 11972 10854 11986 10906
rect 11986 10854 11998 10906
rect 11998 10854 12028 10906
rect 12052 10854 12062 10906
rect 12062 10854 12108 10906
rect 11812 10852 11868 10854
rect 11892 10852 11948 10854
rect 11972 10852 12028 10854
rect 12052 10852 12108 10854
rect 11812 9818 11868 9820
rect 11892 9818 11948 9820
rect 11972 9818 12028 9820
rect 12052 9818 12108 9820
rect 11812 9766 11858 9818
rect 11858 9766 11868 9818
rect 11892 9766 11922 9818
rect 11922 9766 11934 9818
rect 11934 9766 11948 9818
rect 11972 9766 11986 9818
rect 11986 9766 11998 9818
rect 11998 9766 12028 9818
rect 12052 9766 12062 9818
rect 12062 9766 12108 9818
rect 11812 9764 11868 9766
rect 11892 9764 11948 9766
rect 11972 9764 12028 9766
rect 12052 9764 12108 9766
rect 11812 8730 11868 8732
rect 11892 8730 11948 8732
rect 11972 8730 12028 8732
rect 12052 8730 12108 8732
rect 11812 8678 11858 8730
rect 11858 8678 11868 8730
rect 11892 8678 11922 8730
rect 11922 8678 11934 8730
rect 11934 8678 11948 8730
rect 11972 8678 11986 8730
rect 11986 8678 11998 8730
rect 11998 8678 12028 8730
rect 12052 8678 12062 8730
rect 12062 8678 12108 8730
rect 11812 8676 11868 8678
rect 11892 8676 11948 8678
rect 11972 8676 12028 8678
rect 12052 8676 12108 8678
rect 11812 7642 11868 7644
rect 11892 7642 11948 7644
rect 11972 7642 12028 7644
rect 12052 7642 12108 7644
rect 11812 7590 11858 7642
rect 11858 7590 11868 7642
rect 11892 7590 11922 7642
rect 11922 7590 11934 7642
rect 11934 7590 11948 7642
rect 11972 7590 11986 7642
rect 11986 7590 11998 7642
rect 11998 7590 12028 7642
rect 12052 7590 12062 7642
rect 12062 7590 12108 7642
rect 11812 7588 11868 7590
rect 11892 7588 11948 7590
rect 11972 7588 12028 7590
rect 12052 7588 12108 7590
rect 11812 6554 11868 6556
rect 11892 6554 11948 6556
rect 11972 6554 12028 6556
rect 12052 6554 12108 6556
rect 11812 6502 11858 6554
rect 11858 6502 11868 6554
rect 11892 6502 11922 6554
rect 11922 6502 11934 6554
rect 11934 6502 11948 6554
rect 11972 6502 11986 6554
rect 11986 6502 11998 6554
rect 11998 6502 12028 6554
rect 12052 6502 12062 6554
rect 12062 6502 12108 6554
rect 11812 6500 11868 6502
rect 11892 6500 11948 6502
rect 11972 6500 12028 6502
rect 12052 6500 12108 6502
rect 6384 4378 6440 4380
rect 6464 4378 6520 4380
rect 6544 4378 6600 4380
rect 6624 4378 6680 4380
rect 6384 4326 6430 4378
rect 6430 4326 6440 4378
rect 6464 4326 6494 4378
rect 6494 4326 6506 4378
rect 6506 4326 6520 4378
rect 6544 4326 6558 4378
rect 6558 4326 6570 4378
rect 6570 4326 6600 4378
rect 6624 4326 6634 4378
rect 6634 4326 6680 4378
rect 6384 4324 6440 4326
rect 6464 4324 6520 4326
rect 6544 4324 6600 4326
rect 6624 4324 6680 4326
rect 6384 3290 6440 3292
rect 6464 3290 6520 3292
rect 6544 3290 6600 3292
rect 6624 3290 6680 3292
rect 6384 3238 6430 3290
rect 6430 3238 6440 3290
rect 6464 3238 6494 3290
rect 6494 3238 6506 3290
rect 6506 3238 6520 3290
rect 6544 3238 6558 3290
rect 6558 3238 6570 3290
rect 6570 3238 6600 3290
rect 6624 3238 6634 3290
rect 6634 3238 6680 3290
rect 6384 3236 6440 3238
rect 6464 3236 6520 3238
rect 6544 3236 6600 3238
rect 6624 3236 6680 3238
rect 9098 6010 9154 6012
rect 9178 6010 9234 6012
rect 9258 6010 9314 6012
rect 9338 6010 9394 6012
rect 9098 5958 9144 6010
rect 9144 5958 9154 6010
rect 9178 5958 9208 6010
rect 9208 5958 9220 6010
rect 9220 5958 9234 6010
rect 9258 5958 9272 6010
rect 9272 5958 9284 6010
rect 9284 5958 9314 6010
rect 9338 5958 9348 6010
rect 9348 5958 9394 6010
rect 9098 5956 9154 5958
rect 9178 5956 9234 5958
rect 9258 5956 9314 5958
rect 9338 5956 9394 5958
rect 11812 5466 11868 5468
rect 11892 5466 11948 5468
rect 11972 5466 12028 5468
rect 12052 5466 12108 5468
rect 11812 5414 11858 5466
rect 11858 5414 11868 5466
rect 11892 5414 11922 5466
rect 11922 5414 11934 5466
rect 11934 5414 11948 5466
rect 11972 5414 11986 5466
rect 11986 5414 11998 5466
rect 11998 5414 12028 5466
rect 12052 5414 12062 5466
rect 12062 5414 12108 5466
rect 11812 5412 11868 5414
rect 11892 5412 11948 5414
rect 11972 5412 12028 5414
rect 12052 5412 12108 5414
rect 9098 4922 9154 4924
rect 9178 4922 9234 4924
rect 9258 4922 9314 4924
rect 9338 4922 9394 4924
rect 9098 4870 9144 4922
rect 9144 4870 9154 4922
rect 9178 4870 9208 4922
rect 9208 4870 9220 4922
rect 9220 4870 9234 4922
rect 9258 4870 9272 4922
rect 9272 4870 9284 4922
rect 9284 4870 9314 4922
rect 9338 4870 9348 4922
rect 9348 4870 9394 4922
rect 9098 4868 9154 4870
rect 9178 4868 9234 4870
rect 9258 4868 9314 4870
rect 9338 4868 9394 4870
rect 11812 4378 11868 4380
rect 11892 4378 11948 4380
rect 11972 4378 12028 4380
rect 12052 4378 12108 4380
rect 11812 4326 11858 4378
rect 11858 4326 11868 4378
rect 11892 4326 11922 4378
rect 11922 4326 11934 4378
rect 11934 4326 11948 4378
rect 11972 4326 11986 4378
rect 11986 4326 11998 4378
rect 11998 4326 12028 4378
rect 12052 4326 12062 4378
rect 12062 4326 12108 4378
rect 11812 4324 11868 4326
rect 11892 4324 11948 4326
rect 11972 4324 12028 4326
rect 12052 4324 12108 4326
rect 14526 15802 14582 15804
rect 14606 15802 14662 15804
rect 14686 15802 14742 15804
rect 14766 15802 14822 15804
rect 14526 15750 14572 15802
rect 14572 15750 14582 15802
rect 14606 15750 14636 15802
rect 14636 15750 14648 15802
rect 14648 15750 14662 15802
rect 14686 15750 14700 15802
rect 14700 15750 14712 15802
rect 14712 15750 14742 15802
rect 14766 15750 14776 15802
rect 14776 15750 14822 15802
rect 14526 15748 14582 15750
rect 14606 15748 14662 15750
rect 14686 15748 14742 15750
rect 14766 15748 14822 15750
rect 19954 15802 20010 15804
rect 20034 15802 20090 15804
rect 20114 15802 20170 15804
rect 20194 15802 20250 15804
rect 19954 15750 20000 15802
rect 20000 15750 20010 15802
rect 20034 15750 20064 15802
rect 20064 15750 20076 15802
rect 20076 15750 20090 15802
rect 20114 15750 20128 15802
rect 20128 15750 20140 15802
rect 20140 15750 20170 15802
rect 20194 15750 20204 15802
rect 20204 15750 20250 15802
rect 19954 15748 20010 15750
rect 20034 15748 20090 15750
rect 20114 15748 20170 15750
rect 20194 15748 20250 15750
rect 17240 15258 17296 15260
rect 17320 15258 17376 15260
rect 17400 15258 17456 15260
rect 17480 15258 17536 15260
rect 17240 15206 17286 15258
rect 17286 15206 17296 15258
rect 17320 15206 17350 15258
rect 17350 15206 17362 15258
rect 17362 15206 17376 15258
rect 17400 15206 17414 15258
rect 17414 15206 17426 15258
rect 17426 15206 17456 15258
rect 17480 15206 17490 15258
rect 17490 15206 17536 15258
rect 17240 15204 17296 15206
rect 17320 15204 17376 15206
rect 17400 15204 17456 15206
rect 17480 15204 17536 15206
rect 22668 15258 22724 15260
rect 22748 15258 22804 15260
rect 22828 15258 22884 15260
rect 22908 15258 22964 15260
rect 22668 15206 22714 15258
rect 22714 15206 22724 15258
rect 22748 15206 22778 15258
rect 22778 15206 22790 15258
rect 22790 15206 22804 15258
rect 22828 15206 22842 15258
rect 22842 15206 22854 15258
rect 22854 15206 22884 15258
rect 22908 15206 22918 15258
rect 22918 15206 22964 15258
rect 22668 15204 22724 15206
rect 22748 15204 22804 15206
rect 22828 15204 22884 15206
rect 22908 15204 22964 15206
rect 14526 14714 14582 14716
rect 14606 14714 14662 14716
rect 14686 14714 14742 14716
rect 14766 14714 14822 14716
rect 14526 14662 14572 14714
rect 14572 14662 14582 14714
rect 14606 14662 14636 14714
rect 14636 14662 14648 14714
rect 14648 14662 14662 14714
rect 14686 14662 14700 14714
rect 14700 14662 14712 14714
rect 14712 14662 14742 14714
rect 14766 14662 14776 14714
rect 14776 14662 14822 14714
rect 14526 14660 14582 14662
rect 14606 14660 14662 14662
rect 14686 14660 14742 14662
rect 14766 14660 14822 14662
rect 19954 14714 20010 14716
rect 20034 14714 20090 14716
rect 20114 14714 20170 14716
rect 20194 14714 20250 14716
rect 19954 14662 20000 14714
rect 20000 14662 20010 14714
rect 20034 14662 20064 14714
rect 20064 14662 20076 14714
rect 20076 14662 20090 14714
rect 20114 14662 20128 14714
rect 20128 14662 20140 14714
rect 20140 14662 20170 14714
rect 20194 14662 20204 14714
rect 20204 14662 20250 14714
rect 19954 14660 20010 14662
rect 20034 14660 20090 14662
rect 20114 14660 20170 14662
rect 20194 14660 20250 14662
rect 17240 14170 17296 14172
rect 17320 14170 17376 14172
rect 17400 14170 17456 14172
rect 17480 14170 17536 14172
rect 17240 14118 17286 14170
rect 17286 14118 17296 14170
rect 17320 14118 17350 14170
rect 17350 14118 17362 14170
rect 17362 14118 17376 14170
rect 17400 14118 17414 14170
rect 17414 14118 17426 14170
rect 17426 14118 17456 14170
rect 17480 14118 17490 14170
rect 17490 14118 17536 14170
rect 17240 14116 17296 14118
rect 17320 14116 17376 14118
rect 17400 14116 17456 14118
rect 17480 14116 17536 14118
rect 22668 14170 22724 14172
rect 22748 14170 22804 14172
rect 22828 14170 22884 14172
rect 22908 14170 22964 14172
rect 22668 14118 22714 14170
rect 22714 14118 22724 14170
rect 22748 14118 22778 14170
rect 22778 14118 22790 14170
rect 22790 14118 22804 14170
rect 22828 14118 22842 14170
rect 22842 14118 22854 14170
rect 22854 14118 22884 14170
rect 22908 14118 22918 14170
rect 22918 14118 22964 14170
rect 22668 14116 22724 14118
rect 22748 14116 22804 14118
rect 22828 14116 22884 14118
rect 22908 14116 22964 14118
rect 14526 13626 14582 13628
rect 14606 13626 14662 13628
rect 14686 13626 14742 13628
rect 14766 13626 14822 13628
rect 14526 13574 14572 13626
rect 14572 13574 14582 13626
rect 14606 13574 14636 13626
rect 14636 13574 14648 13626
rect 14648 13574 14662 13626
rect 14686 13574 14700 13626
rect 14700 13574 14712 13626
rect 14712 13574 14742 13626
rect 14766 13574 14776 13626
rect 14776 13574 14822 13626
rect 14526 13572 14582 13574
rect 14606 13572 14662 13574
rect 14686 13572 14742 13574
rect 14766 13572 14822 13574
rect 12990 7404 13046 7440
rect 12990 7384 12992 7404
rect 12992 7384 13044 7404
rect 13044 7384 13046 7404
rect 9098 3834 9154 3836
rect 9178 3834 9234 3836
rect 9258 3834 9314 3836
rect 9338 3834 9394 3836
rect 9098 3782 9144 3834
rect 9144 3782 9154 3834
rect 9178 3782 9208 3834
rect 9208 3782 9220 3834
rect 9220 3782 9234 3834
rect 9258 3782 9272 3834
rect 9272 3782 9284 3834
rect 9284 3782 9314 3834
rect 9338 3782 9348 3834
rect 9348 3782 9394 3834
rect 9098 3780 9154 3782
rect 9178 3780 9234 3782
rect 9258 3780 9314 3782
rect 9338 3780 9394 3782
rect 9098 2746 9154 2748
rect 9178 2746 9234 2748
rect 9258 2746 9314 2748
rect 9338 2746 9394 2748
rect 9098 2694 9144 2746
rect 9144 2694 9154 2746
rect 9178 2694 9208 2746
rect 9208 2694 9220 2746
rect 9220 2694 9234 2746
rect 9258 2694 9272 2746
rect 9272 2694 9284 2746
rect 9284 2694 9314 2746
rect 9338 2694 9348 2746
rect 9348 2694 9394 2746
rect 9098 2692 9154 2694
rect 9178 2692 9234 2694
rect 9258 2692 9314 2694
rect 9338 2692 9394 2694
rect 10966 3460 11022 3496
rect 10966 3440 10968 3460
rect 10968 3440 11020 3460
rect 11020 3440 11022 3460
rect 13910 8372 13912 8392
rect 13912 8372 13964 8392
rect 13964 8372 13966 8392
rect 13910 8336 13966 8372
rect 14278 11212 14334 11248
rect 14278 11192 14280 11212
rect 14280 11192 14332 11212
rect 14332 11192 14334 11212
rect 13082 5072 13138 5128
rect 11812 3290 11868 3292
rect 11892 3290 11948 3292
rect 11972 3290 12028 3292
rect 12052 3290 12108 3292
rect 11812 3238 11858 3290
rect 11858 3238 11868 3290
rect 11892 3238 11922 3290
rect 11922 3238 11934 3290
rect 11934 3238 11948 3290
rect 11972 3238 11986 3290
rect 11986 3238 11998 3290
rect 11998 3238 12028 3290
rect 12052 3238 12062 3290
rect 12062 3238 12108 3290
rect 11812 3236 11868 3238
rect 11892 3236 11948 3238
rect 11972 3236 12028 3238
rect 12052 3236 12108 3238
rect 19954 13626 20010 13628
rect 20034 13626 20090 13628
rect 20114 13626 20170 13628
rect 20194 13626 20250 13628
rect 19954 13574 20000 13626
rect 20000 13574 20010 13626
rect 20034 13574 20064 13626
rect 20064 13574 20076 13626
rect 20076 13574 20090 13626
rect 20114 13574 20128 13626
rect 20128 13574 20140 13626
rect 20140 13574 20170 13626
rect 20194 13574 20204 13626
rect 20204 13574 20250 13626
rect 19954 13572 20010 13574
rect 20034 13572 20090 13574
rect 20114 13572 20170 13574
rect 20194 13572 20250 13574
rect 14526 12538 14582 12540
rect 14606 12538 14662 12540
rect 14686 12538 14742 12540
rect 14766 12538 14822 12540
rect 14526 12486 14572 12538
rect 14572 12486 14582 12538
rect 14606 12486 14636 12538
rect 14636 12486 14648 12538
rect 14648 12486 14662 12538
rect 14686 12486 14700 12538
rect 14700 12486 14712 12538
rect 14712 12486 14742 12538
rect 14766 12486 14776 12538
rect 14776 12486 14822 12538
rect 14526 12484 14582 12486
rect 14606 12484 14662 12486
rect 14686 12484 14742 12486
rect 14766 12484 14822 12486
rect 14526 11450 14582 11452
rect 14606 11450 14662 11452
rect 14686 11450 14742 11452
rect 14766 11450 14822 11452
rect 14526 11398 14572 11450
rect 14572 11398 14582 11450
rect 14606 11398 14636 11450
rect 14636 11398 14648 11450
rect 14648 11398 14662 11450
rect 14686 11398 14700 11450
rect 14700 11398 14712 11450
rect 14712 11398 14742 11450
rect 14766 11398 14776 11450
rect 14776 11398 14822 11450
rect 14526 11396 14582 11398
rect 14606 11396 14662 11398
rect 14686 11396 14742 11398
rect 14766 11396 14822 11398
rect 14526 10362 14582 10364
rect 14606 10362 14662 10364
rect 14686 10362 14742 10364
rect 14766 10362 14822 10364
rect 14526 10310 14572 10362
rect 14572 10310 14582 10362
rect 14606 10310 14636 10362
rect 14636 10310 14648 10362
rect 14648 10310 14662 10362
rect 14686 10310 14700 10362
rect 14700 10310 14712 10362
rect 14712 10310 14742 10362
rect 14766 10310 14776 10362
rect 14776 10310 14822 10362
rect 14526 10308 14582 10310
rect 14606 10308 14662 10310
rect 14686 10308 14742 10310
rect 14766 10308 14822 10310
rect 14526 9274 14582 9276
rect 14606 9274 14662 9276
rect 14686 9274 14742 9276
rect 14766 9274 14822 9276
rect 14526 9222 14572 9274
rect 14572 9222 14582 9274
rect 14606 9222 14636 9274
rect 14636 9222 14648 9274
rect 14648 9222 14662 9274
rect 14686 9222 14700 9274
rect 14700 9222 14712 9274
rect 14712 9222 14742 9274
rect 14766 9222 14776 9274
rect 14776 9222 14822 9274
rect 14526 9220 14582 9222
rect 14606 9220 14662 9222
rect 14686 9220 14742 9222
rect 14766 9220 14822 9222
rect 14526 8186 14582 8188
rect 14606 8186 14662 8188
rect 14686 8186 14742 8188
rect 14766 8186 14822 8188
rect 14526 8134 14572 8186
rect 14572 8134 14582 8186
rect 14606 8134 14636 8186
rect 14636 8134 14648 8186
rect 14648 8134 14662 8186
rect 14686 8134 14700 8186
rect 14700 8134 14712 8186
rect 14712 8134 14742 8186
rect 14766 8134 14776 8186
rect 14776 8134 14822 8186
rect 14526 8132 14582 8134
rect 14606 8132 14662 8134
rect 14686 8132 14742 8134
rect 14766 8132 14822 8134
rect 14526 7098 14582 7100
rect 14606 7098 14662 7100
rect 14686 7098 14742 7100
rect 14766 7098 14822 7100
rect 14526 7046 14572 7098
rect 14572 7046 14582 7098
rect 14606 7046 14636 7098
rect 14636 7046 14648 7098
rect 14648 7046 14662 7098
rect 14686 7046 14700 7098
rect 14700 7046 14712 7098
rect 14712 7046 14742 7098
rect 14766 7046 14776 7098
rect 14776 7046 14822 7098
rect 14526 7044 14582 7046
rect 14606 7044 14662 7046
rect 14686 7044 14742 7046
rect 14766 7044 14822 7046
rect 15290 11076 15346 11112
rect 15290 11056 15292 11076
rect 15292 11056 15344 11076
rect 15344 11056 15346 11076
rect 15750 8508 15752 8528
rect 15752 8508 15804 8528
rect 15804 8508 15806 8528
rect 15750 8472 15806 8508
rect 16394 11228 16396 11248
rect 16396 11228 16448 11248
rect 16448 11228 16450 11248
rect 16394 11192 16450 11228
rect 14526 6010 14582 6012
rect 14606 6010 14662 6012
rect 14686 6010 14742 6012
rect 14766 6010 14822 6012
rect 14526 5958 14572 6010
rect 14572 5958 14582 6010
rect 14606 5958 14636 6010
rect 14636 5958 14648 6010
rect 14648 5958 14662 6010
rect 14686 5958 14700 6010
rect 14700 5958 14712 6010
rect 14712 5958 14742 6010
rect 14766 5958 14776 6010
rect 14776 5958 14822 6010
rect 14526 5956 14582 5958
rect 14606 5956 14662 5958
rect 14686 5956 14742 5958
rect 14766 5956 14822 5958
rect 14738 5092 14794 5128
rect 14738 5072 14740 5092
rect 14740 5072 14792 5092
rect 14792 5072 14794 5092
rect 14526 4922 14582 4924
rect 14606 4922 14662 4924
rect 14686 4922 14742 4924
rect 14766 4922 14822 4924
rect 14526 4870 14572 4922
rect 14572 4870 14582 4922
rect 14606 4870 14636 4922
rect 14636 4870 14648 4922
rect 14648 4870 14662 4922
rect 14686 4870 14700 4922
rect 14700 4870 14712 4922
rect 14712 4870 14742 4922
rect 14766 4870 14776 4922
rect 14776 4870 14822 4922
rect 14526 4868 14582 4870
rect 14606 4868 14662 4870
rect 14686 4868 14742 4870
rect 14766 4868 14822 4870
rect 14526 3834 14582 3836
rect 14606 3834 14662 3836
rect 14686 3834 14742 3836
rect 14766 3834 14822 3836
rect 14526 3782 14572 3834
rect 14572 3782 14582 3834
rect 14606 3782 14636 3834
rect 14636 3782 14648 3834
rect 14648 3782 14662 3834
rect 14686 3782 14700 3834
rect 14700 3782 14712 3834
rect 14712 3782 14742 3834
rect 14766 3782 14776 3834
rect 14776 3782 14822 3834
rect 14526 3780 14582 3782
rect 14606 3780 14662 3782
rect 14686 3780 14742 3782
rect 14766 3780 14822 3782
rect 17240 13082 17296 13084
rect 17320 13082 17376 13084
rect 17400 13082 17456 13084
rect 17480 13082 17536 13084
rect 17240 13030 17286 13082
rect 17286 13030 17296 13082
rect 17320 13030 17350 13082
rect 17350 13030 17362 13082
rect 17362 13030 17376 13082
rect 17400 13030 17414 13082
rect 17414 13030 17426 13082
rect 17426 13030 17456 13082
rect 17480 13030 17490 13082
rect 17490 13030 17536 13082
rect 17240 13028 17296 13030
rect 17320 13028 17376 13030
rect 17400 13028 17456 13030
rect 17480 13028 17536 13030
rect 17240 11994 17296 11996
rect 17320 11994 17376 11996
rect 17400 11994 17456 11996
rect 17480 11994 17536 11996
rect 17240 11942 17286 11994
rect 17286 11942 17296 11994
rect 17320 11942 17350 11994
rect 17350 11942 17362 11994
rect 17362 11942 17376 11994
rect 17400 11942 17414 11994
rect 17414 11942 17426 11994
rect 17426 11942 17456 11994
rect 17480 11942 17490 11994
rect 17490 11942 17536 11994
rect 17240 11940 17296 11942
rect 17320 11940 17376 11942
rect 17400 11940 17456 11942
rect 17480 11940 17536 11942
rect 17240 10906 17296 10908
rect 17320 10906 17376 10908
rect 17400 10906 17456 10908
rect 17480 10906 17536 10908
rect 17240 10854 17286 10906
rect 17286 10854 17296 10906
rect 17320 10854 17350 10906
rect 17350 10854 17362 10906
rect 17362 10854 17376 10906
rect 17400 10854 17414 10906
rect 17414 10854 17426 10906
rect 17426 10854 17456 10906
rect 17480 10854 17490 10906
rect 17490 10854 17536 10906
rect 17240 10852 17296 10854
rect 17320 10852 17376 10854
rect 17400 10852 17456 10854
rect 17480 10852 17536 10854
rect 17682 10104 17738 10160
rect 17240 9818 17296 9820
rect 17320 9818 17376 9820
rect 17400 9818 17456 9820
rect 17480 9818 17536 9820
rect 17240 9766 17286 9818
rect 17286 9766 17296 9818
rect 17320 9766 17350 9818
rect 17350 9766 17362 9818
rect 17362 9766 17376 9818
rect 17400 9766 17414 9818
rect 17414 9766 17426 9818
rect 17426 9766 17456 9818
rect 17480 9766 17490 9818
rect 17490 9766 17536 9818
rect 17240 9764 17296 9766
rect 17320 9764 17376 9766
rect 17400 9764 17456 9766
rect 17480 9764 17536 9766
rect 17240 8730 17296 8732
rect 17320 8730 17376 8732
rect 17400 8730 17456 8732
rect 17480 8730 17536 8732
rect 17240 8678 17286 8730
rect 17286 8678 17296 8730
rect 17320 8678 17350 8730
rect 17350 8678 17362 8730
rect 17362 8678 17376 8730
rect 17400 8678 17414 8730
rect 17414 8678 17426 8730
rect 17426 8678 17456 8730
rect 17480 8678 17490 8730
rect 17490 8678 17536 8730
rect 17240 8676 17296 8678
rect 17320 8676 17376 8678
rect 17400 8676 17456 8678
rect 17480 8676 17536 8678
rect 17498 8336 17554 8392
rect 17240 7642 17296 7644
rect 17320 7642 17376 7644
rect 17400 7642 17456 7644
rect 17480 7642 17536 7644
rect 17240 7590 17286 7642
rect 17286 7590 17296 7642
rect 17320 7590 17350 7642
rect 17350 7590 17362 7642
rect 17362 7590 17376 7642
rect 17400 7590 17414 7642
rect 17414 7590 17426 7642
rect 17426 7590 17456 7642
rect 17480 7590 17490 7642
rect 17490 7590 17536 7642
rect 17240 7588 17296 7590
rect 17320 7588 17376 7590
rect 17400 7588 17456 7590
rect 17480 7588 17536 7590
rect 17240 6554 17296 6556
rect 17320 6554 17376 6556
rect 17400 6554 17456 6556
rect 17480 6554 17536 6556
rect 17240 6502 17286 6554
rect 17286 6502 17296 6554
rect 17320 6502 17350 6554
rect 17350 6502 17362 6554
rect 17362 6502 17376 6554
rect 17400 6502 17414 6554
rect 17414 6502 17426 6554
rect 17426 6502 17456 6554
rect 17480 6502 17490 6554
rect 17490 6502 17536 6554
rect 17240 6500 17296 6502
rect 17320 6500 17376 6502
rect 17400 6500 17456 6502
rect 17480 6500 17536 6502
rect 17240 5466 17296 5468
rect 17320 5466 17376 5468
rect 17400 5466 17456 5468
rect 17480 5466 17536 5468
rect 17240 5414 17286 5466
rect 17286 5414 17296 5466
rect 17320 5414 17350 5466
rect 17350 5414 17362 5466
rect 17362 5414 17376 5466
rect 17400 5414 17414 5466
rect 17414 5414 17426 5466
rect 17426 5414 17456 5466
rect 17480 5414 17490 5466
rect 17490 5414 17536 5466
rect 17240 5412 17296 5414
rect 17320 5412 17376 5414
rect 17400 5412 17456 5414
rect 17480 5412 17536 5414
rect 19954 12538 20010 12540
rect 20034 12538 20090 12540
rect 20114 12538 20170 12540
rect 20194 12538 20250 12540
rect 19954 12486 20000 12538
rect 20000 12486 20010 12538
rect 20034 12486 20064 12538
rect 20064 12486 20076 12538
rect 20076 12486 20090 12538
rect 20114 12486 20128 12538
rect 20128 12486 20140 12538
rect 20140 12486 20170 12538
rect 20194 12486 20204 12538
rect 20204 12486 20250 12538
rect 19954 12484 20010 12486
rect 20034 12484 20090 12486
rect 20114 12484 20170 12486
rect 20194 12484 20250 12486
rect 17866 8336 17922 8392
rect 19154 8492 19210 8528
rect 19154 8472 19156 8492
rect 19156 8472 19208 8492
rect 19208 8472 19210 8492
rect 22668 13082 22724 13084
rect 22748 13082 22804 13084
rect 22828 13082 22884 13084
rect 22908 13082 22964 13084
rect 22668 13030 22714 13082
rect 22714 13030 22724 13082
rect 22748 13030 22778 13082
rect 22778 13030 22790 13082
rect 22790 13030 22804 13082
rect 22828 13030 22842 13082
rect 22842 13030 22854 13082
rect 22854 13030 22884 13082
rect 22908 13030 22918 13082
rect 22918 13030 22964 13082
rect 22668 13028 22724 13030
rect 22748 13028 22804 13030
rect 22828 13028 22884 13030
rect 22908 13028 22964 13030
rect 19954 11450 20010 11452
rect 20034 11450 20090 11452
rect 20114 11450 20170 11452
rect 20194 11450 20250 11452
rect 19954 11398 20000 11450
rect 20000 11398 20010 11450
rect 20034 11398 20064 11450
rect 20064 11398 20076 11450
rect 20076 11398 20090 11450
rect 20114 11398 20128 11450
rect 20128 11398 20140 11450
rect 20140 11398 20170 11450
rect 20194 11398 20204 11450
rect 20204 11398 20250 11450
rect 19954 11396 20010 11398
rect 20034 11396 20090 11398
rect 20114 11396 20170 11398
rect 20194 11396 20250 11398
rect 19954 10362 20010 10364
rect 20034 10362 20090 10364
rect 20114 10362 20170 10364
rect 20194 10362 20250 10364
rect 19954 10310 20000 10362
rect 20000 10310 20010 10362
rect 20034 10310 20064 10362
rect 20064 10310 20076 10362
rect 20076 10310 20090 10362
rect 20114 10310 20128 10362
rect 20128 10310 20140 10362
rect 20140 10310 20170 10362
rect 20194 10310 20204 10362
rect 20204 10310 20250 10362
rect 19954 10308 20010 10310
rect 20034 10308 20090 10310
rect 20114 10308 20170 10310
rect 20194 10308 20250 10310
rect 17240 4378 17296 4380
rect 17320 4378 17376 4380
rect 17400 4378 17456 4380
rect 17480 4378 17536 4380
rect 17240 4326 17286 4378
rect 17286 4326 17296 4378
rect 17320 4326 17350 4378
rect 17350 4326 17362 4378
rect 17362 4326 17376 4378
rect 17400 4326 17414 4378
rect 17414 4326 17426 4378
rect 17426 4326 17456 4378
rect 17480 4326 17490 4378
rect 17490 4326 17536 4378
rect 17240 4324 17296 4326
rect 17320 4324 17376 4326
rect 17400 4324 17456 4326
rect 17480 4324 17536 4326
rect 19954 9274 20010 9276
rect 20034 9274 20090 9276
rect 20114 9274 20170 9276
rect 20194 9274 20250 9276
rect 19954 9222 20000 9274
rect 20000 9222 20010 9274
rect 20034 9222 20064 9274
rect 20064 9222 20076 9274
rect 20076 9222 20090 9274
rect 20114 9222 20128 9274
rect 20128 9222 20140 9274
rect 20140 9222 20170 9274
rect 20194 9222 20204 9274
rect 20204 9222 20250 9274
rect 19954 9220 20010 9222
rect 20034 9220 20090 9222
rect 20114 9220 20170 9222
rect 20194 9220 20250 9222
rect 19954 8186 20010 8188
rect 20034 8186 20090 8188
rect 20114 8186 20170 8188
rect 20194 8186 20250 8188
rect 19954 8134 20000 8186
rect 20000 8134 20010 8186
rect 20034 8134 20064 8186
rect 20064 8134 20076 8186
rect 20076 8134 20090 8186
rect 20114 8134 20128 8186
rect 20128 8134 20140 8186
rect 20140 8134 20170 8186
rect 20194 8134 20204 8186
rect 20204 8134 20250 8186
rect 19954 8132 20010 8134
rect 20034 8132 20090 8134
rect 20114 8132 20170 8134
rect 20194 8132 20250 8134
rect 19954 7098 20010 7100
rect 20034 7098 20090 7100
rect 20114 7098 20170 7100
rect 20194 7098 20250 7100
rect 19954 7046 20000 7098
rect 20000 7046 20010 7098
rect 20034 7046 20064 7098
rect 20064 7046 20076 7098
rect 20076 7046 20090 7098
rect 20114 7046 20128 7098
rect 20128 7046 20140 7098
rect 20140 7046 20170 7098
rect 20194 7046 20204 7098
rect 20204 7046 20250 7098
rect 19954 7044 20010 7046
rect 20034 7044 20090 7046
rect 20114 7044 20170 7046
rect 20194 7044 20250 7046
rect 22668 11994 22724 11996
rect 22748 11994 22804 11996
rect 22828 11994 22884 11996
rect 22908 11994 22964 11996
rect 22668 11942 22714 11994
rect 22714 11942 22724 11994
rect 22748 11942 22778 11994
rect 22778 11942 22790 11994
rect 22790 11942 22804 11994
rect 22828 11942 22842 11994
rect 22842 11942 22854 11994
rect 22854 11942 22884 11994
rect 22908 11942 22918 11994
rect 22918 11942 22964 11994
rect 22668 11940 22724 11942
rect 22748 11940 22804 11942
rect 22828 11940 22884 11942
rect 22908 11940 22964 11942
rect 22668 10906 22724 10908
rect 22748 10906 22804 10908
rect 22828 10906 22884 10908
rect 22908 10906 22964 10908
rect 22668 10854 22714 10906
rect 22714 10854 22724 10906
rect 22748 10854 22778 10906
rect 22778 10854 22790 10906
rect 22790 10854 22804 10906
rect 22828 10854 22842 10906
rect 22842 10854 22854 10906
rect 22854 10854 22884 10906
rect 22908 10854 22918 10906
rect 22918 10854 22964 10906
rect 22668 10852 22724 10854
rect 22748 10852 22804 10854
rect 22828 10852 22884 10854
rect 22908 10852 22964 10854
rect 22668 9818 22724 9820
rect 22748 9818 22804 9820
rect 22828 9818 22884 9820
rect 22908 9818 22964 9820
rect 22668 9766 22714 9818
rect 22714 9766 22724 9818
rect 22748 9766 22778 9818
rect 22778 9766 22790 9818
rect 22790 9766 22804 9818
rect 22828 9766 22842 9818
rect 22842 9766 22854 9818
rect 22854 9766 22884 9818
rect 22908 9766 22918 9818
rect 22918 9766 22964 9818
rect 22668 9764 22724 9766
rect 22748 9764 22804 9766
rect 22828 9764 22884 9766
rect 22908 9764 22964 9766
rect 22668 8730 22724 8732
rect 22748 8730 22804 8732
rect 22828 8730 22884 8732
rect 22908 8730 22964 8732
rect 22668 8678 22714 8730
rect 22714 8678 22724 8730
rect 22748 8678 22778 8730
rect 22778 8678 22790 8730
rect 22790 8678 22804 8730
rect 22828 8678 22842 8730
rect 22842 8678 22854 8730
rect 22854 8678 22884 8730
rect 22908 8678 22918 8730
rect 22918 8678 22964 8730
rect 22668 8676 22724 8678
rect 22748 8676 22804 8678
rect 22828 8676 22884 8678
rect 22908 8676 22964 8678
rect 22668 7642 22724 7644
rect 22748 7642 22804 7644
rect 22828 7642 22884 7644
rect 22908 7642 22964 7644
rect 22668 7590 22714 7642
rect 22714 7590 22724 7642
rect 22748 7590 22778 7642
rect 22778 7590 22790 7642
rect 22790 7590 22804 7642
rect 22828 7590 22842 7642
rect 22842 7590 22854 7642
rect 22854 7590 22884 7642
rect 22908 7590 22918 7642
rect 22918 7590 22964 7642
rect 22668 7588 22724 7590
rect 22748 7588 22804 7590
rect 22828 7588 22884 7590
rect 22908 7588 22964 7590
rect 22668 6554 22724 6556
rect 22748 6554 22804 6556
rect 22828 6554 22884 6556
rect 22908 6554 22964 6556
rect 22668 6502 22714 6554
rect 22714 6502 22724 6554
rect 22748 6502 22778 6554
rect 22778 6502 22790 6554
rect 22790 6502 22804 6554
rect 22828 6502 22842 6554
rect 22842 6502 22854 6554
rect 22854 6502 22884 6554
rect 22908 6502 22918 6554
rect 22918 6502 22964 6554
rect 22668 6500 22724 6502
rect 22748 6500 22804 6502
rect 22828 6500 22884 6502
rect 22908 6500 22964 6502
rect 19954 6010 20010 6012
rect 20034 6010 20090 6012
rect 20114 6010 20170 6012
rect 20194 6010 20250 6012
rect 19954 5958 20000 6010
rect 20000 5958 20010 6010
rect 20034 5958 20064 6010
rect 20064 5958 20076 6010
rect 20076 5958 20090 6010
rect 20114 5958 20128 6010
rect 20128 5958 20140 6010
rect 20140 5958 20170 6010
rect 20194 5958 20204 6010
rect 20204 5958 20250 6010
rect 19954 5956 20010 5958
rect 20034 5956 20090 5958
rect 20114 5956 20170 5958
rect 20194 5956 20250 5958
rect 22668 5466 22724 5468
rect 22748 5466 22804 5468
rect 22828 5466 22884 5468
rect 22908 5466 22964 5468
rect 22668 5414 22714 5466
rect 22714 5414 22724 5466
rect 22748 5414 22778 5466
rect 22778 5414 22790 5466
rect 22790 5414 22804 5466
rect 22828 5414 22842 5466
rect 22842 5414 22854 5466
rect 22854 5414 22884 5466
rect 22908 5414 22918 5466
rect 22918 5414 22964 5466
rect 22668 5412 22724 5414
rect 22748 5412 22804 5414
rect 22828 5412 22884 5414
rect 22908 5412 22964 5414
rect 19954 4922 20010 4924
rect 20034 4922 20090 4924
rect 20114 4922 20170 4924
rect 20194 4922 20250 4924
rect 19954 4870 20000 4922
rect 20000 4870 20010 4922
rect 20034 4870 20064 4922
rect 20064 4870 20076 4922
rect 20076 4870 20090 4922
rect 20114 4870 20128 4922
rect 20128 4870 20140 4922
rect 20140 4870 20170 4922
rect 20194 4870 20204 4922
rect 20204 4870 20250 4922
rect 19954 4868 20010 4870
rect 20034 4868 20090 4870
rect 20114 4868 20170 4870
rect 20194 4868 20250 4870
rect 22668 4378 22724 4380
rect 22748 4378 22804 4380
rect 22828 4378 22884 4380
rect 22908 4378 22964 4380
rect 22668 4326 22714 4378
rect 22714 4326 22724 4378
rect 22748 4326 22778 4378
rect 22778 4326 22790 4378
rect 22790 4326 22804 4378
rect 22828 4326 22842 4378
rect 22842 4326 22854 4378
rect 22854 4326 22884 4378
rect 22908 4326 22918 4378
rect 22918 4326 22964 4378
rect 22668 4324 22724 4326
rect 22748 4324 22804 4326
rect 22828 4324 22884 4326
rect 22908 4324 22964 4326
rect 19954 3834 20010 3836
rect 20034 3834 20090 3836
rect 20114 3834 20170 3836
rect 20194 3834 20250 3836
rect 19954 3782 20000 3834
rect 20000 3782 20010 3834
rect 20034 3782 20064 3834
rect 20064 3782 20076 3834
rect 20076 3782 20090 3834
rect 20114 3782 20128 3834
rect 20128 3782 20140 3834
rect 20140 3782 20170 3834
rect 20194 3782 20204 3834
rect 20204 3782 20250 3834
rect 19954 3780 20010 3782
rect 20034 3780 20090 3782
rect 20114 3780 20170 3782
rect 20194 3780 20250 3782
rect 19430 3440 19486 3496
rect 17240 3290 17296 3292
rect 17320 3290 17376 3292
rect 17400 3290 17456 3292
rect 17480 3290 17536 3292
rect 17240 3238 17286 3290
rect 17286 3238 17296 3290
rect 17320 3238 17350 3290
rect 17350 3238 17362 3290
rect 17362 3238 17376 3290
rect 17400 3238 17414 3290
rect 17414 3238 17426 3290
rect 17426 3238 17456 3290
rect 17480 3238 17490 3290
rect 17490 3238 17536 3290
rect 17240 3236 17296 3238
rect 17320 3236 17376 3238
rect 17400 3236 17456 3238
rect 17480 3236 17536 3238
rect 22668 3290 22724 3292
rect 22748 3290 22804 3292
rect 22828 3290 22884 3292
rect 22908 3290 22964 3292
rect 22668 3238 22714 3290
rect 22714 3238 22724 3290
rect 22748 3238 22778 3290
rect 22778 3238 22790 3290
rect 22790 3238 22804 3290
rect 22828 3238 22842 3290
rect 22842 3238 22854 3290
rect 22854 3238 22884 3290
rect 22908 3238 22918 3290
rect 22918 3238 22964 3290
rect 22668 3236 22724 3238
rect 22748 3236 22804 3238
rect 22828 3236 22884 3238
rect 22908 3236 22964 3238
rect 14526 2746 14582 2748
rect 14606 2746 14662 2748
rect 14686 2746 14742 2748
rect 14766 2746 14822 2748
rect 14526 2694 14572 2746
rect 14572 2694 14582 2746
rect 14606 2694 14636 2746
rect 14636 2694 14648 2746
rect 14648 2694 14662 2746
rect 14686 2694 14700 2746
rect 14700 2694 14712 2746
rect 14712 2694 14742 2746
rect 14766 2694 14776 2746
rect 14776 2694 14822 2746
rect 14526 2692 14582 2694
rect 14606 2692 14662 2694
rect 14686 2692 14742 2694
rect 14766 2692 14822 2694
rect 19954 2746 20010 2748
rect 20034 2746 20090 2748
rect 20114 2746 20170 2748
rect 20194 2746 20250 2748
rect 19954 2694 20000 2746
rect 20000 2694 20010 2746
rect 20034 2694 20064 2746
rect 20064 2694 20076 2746
rect 20076 2694 20090 2746
rect 20114 2694 20128 2746
rect 20128 2694 20140 2746
rect 20140 2694 20170 2746
rect 20194 2694 20204 2746
rect 20204 2694 20250 2746
rect 19954 2692 20010 2694
rect 20034 2692 20090 2694
rect 20114 2692 20170 2694
rect 20194 2692 20250 2694
rect 6384 2202 6440 2204
rect 6464 2202 6520 2204
rect 6544 2202 6600 2204
rect 6624 2202 6680 2204
rect 6384 2150 6430 2202
rect 6430 2150 6440 2202
rect 6464 2150 6494 2202
rect 6494 2150 6506 2202
rect 6506 2150 6520 2202
rect 6544 2150 6558 2202
rect 6558 2150 6570 2202
rect 6570 2150 6600 2202
rect 6624 2150 6634 2202
rect 6634 2150 6680 2202
rect 6384 2148 6440 2150
rect 6464 2148 6520 2150
rect 6544 2148 6600 2150
rect 6624 2148 6680 2150
rect 11812 2202 11868 2204
rect 11892 2202 11948 2204
rect 11972 2202 12028 2204
rect 12052 2202 12108 2204
rect 11812 2150 11858 2202
rect 11858 2150 11868 2202
rect 11892 2150 11922 2202
rect 11922 2150 11934 2202
rect 11934 2150 11948 2202
rect 11972 2150 11986 2202
rect 11986 2150 11998 2202
rect 11998 2150 12028 2202
rect 12052 2150 12062 2202
rect 12062 2150 12108 2202
rect 11812 2148 11868 2150
rect 11892 2148 11948 2150
rect 11972 2148 12028 2150
rect 12052 2148 12108 2150
rect 17240 2202 17296 2204
rect 17320 2202 17376 2204
rect 17400 2202 17456 2204
rect 17480 2202 17536 2204
rect 17240 2150 17286 2202
rect 17286 2150 17296 2202
rect 17320 2150 17350 2202
rect 17350 2150 17362 2202
rect 17362 2150 17376 2202
rect 17400 2150 17414 2202
rect 17414 2150 17426 2202
rect 17426 2150 17456 2202
rect 17480 2150 17490 2202
rect 17490 2150 17536 2202
rect 17240 2148 17296 2150
rect 17320 2148 17376 2150
rect 17400 2148 17456 2150
rect 17480 2148 17536 2150
rect 22668 2202 22724 2204
rect 22748 2202 22804 2204
rect 22828 2202 22884 2204
rect 22908 2202 22964 2204
rect 22668 2150 22714 2202
rect 22714 2150 22724 2202
rect 22748 2150 22778 2202
rect 22778 2150 22790 2202
rect 22790 2150 22804 2202
rect 22828 2150 22842 2202
rect 22842 2150 22854 2202
rect 22854 2150 22884 2202
rect 22908 2150 22918 2202
rect 22918 2150 22964 2202
rect 22668 2148 22724 2150
rect 22748 2148 22804 2150
rect 22828 2148 22884 2150
rect 22908 2148 22964 2150
<< metal3 >>
rect 6374 21792 6690 21793
rect 6374 21728 6380 21792
rect 6444 21728 6460 21792
rect 6524 21728 6540 21792
rect 6604 21728 6620 21792
rect 6684 21728 6690 21792
rect 6374 21727 6690 21728
rect 11802 21792 12118 21793
rect 11802 21728 11808 21792
rect 11872 21728 11888 21792
rect 11952 21728 11968 21792
rect 12032 21728 12048 21792
rect 12112 21728 12118 21792
rect 11802 21727 12118 21728
rect 17230 21792 17546 21793
rect 17230 21728 17236 21792
rect 17300 21728 17316 21792
rect 17380 21728 17396 21792
rect 17460 21728 17476 21792
rect 17540 21728 17546 21792
rect 17230 21727 17546 21728
rect 22658 21792 22974 21793
rect 22658 21728 22664 21792
rect 22728 21728 22744 21792
rect 22808 21728 22824 21792
rect 22888 21728 22904 21792
rect 22968 21728 22974 21792
rect 22658 21727 22974 21728
rect 3660 21248 3976 21249
rect 3660 21184 3666 21248
rect 3730 21184 3746 21248
rect 3810 21184 3826 21248
rect 3890 21184 3906 21248
rect 3970 21184 3976 21248
rect 3660 21183 3976 21184
rect 9088 21248 9404 21249
rect 9088 21184 9094 21248
rect 9158 21184 9174 21248
rect 9238 21184 9254 21248
rect 9318 21184 9334 21248
rect 9398 21184 9404 21248
rect 9088 21183 9404 21184
rect 14516 21248 14832 21249
rect 14516 21184 14522 21248
rect 14586 21184 14602 21248
rect 14666 21184 14682 21248
rect 14746 21184 14762 21248
rect 14826 21184 14832 21248
rect 14516 21183 14832 21184
rect 19944 21248 20260 21249
rect 19944 21184 19950 21248
rect 20014 21184 20030 21248
rect 20094 21184 20110 21248
rect 20174 21184 20190 21248
rect 20254 21184 20260 21248
rect 19944 21183 20260 21184
rect 6374 20704 6690 20705
rect 6374 20640 6380 20704
rect 6444 20640 6460 20704
rect 6524 20640 6540 20704
rect 6604 20640 6620 20704
rect 6684 20640 6690 20704
rect 6374 20639 6690 20640
rect 11802 20704 12118 20705
rect 11802 20640 11808 20704
rect 11872 20640 11888 20704
rect 11952 20640 11968 20704
rect 12032 20640 12048 20704
rect 12112 20640 12118 20704
rect 11802 20639 12118 20640
rect 17230 20704 17546 20705
rect 17230 20640 17236 20704
rect 17300 20640 17316 20704
rect 17380 20640 17396 20704
rect 17460 20640 17476 20704
rect 17540 20640 17546 20704
rect 17230 20639 17546 20640
rect 22658 20704 22974 20705
rect 22658 20640 22664 20704
rect 22728 20640 22744 20704
rect 22808 20640 22824 20704
rect 22888 20640 22904 20704
rect 22968 20640 22974 20704
rect 22658 20639 22974 20640
rect 3660 20160 3976 20161
rect 3660 20096 3666 20160
rect 3730 20096 3746 20160
rect 3810 20096 3826 20160
rect 3890 20096 3906 20160
rect 3970 20096 3976 20160
rect 3660 20095 3976 20096
rect 9088 20160 9404 20161
rect 9088 20096 9094 20160
rect 9158 20096 9174 20160
rect 9238 20096 9254 20160
rect 9318 20096 9334 20160
rect 9398 20096 9404 20160
rect 9088 20095 9404 20096
rect 14516 20160 14832 20161
rect 14516 20096 14522 20160
rect 14586 20096 14602 20160
rect 14666 20096 14682 20160
rect 14746 20096 14762 20160
rect 14826 20096 14832 20160
rect 14516 20095 14832 20096
rect 19944 20160 20260 20161
rect 19944 20096 19950 20160
rect 20014 20096 20030 20160
rect 20094 20096 20110 20160
rect 20174 20096 20190 20160
rect 20254 20096 20260 20160
rect 19944 20095 20260 20096
rect 0 19818 800 19848
rect 933 19818 999 19821
rect 0 19816 999 19818
rect 0 19760 938 19816
rect 994 19760 999 19816
rect 0 19758 999 19760
rect 0 19728 800 19758
rect 933 19755 999 19758
rect 6374 19616 6690 19617
rect 6374 19552 6380 19616
rect 6444 19552 6460 19616
rect 6524 19552 6540 19616
rect 6604 19552 6620 19616
rect 6684 19552 6690 19616
rect 6374 19551 6690 19552
rect 11802 19616 12118 19617
rect 11802 19552 11808 19616
rect 11872 19552 11888 19616
rect 11952 19552 11968 19616
rect 12032 19552 12048 19616
rect 12112 19552 12118 19616
rect 11802 19551 12118 19552
rect 17230 19616 17546 19617
rect 17230 19552 17236 19616
rect 17300 19552 17316 19616
rect 17380 19552 17396 19616
rect 17460 19552 17476 19616
rect 17540 19552 17546 19616
rect 17230 19551 17546 19552
rect 22658 19616 22974 19617
rect 22658 19552 22664 19616
rect 22728 19552 22744 19616
rect 22808 19552 22824 19616
rect 22888 19552 22904 19616
rect 22968 19552 22974 19616
rect 22658 19551 22974 19552
rect 3660 19072 3976 19073
rect 3660 19008 3666 19072
rect 3730 19008 3746 19072
rect 3810 19008 3826 19072
rect 3890 19008 3906 19072
rect 3970 19008 3976 19072
rect 3660 19007 3976 19008
rect 9088 19072 9404 19073
rect 9088 19008 9094 19072
rect 9158 19008 9174 19072
rect 9238 19008 9254 19072
rect 9318 19008 9334 19072
rect 9398 19008 9404 19072
rect 9088 19007 9404 19008
rect 14516 19072 14832 19073
rect 14516 19008 14522 19072
rect 14586 19008 14602 19072
rect 14666 19008 14682 19072
rect 14746 19008 14762 19072
rect 14826 19008 14832 19072
rect 14516 19007 14832 19008
rect 19944 19072 20260 19073
rect 19944 19008 19950 19072
rect 20014 19008 20030 19072
rect 20094 19008 20110 19072
rect 20174 19008 20190 19072
rect 20254 19008 20260 19072
rect 19944 19007 20260 19008
rect 6374 18528 6690 18529
rect 6374 18464 6380 18528
rect 6444 18464 6460 18528
rect 6524 18464 6540 18528
rect 6604 18464 6620 18528
rect 6684 18464 6690 18528
rect 6374 18463 6690 18464
rect 11802 18528 12118 18529
rect 11802 18464 11808 18528
rect 11872 18464 11888 18528
rect 11952 18464 11968 18528
rect 12032 18464 12048 18528
rect 12112 18464 12118 18528
rect 11802 18463 12118 18464
rect 17230 18528 17546 18529
rect 17230 18464 17236 18528
rect 17300 18464 17316 18528
rect 17380 18464 17396 18528
rect 17460 18464 17476 18528
rect 17540 18464 17546 18528
rect 17230 18463 17546 18464
rect 22658 18528 22974 18529
rect 22658 18464 22664 18528
rect 22728 18464 22744 18528
rect 22808 18464 22824 18528
rect 22888 18464 22904 18528
rect 22968 18464 22974 18528
rect 22658 18463 22974 18464
rect 3660 17984 3976 17985
rect 3660 17920 3666 17984
rect 3730 17920 3746 17984
rect 3810 17920 3826 17984
rect 3890 17920 3906 17984
rect 3970 17920 3976 17984
rect 3660 17919 3976 17920
rect 9088 17984 9404 17985
rect 9088 17920 9094 17984
rect 9158 17920 9174 17984
rect 9238 17920 9254 17984
rect 9318 17920 9334 17984
rect 9398 17920 9404 17984
rect 9088 17919 9404 17920
rect 14516 17984 14832 17985
rect 14516 17920 14522 17984
rect 14586 17920 14602 17984
rect 14666 17920 14682 17984
rect 14746 17920 14762 17984
rect 14826 17920 14832 17984
rect 14516 17919 14832 17920
rect 19944 17984 20260 17985
rect 19944 17920 19950 17984
rect 20014 17920 20030 17984
rect 20094 17920 20110 17984
rect 20174 17920 20190 17984
rect 20254 17920 20260 17984
rect 19944 17919 20260 17920
rect 6374 17440 6690 17441
rect 6374 17376 6380 17440
rect 6444 17376 6460 17440
rect 6524 17376 6540 17440
rect 6604 17376 6620 17440
rect 6684 17376 6690 17440
rect 6374 17375 6690 17376
rect 11802 17440 12118 17441
rect 11802 17376 11808 17440
rect 11872 17376 11888 17440
rect 11952 17376 11968 17440
rect 12032 17376 12048 17440
rect 12112 17376 12118 17440
rect 11802 17375 12118 17376
rect 17230 17440 17546 17441
rect 17230 17376 17236 17440
rect 17300 17376 17316 17440
rect 17380 17376 17396 17440
rect 17460 17376 17476 17440
rect 17540 17376 17546 17440
rect 17230 17375 17546 17376
rect 22658 17440 22974 17441
rect 22658 17376 22664 17440
rect 22728 17376 22744 17440
rect 22808 17376 22824 17440
rect 22888 17376 22904 17440
rect 22968 17376 22974 17440
rect 22658 17375 22974 17376
rect 3660 16896 3976 16897
rect 3660 16832 3666 16896
rect 3730 16832 3746 16896
rect 3810 16832 3826 16896
rect 3890 16832 3906 16896
rect 3970 16832 3976 16896
rect 3660 16831 3976 16832
rect 9088 16896 9404 16897
rect 9088 16832 9094 16896
rect 9158 16832 9174 16896
rect 9238 16832 9254 16896
rect 9318 16832 9334 16896
rect 9398 16832 9404 16896
rect 9088 16831 9404 16832
rect 14516 16896 14832 16897
rect 14516 16832 14522 16896
rect 14586 16832 14602 16896
rect 14666 16832 14682 16896
rect 14746 16832 14762 16896
rect 14826 16832 14832 16896
rect 14516 16831 14832 16832
rect 19944 16896 20260 16897
rect 19944 16832 19950 16896
rect 20014 16832 20030 16896
rect 20094 16832 20110 16896
rect 20174 16832 20190 16896
rect 20254 16832 20260 16896
rect 19944 16831 20260 16832
rect 6374 16352 6690 16353
rect 6374 16288 6380 16352
rect 6444 16288 6460 16352
rect 6524 16288 6540 16352
rect 6604 16288 6620 16352
rect 6684 16288 6690 16352
rect 6374 16287 6690 16288
rect 11802 16352 12118 16353
rect 11802 16288 11808 16352
rect 11872 16288 11888 16352
rect 11952 16288 11968 16352
rect 12032 16288 12048 16352
rect 12112 16288 12118 16352
rect 11802 16287 12118 16288
rect 17230 16352 17546 16353
rect 17230 16288 17236 16352
rect 17300 16288 17316 16352
rect 17380 16288 17396 16352
rect 17460 16288 17476 16352
rect 17540 16288 17546 16352
rect 17230 16287 17546 16288
rect 22658 16352 22974 16353
rect 22658 16288 22664 16352
rect 22728 16288 22744 16352
rect 22808 16288 22824 16352
rect 22888 16288 22904 16352
rect 22968 16288 22974 16352
rect 22658 16287 22974 16288
rect 3660 15808 3976 15809
rect 3660 15744 3666 15808
rect 3730 15744 3746 15808
rect 3810 15744 3826 15808
rect 3890 15744 3906 15808
rect 3970 15744 3976 15808
rect 3660 15743 3976 15744
rect 9088 15808 9404 15809
rect 9088 15744 9094 15808
rect 9158 15744 9174 15808
rect 9238 15744 9254 15808
rect 9318 15744 9334 15808
rect 9398 15744 9404 15808
rect 9088 15743 9404 15744
rect 14516 15808 14832 15809
rect 14516 15744 14522 15808
rect 14586 15744 14602 15808
rect 14666 15744 14682 15808
rect 14746 15744 14762 15808
rect 14826 15744 14832 15808
rect 14516 15743 14832 15744
rect 19944 15808 20260 15809
rect 19944 15744 19950 15808
rect 20014 15744 20030 15808
rect 20094 15744 20110 15808
rect 20174 15744 20190 15808
rect 20254 15744 20260 15808
rect 19944 15743 20260 15744
rect 6374 15264 6690 15265
rect 6374 15200 6380 15264
rect 6444 15200 6460 15264
rect 6524 15200 6540 15264
rect 6604 15200 6620 15264
rect 6684 15200 6690 15264
rect 6374 15199 6690 15200
rect 11802 15264 12118 15265
rect 11802 15200 11808 15264
rect 11872 15200 11888 15264
rect 11952 15200 11968 15264
rect 12032 15200 12048 15264
rect 12112 15200 12118 15264
rect 11802 15199 12118 15200
rect 17230 15264 17546 15265
rect 17230 15200 17236 15264
rect 17300 15200 17316 15264
rect 17380 15200 17396 15264
rect 17460 15200 17476 15264
rect 17540 15200 17546 15264
rect 17230 15199 17546 15200
rect 22658 15264 22974 15265
rect 22658 15200 22664 15264
rect 22728 15200 22744 15264
rect 22808 15200 22824 15264
rect 22888 15200 22904 15264
rect 22968 15200 22974 15264
rect 22658 15199 22974 15200
rect 3660 14720 3976 14721
rect 3660 14656 3666 14720
rect 3730 14656 3746 14720
rect 3810 14656 3826 14720
rect 3890 14656 3906 14720
rect 3970 14656 3976 14720
rect 3660 14655 3976 14656
rect 9088 14720 9404 14721
rect 9088 14656 9094 14720
rect 9158 14656 9174 14720
rect 9238 14656 9254 14720
rect 9318 14656 9334 14720
rect 9398 14656 9404 14720
rect 9088 14655 9404 14656
rect 14516 14720 14832 14721
rect 14516 14656 14522 14720
rect 14586 14656 14602 14720
rect 14666 14656 14682 14720
rect 14746 14656 14762 14720
rect 14826 14656 14832 14720
rect 14516 14655 14832 14656
rect 19944 14720 20260 14721
rect 19944 14656 19950 14720
rect 20014 14656 20030 14720
rect 20094 14656 20110 14720
rect 20174 14656 20190 14720
rect 20254 14656 20260 14720
rect 19944 14655 20260 14656
rect 6374 14176 6690 14177
rect 6374 14112 6380 14176
rect 6444 14112 6460 14176
rect 6524 14112 6540 14176
rect 6604 14112 6620 14176
rect 6684 14112 6690 14176
rect 6374 14111 6690 14112
rect 11802 14176 12118 14177
rect 11802 14112 11808 14176
rect 11872 14112 11888 14176
rect 11952 14112 11968 14176
rect 12032 14112 12048 14176
rect 12112 14112 12118 14176
rect 11802 14111 12118 14112
rect 17230 14176 17546 14177
rect 17230 14112 17236 14176
rect 17300 14112 17316 14176
rect 17380 14112 17396 14176
rect 17460 14112 17476 14176
rect 17540 14112 17546 14176
rect 17230 14111 17546 14112
rect 22658 14176 22974 14177
rect 22658 14112 22664 14176
rect 22728 14112 22744 14176
rect 22808 14112 22824 14176
rect 22888 14112 22904 14176
rect 22968 14112 22974 14176
rect 22658 14111 22974 14112
rect 3660 13632 3976 13633
rect 3660 13568 3666 13632
rect 3730 13568 3746 13632
rect 3810 13568 3826 13632
rect 3890 13568 3906 13632
rect 3970 13568 3976 13632
rect 3660 13567 3976 13568
rect 9088 13632 9404 13633
rect 9088 13568 9094 13632
rect 9158 13568 9174 13632
rect 9238 13568 9254 13632
rect 9318 13568 9334 13632
rect 9398 13568 9404 13632
rect 9088 13567 9404 13568
rect 14516 13632 14832 13633
rect 14516 13568 14522 13632
rect 14586 13568 14602 13632
rect 14666 13568 14682 13632
rect 14746 13568 14762 13632
rect 14826 13568 14832 13632
rect 14516 13567 14832 13568
rect 19944 13632 20260 13633
rect 19944 13568 19950 13632
rect 20014 13568 20030 13632
rect 20094 13568 20110 13632
rect 20174 13568 20190 13632
rect 20254 13568 20260 13632
rect 19944 13567 20260 13568
rect 6374 13088 6690 13089
rect 6374 13024 6380 13088
rect 6444 13024 6460 13088
rect 6524 13024 6540 13088
rect 6604 13024 6620 13088
rect 6684 13024 6690 13088
rect 6374 13023 6690 13024
rect 11802 13088 12118 13089
rect 11802 13024 11808 13088
rect 11872 13024 11888 13088
rect 11952 13024 11968 13088
rect 12032 13024 12048 13088
rect 12112 13024 12118 13088
rect 11802 13023 12118 13024
rect 17230 13088 17546 13089
rect 17230 13024 17236 13088
rect 17300 13024 17316 13088
rect 17380 13024 17396 13088
rect 17460 13024 17476 13088
rect 17540 13024 17546 13088
rect 17230 13023 17546 13024
rect 22658 13088 22974 13089
rect 22658 13024 22664 13088
rect 22728 13024 22744 13088
rect 22808 13024 22824 13088
rect 22888 13024 22904 13088
rect 22968 13024 22974 13088
rect 22658 13023 22974 13024
rect 3660 12544 3976 12545
rect 3660 12480 3666 12544
rect 3730 12480 3746 12544
rect 3810 12480 3826 12544
rect 3890 12480 3906 12544
rect 3970 12480 3976 12544
rect 3660 12479 3976 12480
rect 9088 12544 9404 12545
rect 9088 12480 9094 12544
rect 9158 12480 9174 12544
rect 9238 12480 9254 12544
rect 9318 12480 9334 12544
rect 9398 12480 9404 12544
rect 9088 12479 9404 12480
rect 14516 12544 14832 12545
rect 14516 12480 14522 12544
rect 14586 12480 14602 12544
rect 14666 12480 14682 12544
rect 14746 12480 14762 12544
rect 14826 12480 14832 12544
rect 14516 12479 14832 12480
rect 19944 12544 20260 12545
rect 19944 12480 19950 12544
rect 20014 12480 20030 12544
rect 20094 12480 20110 12544
rect 20174 12480 20190 12544
rect 20254 12480 20260 12544
rect 19944 12479 20260 12480
rect 6374 12000 6690 12001
rect 0 11930 800 11960
rect 6374 11936 6380 12000
rect 6444 11936 6460 12000
rect 6524 11936 6540 12000
rect 6604 11936 6620 12000
rect 6684 11936 6690 12000
rect 6374 11935 6690 11936
rect 11802 12000 12118 12001
rect 11802 11936 11808 12000
rect 11872 11936 11888 12000
rect 11952 11936 11968 12000
rect 12032 11936 12048 12000
rect 12112 11936 12118 12000
rect 11802 11935 12118 11936
rect 17230 12000 17546 12001
rect 17230 11936 17236 12000
rect 17300 11936 17316 12000
rect 17380 11936 17396 12000
rect 17460 11936 17476 12000
rect 17540 11936 17546 12000
rect 17230 11935 17546 11936
rect 22658 12000 22974 12001
rect 22658 11936 22664 12000
rect 22728 11936 22744 12000
rect 22808 11936 22824 12000
rect 22888 11936 22904 12000
rect 22968 11936 22974 12000
rect 22658 11935 22974 11936
rect 933 11930 999 11933
rect 0 11928 999 11930
rect 0 11872 938 11928
rect 994 11872 999 11928
rect 0 11870 999 11872
rect 0 11840 800 11870
rect 933 11867 999 11870
rect 3660 11456 3976 11457
rect 3660 11392 3666 11456
rect 3730 11392 3746 11456
rect 3810 11392 3826 11456
rect 3890 11392 3906 11456
rect 3970 11392 3976 11456
rect 3660 11391 3976 11392
rect 9088 11456 9404 11457
rect 9088 11392 9094 11456
rect 9158 11392 9174 11456
rect 9238 11392 9254 11456
rect 9318 11392 9334 11456
rect 9398 11392 9404 11456
rect 9088 11391 9404 11392
rect 14516 11456 14832 11457
rect 14516 11392 14522 11456
rect 14586 11392 14602 11456
rect 14666 11392 14682 11456
rect 14746 11392 14762 11456
rect 14826 11392 14832 11456
rect 14516 11391 14832 11392
rect 19944 11456 20260 11457
rect 19944 11392 19950 11456
rect 20014 11392 20030 11456
rect 20094 11392 20110 11456
rect 20174 11392 20190 11456
rect 20254 11392 20260 11456
rect 19944 11391 20260 11392
rect 14273 11250 14339 11253
rect 16389 11250 16455 11253
rect 14273 11248 16455 11250
rect 14273 11192 14278 11248
rect 14334 11192 16394 11248
rect 16450 11192 16455 11248
rect 14273 11190 16455 11192
rect 14273 11187 14339 11190
rect 16389 11187 16455 11190
rect 15142 11052 15148 11116
rect 15212 11114 15218 11116
rect 15285 11114 15351 11117
rect 15212 11112 15351 11114
rect 15212 11056 15290 11112
rect 15346 11056 15351 11112
rect 15212 11054 15351 11056
rect 15212 11052 15218 11054
rect 15285 11051 15351 11054
rect 6374 10912 6690 10913
rect 6374 10848 6380 10912
rect 6444 10848 6460 10912
rect 6524 10848 6540 10912
rect 6604 10848 6620 10912
rect 6684 10848 6690 10912
rect 6374 10847 6690 10848
rect 11802 10912 12118 10913
rect 11802 10848 11808 10912
rect 11872 10848 11888 10912
rect 11952 10848 11968 10912
rect 12032 10848 12048 10912
rect 12112 10848 12118 10912
rect 11802 10847 12118 10848
rect 17230 10912 17546 10913
rect 17230 10848 17236 10912
rect 17300 10848 17316 10912
rect 17380 10848 17396 10912
rect 17460 10848 17476 10912
rect 17540 10848 17546 10912
rect 17230 10847 17546 10848
rect 22658 10912 22974 10913
rect 22658 10848 22664 10912
rect 22728 10848 22744 10912
rect 22808 10848 22824 10912
rect 22888 10848 22904 10912
rect 22968 10848 22974 10912
rect 22658 10847 22974 10848
rect 3660 10368 3976 10369
rect 3660 10304 3666 10368
rect 3730 10304 3746 10368
rect 3810 10304 3826 10368
rect 3890 10304 3906 10368
rect 3970 10304 3976 10368
rect 3660 10303 3976 10304
rect 9088 10368 9404 10369
rect 9088 10304 9094 10368
rect 9158 10304 9174 10368
rect 9238 10304 9254 10368
rect 9318 10304 9334 10368
rect 9398 10304 9404 10368
rect 9088 10303 9404 10304
rect 14516 10368 14832 10369
rect 14516 10304 14522 10368
rect 14586 10304 14602 10368
rect 14666 10304 14682 10368
rect 14746 10304 14762 10368
rect 14826 10304 14832 10368
rect 14516 10303 14832 10304
rect 19944 10368 20260 10369
rect 19944 10304 19950 10368
rect 20014 10304 20030 10368
rect 20094 10304 20110 10368
rect 20174 10304 20190 10368
rect 20254 10304 20260 10368
rect 19944 10303 20260 10304
rect 10961 10162 11027 10165
rect 17677 10162 17743 10165
rect 10961 10160 17743 10162
rect 10961 10104 10966 10160
rect 11022 10104 17682 10160
rect 17738 10104 17743 10160
rect 10961 10102 17743 10104
rect 10961 10099 11027 10102
rect 17677 10099 17743 10102
rect 6374 9824 6690 9825
rect 6374 9760 6380 9824
rect 6444 9760 6460 9824
rect 6524 9760 6540 9824
rect 6604 9760 6620 9824
rect 6684 9760 6690 9824
rect 6374 9759 6690 9760
rect 11802 9824 12118 9825
rect 11802 9760 11808 9824
rect 11872 9760 11888 9824
rect 11952 9760 11968 9824
rect 12032 9760 12048 9824
rect 12112 9760 12118 9824
rect 11802 9759 12118 9760
rect 17230 9824 17546 9825
rect 17230 9760 17236 9824
rect 17300 9760 17316 9824
rect 17380 9760 17396 9824
rect 17460 9760 17476 9824
rect 17540 9760 17546 9824
rect 17230 9759 17546 9760
rect 22658 9824 22974 9825
rect 22658 9760 22664 9824
rect 22728 9760 22744 9824
rect 22808 9760 22824 9824
rect 22888 9760 22904 9824
rect 22968 9760 22974 9824
rect 22658 9759 22974 9760
rect 3660 9280 3976 9281
rect 3660 9216 3666 9280
rect 3730 9216 3746 9280
rect 3810 9216 3826 9280
rect 3890 9216 3906 9280
rect 3970 9216 3976 9280
rect 3660 9215 3976 9216
rect 9088 9280 9404 9281
rect 9088 9216 9094 9280
rect 9158 9216 9174 9280
rect 9238 9216 9254 9280
rect 9318 9216 9334 9280
rect 9398 9216 9404 9280
rect 9088 9215 9404 9216
rect 14516 9280 14832 9281
rect 14516 9216 14522 9280
rect 14586 9216 14602 9280
rect 14666 9216 14682 9280
rect 14746 9216 14762 9280
rect 14826 9216 14832 9280
rect 14516 9215 14832 9216
rect 19944 9280 20260 9281
rect 19944 9216 19950 9280
rect 20014 9216 20030 9280
rect 20094 9216 20110 9280
rect 20174 9216 20190 9280
rect 20254 9216 20260 9280
rect 19944 9215 20260 9216
rect 6374 8736 6690 8737
rect 6374 8672 6380 8736
rect 6444 8672 6460 8736
rect 6524 8672 6540 8736
rect 6604 8672 6620 8736
rect 6684 8672 6690 8736
rect 6374 8671 6690 8672
rect 11802 8736 12118 8737
rect 11802 8672 11808 8736
rect 11872 8672 11888 8736
rect 11952 8672 11968 8736
rect 12032 8672 12048 8736
rect 12112 8672 12118 8736
rect 11802 8671 12118 8672
rect 17230 8736 17546 8737
rect 17230 8672 17236 8736
rect 17300 8672 17316 8736
rect 17380 8672 17396 8736
rect 17460 8672 17476 8736
rect 17540 8672 17546 8736
rect 17230 8671 17546 8672
rect 22658 8736 22974 8737
rect 22658 8672 22664 8736
rect 22728 8672 22744 8736
rect 22808 8672 22824 8736
rect 22888 8672 22904 8736
rect 22968 8672 22974 8736
rect 22658 8671 22974 8672
rect 15745 8530 15811 8533
rect 19149 8530 19215 8533
rect 15745 8528 19215 8530
rect 15745 8472 15750 8528
rect 15806 8472 19154 8528
rect 19210 8472 19215 8528
rect 15745 8470 19215 8472
rect 15745 8467 15811 8470
rect 19149 8467 19215 8470
rect 13905 8394 13971 8397
rect 17493 8394 17559 8397
rect 17861 8394 17927 8397
rect 13905 8392 17927 8394
rect 13905 8336 13910 8392
rect 13966 8336 17498 8392
rect 17554 8336 17866 8392
rect 17922 8336 17927 8392
rect 13905 8334 17927 8336
rect 13905 8331 13971 8334
rect 17493 8331 17559 8334
rect 17861 8331 17927 8334
rect 3660 8192 3976 8193
rect 3660 8128 3666 8192
rect 3730 8128 3746 8192
rect 3810 8128 3826 8192
rect 3890 8128 3906 8192
rect 3970 8128 3976 8192
rect 3660 8127 3976 8128
rect 9088 8192 9404 8193
rect 9088 8128 9094 8192
rect 9158 8128 9174 8192
rect 9238 8128 9254 8192
rect 9318 8128 9334 8192
rect 9398 8128 9404 8192
rect 9088 8127 9404 8128
rect 14516 8192 14832 8193
rect 14516 8128 14522 8192
rect 14586 8128 14602 8192
rect 14666 8128 14682 8192
rect 14746 8128 14762 8192
rect 14826 8128 14832 8192
rect 14516 8127 14832 8128
rect 19944 8192 20260 8193
rect 19944 8128 19950 8192
rect 20014 8128 20030 8192
rect 20094 8128 20110 8192
rect 20174 8128 20190 8192
rect 20254 8128 20260 8192
rect 19944 8127 20260 8128
rect 6374 7648 6690 7649
rect 6374 7584 6380 7648
rect 6444 7584 6460 7648
rect 6524 7584 6540 7648
rect 6604 7584 6620 7648
rect 6684 7584 6690 7648
rect 6374 7583 6690 7584
rect 11802 7648 12118 7649
rect 11802 7584 11808 7648
rect 11872 7584 11888 7648
rect 11952 7584 11968 7648
rect 12032 7584 12048 7648
rect 12112 7584 12118 7648
rect 11802 7583 12118 7584
rect 17230 7648 17546 7649
rect 17230 7584 17236 7648
rect 17300 7584 17316 7648
rect 17380 7584 17396 7648
rect 17460 7584 17476 7648
rect 17540 7584 17546 7648
rect 17230 7583 17546 7584
rect 22658 7648 22974 7649
rect 22658 7584 22664 7648
rect 22728 7584 22744 7648
rect 22808 7584 22824 7648
rect 22888 7584 22904 7648
rect 22968 7584 22974 7648
rect 22658 7583 22974 7584
rect 12985 7442 13051 7445
rect 15142 7442 15148 7444
rect 12985 7440 15148 7442
rect 12985 7384 12990 7440
rect 13046 7384 15148 7440
rect 12985 7382 15148 7384
rect 12985 7379 13051 7382
rect 15142 7380 15148 7382
rect 15212 7380 15218 7444
rect 3660 7104 3976 7105
rect 3660 7040 3666 7104
rect 3730 7040 3746 7104
rect 3810 7040 3826 7104
rect 3890 7040 3906 7104
rect 3970 7040 3976 7104
rect 3660 7039 3976 7040
rect 9088 7104 9404 7105
rect 9088 7040 9094 7104
rect 9158 7040 9174 7104
rect 9238 7040 9254 7104
rect 9318 7040 9334 7104
rect 9398 7040 9404 7104
rect 9088 7039 9404 7040
rect 14516 7104 14832 7105
rect 14516 7040 14522 7104
rect 14586 7040 14602 7104
rect 14666 7040 14682 7104
rect 14746 7040 14762 7104
rect 14826 7040 14832 7104
rect 14516 7039 14832 7040
rect 19944 7104 20260 7105
rect 19944 7040 19950 7104
rect 20014 7040 20030 7104
rect 20094 7040 20110 7104
rect 20174 7040 20190 7104
rect 20254 7040 20260 7104
rect 19944 7039 20260 7040
rect 6374 6560 6690 6561
rect 6374 6496 6380 6560
rect 6444 6496 6460 6560
rect 6524 6496 6540 6560
rect 6604 6496 6620 6560
rect 6684 6496 6690 6560
rect 6374 6495 6690 6496
rect 11802 6560 12118 6561
rect 11802 6496 11808 6560
rect 11872 6496 11888 6560
rect 11952 6496 11968 6560
rect 12032 6496 12048 6560
rect 12112 6496 12118 6560
rect 11802 6495 12118 6496
rect 17230 6560 17546 6561
rect 17230 6496 17236 6560
rect 17300 6496 17316 6560
rect 17380 6496 17396 6560
rect 17460 6496 17476 6560
rect 17540 6496 17546 6560
rect 17230 6495 17546 6496
rect 22658 6560 22974 6561
rect 22658 6496 22664 6560
rect 22728 6496 22744 6560
rect 22808 6496 22824 6560
rect 22888 6496 22904 6560
rect 22968 6496 22974 6560
rect 22658 6495 22974 6496
rect 3660 6016 3976 6017
rect 3660 5952 3666 6016
rect 3730 5952 3746 6016
rect 3810 5952 3826 6016
rect 3890 5952 3906 6016
rect 3970 5952 3976 6016
rect 3660 5951 3976 5952
rect 9088 6016 9404 6017
rect 9088 5952 9094 6016
rect 9158 5952 9174 6016
rect 9238 5952 9254 6016
rect 9318 5952 9334 6016
rect 9398 5952 9404 6016
rect 9088 5951 9404 5952
rect 14516 6016 14832 6017
rect 14516 5952 14522 6016
rect 14586 5952 14602 6016
rect 14666 5952 14682 6016
rect 14746 5952 14762 6016
rect 14826 5952 14832 6016
rect 14516 5951 14832 5952
rect 19944 6016 20260 6017
rect 19944 5952 19950 6016
rect 20014 5952 20030 6016
rect 20094 5952 20110 6016
rect 20174 5952 20190 6016
rect 20254 5952 20260 6016
rect 19944 5951 20260 5952
rect 6374 5472 6690 5473
rect 6374 5408 6380 5472
rect 6444 5408 6460 5472
rect 6524 5408 6540 5472
rect 6604 5408 6620 5472
rect 6684 5408 6690 5472
rect 6374 5407 6690 5408
rect 11802 5472 12118 5473
rect 11802 5408 11808 5472
rect 11872 5408 11888 5472
rect 11952 5408 11968 5472
rect 12032 5408 12048 5472
rect 12112 5408 12118 5472
rect 11802 5407 12118 5408
rect 17230 5472 17546 5473
rect 17230 5408 17236 5472
rect 17300 5408 17316 5472
rect 17380 5408 17396 5472
rect 17460 5408 17476 5472
rect 17540 5408 17546 5472
rect 17230 5407 17546 5408
rect 22658 5472 22974 5473
rect 22658 5408 22664 5472
rect 22728 5408 22744 5472
rect 22808 5408 22824 5472
rect 22888 5408 22904 5472
rect 22968 5408 22974 5472
rect 22658 5407 22974 5408
rect 13077 5130 13143 5133
rect 14733 5130 14799 5133
rect 13077 5128 14799 5130
rect 13077 5072 13082 5128
rect 13138 5072 14738 5128
rect 14794 5072 14799 5128
rect 13077 5070 14799 5072
rect 13077 5067 13143 5070
rect 14733 5067 14799 5070
rect 3660 4928 3976 4929
rect 3660 4864 3666 4928
rect 3730 4864 3746 4928
rect 3810 4864 3826 4928
rect 3890 4864 3906 4928
rect 3970 4864 3976 4928
rect 3660 4863 3976 4864
rect 9088 4928 9404 4929
rect 9088 4864 9094 4928
rect 9158 4864 9174 4928
rect 9238 4864 9254 4928
rect 9318 4864 9334 4928
rect 9398 4864 9404 4928
rect 9088 4863 9404 4864
rect 14516 4928 14832 4929
rect 14516 4864 14522 4928
rect 14586 4864 14602 4928
rect 14666 4864 14682 4928
rect 14746 4864 14762 4928
rect 14826 4864 14832 4928
rect 14516 4863 14832 4864
rect 19944 4928 20260 4929
rect 19944 4864 19950 4928
rect 20014 4864 20030 4928
rect 20094 4864 20110 4928
rect 20174 4864 20190 4928
rect 20254 4864 20260 4928
rect 19944 4863 20260 4864
rect 6374 4384 6690 4385
rect 6374 4320 6380 4384
rect 6444 4320 6460 4384
rect 6524 4320 6540 4384
rect 6604 4320 6620 4384
rect 6684 4320 6690 4384
rect 6374 4319 6690 4320
rect 11802 4384 12118 4385
rect 11802 4320 11808 4384
rect 11872 4320 11888 4384
rect 11952 4320 11968 4384
rect 12032 4320 12048 4384
rect 12112 4320 12118 4384
rect 11802 4319 12118 4320
rect 17230 4384 17546 4385
rect 17230 4320 17236 4384
rect 17300 4320 17316 4384
rect 17380 4320 17396 4384
rect 17460 4320 17476 4384
rect 17540 4320 17546 4384
rect 17230 4319 17546 4320
rect 22658 4384 22974 4385
rect 22658 4320 22664 4384
rect 22728 4320 22744 4384
rect 22808 4320 22824 4384
rect 22888 4320 22904 4384
rect 22968 4320 22974 4384
rect 22658 4319 22974 4320
rect 0 4042 800 4072
rect 3141 4042 3207 4045
rect 0 4040 3207 4042
rect 0 3984 3146 4040
rect 3202 3984 3207 4040
rect 0 3982 3207 3984
rect 0 3952 800 3982
rect 3141 3979 3207 3982
rect 3660 3840 3976 3841
rect 3660 3776 3666 3840
rect 3730 3776 3746 3840
rect 3810 3776 3826 3840
rect 3890 3776 3906 3840
rect 3970 3776 3976 3840
rect 3660 3775 3976 3776
rect 9088 3840 9404 3841
rect 9088 3776 9094 3840
rect 9158 3776 9174 3840
rect 9238 3776 9254 3840
rect 9318 3776 9334 3840
rect 9398 3776 9404 3840
rect 9088 3775 9404 3776
rect 14516 3840 14832 3841
rect 14516 3776 14522 3840
rect 14586 3776 14602 3840
rect 14666 3776 14682 3840
rect 14746 3776 14762 3840
rect 14826 3776 14832 3840
rect 14516 3775 14832 3776
rect 19944 3840 20260 3841
rect 19944 3776 19950 3840
rect 20014 3776 20030 3840
rect 20094 3776 20110 3840
rect 20174 3776 20190 3840
rect 20254 3776 20260 3840
rect 19944 3775 20260 3776
rect 10961 3498 11027 3501
rect 19425 3498 19491 3501
rect 10961 3496 19491 3498
rect 10961 3440 10966 3496
rect 11022 3440 19430 3496
rect 19486 3440 19491 3496
rect 10961 3438 19491 3440
rect 10961 3435 11027 3438
rect 19425 3435 19491 3438
rect 6374 3296 6690 3297
rect 6374 3232 6380 3296
rect 6444 3232 6460 3296
rect 6524 3232 6540 3296
rect 6604 3232 6620 3296
rect 6684 3232 6690 3296
rect 6374 3231 6690 3232
rect 11802 3296 12118 3297
rect 11802 3232 11808 3296
rect 11872 3232 11888 3296
rect 11952 3232 11968 3296
rect 12032 3232 12048 3296
rect 12112 3232 12118 3296
rect 11802 3231 12118 3232
rect 17230 3296 17546 3297
rect 17230 3232 17236 3296
rect 17300 3232 17316 3296
rect 17380 3232 17396 3296
rect 17460 3232 17476 3296
rect 17540 3232 17546 3296
rect 17230 3231 17546 3232
rect 22658 3296 22974 3297
rect 22658 3232 22664 3296
rect 22728 3232 22744 3296
rect 22808 3232 22824 3296
rect 22888 3232 22904 3296
rect 22968 3232 22974 3296
rect 22658 3231 22974 3232
rect 3660 2752 3976 2753
rect 3660 2688 3666 2752
rect 3730 2688 3746 2752
rect 3810 2688 3826 2752
rect 3890 2688 3906 2752
rect 3970 2688 3976 2752
rect 3660 2687 3976 2688
rect 9088 2752 9404 2753
rect 9088 2688 9094 2752
rect 9158 2688 9174 2752
rect 9238 2688 9254 2752
rect 9318 2688 9334 2752
rect 9398 2688 9404 2752
rect 9088 2687 9404 2688
rect 14516 2752 14832 2753
rect 14516 2688 14522 2752
rect 14586 2688 14602 2752
rect 14666 2688 14682 2752
rect 14746 2688 14762 2752
rect 14826 2688 14832 2752
rect 14516 2687 14832 2688
rect 19944 2752 20260 2753
rect 19944 2688 19950 2752
rect 20014 2688 20030 2752
rect 20094 2688 20110 2752
rect 20174 2688 20190 2752
rect 20254 2688 20260 2752
rect 19944 2687 20260 2688
rect 6374 2208 6690 2209
rect 6374 2144 6380 2208
rect 6444 2144 6460 2208
rect 6524 2144 6540 2208
rect 6604 2144 6620 2208
rect 6684 2144 6690 2208
rect 6374 2143 6690 2144
rect 11802 2208 12118 2209
rect 11802 2144 11808 2208
rect 11872 2144 11888 2208
rect 11952 2144 11968 2208
rect 12032 2144 12048 2208
rect 12112 2144 12118 2208
rect 11802 2143 12118 2144
rect 17230 2208 17546 2209
rect 17230 2144 17236 2208
rect 17300 2144 17316 2208
rect 17380 2144 17396 2208
rect 17460 2144 17476 2208
rect 17540 2144 17546 2208
rect 17230 2143 17546 2144
rect 22658 2208 22974 2209
rect 22658 2144 22664 2208
rect 22728 2144 22744 2208
rect 22808 2144 22824 2208
rect 22888 2144 22904 2208
rect 22968 2144 22974 2208
rect 22658 2143 22974 2144
<< via3 >>
rect 6380 21788 6444 21792
rect 6380 21732 6384 21788
rect 6384 21732 6440 21788
rect 6440 21732 6444 21788
rect 6380 21728 6444 21732
rect 6460 21788 6524 21792
rect 6460 21732 6464 21788
rect 6464 21732 6520 21788
rect 6520 21732 6524 21788
rect 6460 21728 6524 21732
rect 6540 21788 6604 21792
rect 6540 21732 6544 21788
rect 6544 21732 6600 21788
rect 6600 21732 6604 21788
rect 6540 21728 6604 21732
rect 6620 21788 6684 21792
rect 6620 21732 6624 21788
rect 6624 21732 6680 21788
rect 6680 21732 6684 21788
rect 6620 21728 6684 21732
rect 11808 21788 11872 21792
rect 11808 21732 11812 21788
rect 11812 21732 11868 21788
rect 11868 21732 11872 21788
rect 11808 21728 11872 21732
rect 11888 21788 11952 21792
rect 11888 21732 11892 21788
rect 11892 21732 11948 21788
rect 11948 21732 11952 21788
rect 11888 21728 11952 21732
rect 11968 21788 12032 21792
rect 11968 21732 11972 21788
rect 11972 21732 12028 21788
rect 12028 21732 12032 21788
rect 11968 21728 12032 21732
rect 12048 21788 12112 21792
rect 12048 21732 12052 21788
rect 12052 21732 12108 21788
rect 12108 21732 12112 21788
rect 12048 21728 12112 21732
rect 17236 21788 17300 21792
rect 17236 21732 17240 21788
rect 17240 21732 17296 21788
rect 17296 21732 17300 21788
rect 17236 21728 17300 21732
rect 17316 21788 17380 21792
rect 17316 21732 17320 21788
rect 17320 21732 17376 21788
rect 17376 21732 17380 21788
rect 17316 21728 17380 21732
rect 17396 21788 17460 21792
rect 17396 21732 17400 21788
rect 17400 21732 17456 21788
rect 17456 21732 17460 21788
rect 17396 21728 17460 21732
rect 17476 21788 17540 21792
rect 17476 21732 17480 21788
rect 17480 21732 17536 21788
rect 17536 21732 17540 21788
rect 17476 21728 17540 21732
rect 22664 21788 22728 21792
rect 22664 21732 22668 21788
rect 22668 21732 22724 21788
rect 22724 21732 22728 21788
rect 22664 21728 22728 21732
rect 22744 21788 22808 21792
rect 22744 21732 22748 21788
rect 22748 21732 22804 21788
rect 22804 21732 22808 21788
rect 22744 21728 22808 21732
rect 22824 21788 22888 21792
rect 22824 21732 22828 21788
rect 22828 21732 22884 21788
rect 22884 21732 22888 21788
rect 22824 21728 22888 21732
rect 22904 21788 22968 21792
rect 22904 21732 22908 21788
rect 22908 21732 22964 21788
rect 22964 21732 22968 21788
rect 22904 21728 22968 21732
rect 3666 21244 3730 21248
rect 3666 21188 3670 21244
rect 3670 21188 3726 21244
rect 3726 21188 3730 21244
rect 3666 21184 3730 21188
rect 3746 21244 3810 21248
rect 3746 21188 3750 21244
rect 3750 21188 3806 21244
rect 3806 21188 3810 21244
rect 3746 21184 3810 21188
rect 3826 21244 3890 21248
rect 3826 21188 3830 21244
rect 3830 21188 3886 21244
rect 3886 21188 3890 21244
rect 3826 21184 3890 21188
rect 3906 21244 3970 21248
rect 3906 21188 3910 21244
rect 3910 21188 3966 21244
rect 3966 21188 3970 21244
rect 3906 21184 3970 21188
rect 9094 21244 9158 21248
rect 9094 21188 9098 21244
rect 9098 21188 9154 21244
rect 9154 21188 9158 21244
rect 9094 21184 9158 21188
rect 9174 21244 9238 21248
rect 9174 21188 9178 21244
rect 9178 21188 9234 21244
rect 9234 21188 9238 21244
rect 9174 21184 9238 21188
rect 9254 21244 9318 21248
rect 9254 21188 9258 21244
rect 9258 21188 9314 21244
rect 9314 21188 9318 21244
rect 9254 21184 9318 21188
rect 9334 21244 9398 21248
rect 9334 21188 9338 21244
rect 9338 21188 9394 21244
rect 9394 21188 9398 21244
rect 9334 21184 9398 21188
rect 14522 21244 14586 21248
rect 14522 21188 14526 21244
rect 14526 21188 14582 21244
rect 14582 21188 14586 21244
rect 14522 21184 14586 21188
rect 14602 21244 14666 21248
rect 14602 21188 14606 21244
rect 14606 21188 14662 21244
rect 14662 21188 14666 21244
rect 14602 21184 14666 21188
rect 14682 21244 14746 21248
rect 14682 21188 14686 21244
rect 14686 21188 14742 21244
rect 14742 21188 14746 21244
rect 14682 21184 14746 21188
rect 14762 21244 14826 21248
rect 14762 21188 14766 21244
rect 14766 21188 14822 21244
rect 14822 21188 14826 21244
rect 14762 21184 14826 21188
rect 19950 21244 20014 21248
rect 19950 21188 19954 21244
rect 19954 21188 20010 21244
rect 20010 21188 20014 21244
rect 19950 21184 20014 21188
rect 20030 21244 20094 21248
rect 20030 21188 20034 21244
rect 20034 21188 20090 21244
rect 20090 21188 20094 21244
rect 20030 21184 20094 21188
rect 20110 21244 20174 21248
rect 20110 21188 20114 21244
rect 20114 21188 20170 21244
rect 20170 21188 20174 21244
rect 20110 21184 20174 21188
rect 20190 21244 20254 21248
rect 20190 21188 20194 21244
rect 20194 21188 20250 21244
rect 20250 21188 20254 21244
rect 20190 21184 20254 21188
rect 6380 20700 6444 20704
rect 6380 20644 6384 20700
rect 6384 20644 6440 20700
rect 6440 20644 6444 20700
rect 6380 20640 6444 20644
rect 6460 20700 6524 20704
rect 6460 20644 6464 20700
rect 6464 20644 6520 20700
rect 6520 20644 6524 20700
rect 6460 20640 6524 20644
rect 6540 20700 6604 20704
rect 6540 20644 6544 20700
rect 6544 20644 6600 20700
rect 6600 20644 6604 20700
rect 6540 20640 6604 20644
rect 6620 20700 6684 20704
rect 6620 20644 6624 20700
rect 6624 20644 6680 20700
rect 6680 20644 6684 20700
rect 6620 20640 6684 20644
rect 11808 20700 11872 20704
rect 11808 20644 11812 20700
rect 11812 20644 11868 20700
rect 11868 20644 11872 20700
rect 11808 20640 11872 20644
rect 11888 20700 11952 20704
rect 11888 20644 11892 20700
rect 11892 20644 11948 20700
rect 11948 20644 11952 20700
rect 11888 20640 11952 20644
rect 11968 20700 12032 20704
rect 11968 20644 11972 20700
rect 11972 20644 12028 20700
rect 12028 20644 12032 20700
rect 11968 20640 12032 20644
rect 12048 20700 12112 20704
rect 12048 20644 12052 20700
rect 12052 20644 12108 20700
rect 12108 20644 12112 20700
rect 12048 20640 12112 20644
rect 17236 20700 17300 20704
rect 17236 20644 17240 20700
rect 17240 20644 17296 20700
rect 17296 20644 17300 20700
rect 17236 20640 17300 20644
rect 17316 20700 17380 20704
rect 17316 20644 17320 20700
rect 17320 20644 17376 20700
rect 17376 20644 17380 20700
rect 17316 20640 17380 20644
rect 17396 20700 17460 20704
rect 17396 20644 17400 20700
rect 17400 20644 17456 20700
rect 17456 20644 17460 20700
rect 17396 20640 17460 20644
rect 17476 20700 17540 20704
rect 17476 20644 17480 20700
rect 17480 20644 17536 20700
rect 17536 20644 17540 20700
rect 17476 20640 17540 20644
rect 22664 20700 22728 20704
rect 22664 20644 22668 20700
rect 22668 20644 22724 20700
rect 22724 20644 22728 20700
rect 22664 20640 22728 20644
rect 22744 20700 22808 20704
rect 22744 20644 22748 20700
rect 22748 20644 22804 20700
rect 22804 20644 22808 20700
rect 22744 20640 22808 20644
rect 22824 20700 22888 20704
rect 22824 20644 22828 20700
rect 22828 20644 22884 20700
rect 22884 20644 22888 20700
rect 22824 20640 22888 20644
rect 22904 20700 22968 20704
rect 22904 20644 22908 20700
rect 22908 20644 22964 20700
rect 22964 20644 22968 20700
rect 22904 20640 22968 20644
rect 3666 20156 3730 20160
rect 3666 20100 3670 20156
rect 3670 20100 3726 20156
rect 3726 20100 3730 20156
rect 3666 20096 3730 20100
rect 3746 20156 3810 20160
rect 3746 20100 3750 20156
rect 3750 20100 3806 20156
rect 3806 20100 3810 20156
rect 3746 20096 3810 20100
rect 3826 20156 3890 20160
rect 3826 20100 3830 20156
rect 3830 20100 3886 20156
rect 3886 20100 3890 20156
rect 3826 20096 3890 20100
rect 3906 20156 3970 20160
rect 3906 20100 3910 20156
rect 3910 20100 3966 20156
rect 3966 20100 3970 20156
rect 3906 20096 3970 20100
rect 9094 20156 9158 20160
rect 9094 20100 9098 20156
rect 9098 20100 9154 20156
rect 9154 20100 9158 20156
rect 9094 20096 9158 20100
rect 9174 20156 9238 20160
rect 9174 20100 9178 20156
rect 9178 20100 9234 20156
rect 9234 20100 9238 20156
rect 9174 20096 9238 20100
rect 9254 20156 9318 20160
rect 9254 20100 9258 20156
rect 9258 20100 9314 20156
rect 9314 20100 9318 20156
rect 9254 20096 9318 20100
rect 9334 20156 9398 20160
rect 9334 20100 9338 20156
rect 9338 20100 9394 20156
rect 9394 20100 9398 20156
rect 9334 20096 9398 20100
rect 14522 20156 14586 20160
rect 14522 20100 14526 20156
rect 14526 20100 14582 20156
rect 14582 20100 14586 20156
rect 14522 20096 14586 20100
rect 14602 20156 14666 20160
rect 14602 20100 14606 20156
rect 14606 20100 14662 20156
rect 14662 20100 14666 20156
rect 14602 20096 14666 20100
rect 14682 20156 14746 20160
rect 14682 20100 14686 20156
rect 14686 20100 14742 20156
rect 14742 20100 14746 20156
rect 14682 20096 14746 20100
rect 14762 20156 14826 20160
rect 14762 20100 14766 20156
rect 14766 20100 14822 20156
rect 14822 20100 14826 20156
rect 14762 20096 14826 20100
rect 19950 20156 20014 20160
rect 19950 20100 19954 20156
rect 19954 20100 20010 20156
rect 20010 20100 20014 20156
rect 19950 20096 20014 20100
rect 20030 20156 20094 20160
rect 20030 20100 20034 20156
rect 20034 20100 20090 20156
rect 20090 20100 20094 20156
rect 20030 20096 20094 20100
rect 20110 20156 20174 20160
rect 20110 20100 20114 20156
rect 20114 20100 20170 20156
rect 20170 20100 20174 20156
rect 20110 20096 20174 20100
rect 20190 20156 20254 20160
rect 20190 20100 20194 20156
rect 20194 20100 20250 20156
rect 20250 20100 20254 20156
rect 20190 20096 20254 20100
rect 6380 19612 6444 19616
rect 6380 19556 6384 19612
rect 6384 19556 6440 19612
rect 6440 19556 6444 19612
rect 6380 19552 6444 19556
rect 6460 19612 6524 19616
rect 6460 19556 6464 19612
rect 6464 19556 6520 19612
rect 6520 19556 6524 19612
rect 6460 19552 6524 19556
rect 6540 19612 6604 19616
rect 6540 19556 6544 19612
rect 6544 19556 6600 19612
rect 6600 19556 6604 19612
rect 6540 19552 6604 19556
rect 6620 19612 6684 19616
rect 6620 19556 6624 19612
rect 6624 19556 6680 19612
rect 6680 19556 6684 19612
rect 6620 19552 6684 19556
rect 11808 19612 11872 19616
rect 11808 19556 11812 19612
rect 11812 19556 11868 19612
rect 11868 19556 11872 19612
rect 11808 19552 11872 19556
rect 11888 19612 11952 19616
rect 11888 19556 11892 19612
rect 11892 19556 11948 19612
rect 11948 19556 11952 19612
rect 11888 19552 11952 19556
rect 11968 19612 12032 19616
rect 11968 19556 11972 19612
rect 11972 19556 12028 19612
rect 12028 19556 12032 19612
rect 11968 19552 12032 19556
rect 12048 19612 12112 19616
rect 12048 19556 12052 19612
rect 12052 19556 12108 19612
rect 12108 19556 12112 19612
rect 12048 19552 12112 19556
rect 17236 19612 17300 19616
rect 17236 19556 17240 19612
rect 17240 19556 17296 19612
rect 17296 19556 17300 19612
rect 17236 19552 17300 19556
rect 17316 19612 17380 19616
rect 17316 19556 17320 19612
rect 17320 19556 17376 19612
rect 17376 19556 17380 19612
rect 17316 19552 17380 19556
rect 17396 19612 17460 19616
rect 17396 19556 17400 19612
rect 17400 19556 17456 19612
rect 17456 19556 17460 19612
rect 17396 19552 17460 19556
rect 17476 19612 17540 19616
rect 17476 19556 17480 19612
rect 17480 19556 17536 19612
rect 17536 19556 17540 19612
rect 17476 19552 17540 19556
rect 22664 19612 22728 19616
rect 22664 19556 22668 19612
rect 22668 19556 22724 19612
rect 22724 19556 22728 19612
rect 22664 19552 22728 19556
rect 22744 19612 22808 19616
rect 22744 19556 22748 19612
rect 22748 19556 22804 19612
rect 22804 19556 22808 19612
rect 22744 19552 22808 19556
rect 22824 19612 22888 19616
rect 22824 19556 22828 19612
rect 22828 19556 22884 19612
rect 22884 19556 22888 19612
rect 22824 19552 22888 19556
rect 22904 19612 22968 19616
rect 22904 19556 22908 19612
rect 22908 19556 22964 19612
rect 22964 19556 22968 19612
rect 22904 19552 22968 19556
rect 3666 19068 3730 19072
rect 3666 19012 3670 19068
rect 3670 19012 3726 19068
rect 3726 19012 3730 19068
rect 3666 19008 3730 19012
rect 3746 19068 3810 19072
rect 3746 19012 3750 19068
rect 3750 19012 3806 19068
rect 3806 19012 3810 19068
rect 3746 19008 3810 19012
rect 3826 19068 3890 19072
rect 3826 19012 3830 19068
rect 3830 19012 3886 19068
rect 3886 19012 3890 19068
rect 3826 19008 3890 19012
rect 3906 19068 3970 19072
rect 3906 19012 3910 19068
rect 3910 19012 3966 19068
rect 3966 19012 3970 19068
rect 3906 19008 3970 19012
rect 9094 19068 9158 19072
rect 9094 19012 9098 19068
rect 9098 19012 9154 19068
rect 9154 19012 9158 19068
rect 9094 19008 9158 19012
rect 9174 19068 9238 19072
rect 9174 19012 9178 19068
rect 9178 19012 9234 19068
rect 9234 19012 9238 19068
rect 9174 19008 9238 19012
rect 9254 19068 9318 19072
rect 9254 19012 9258 19068
rect 9258 19012 9314 19068
rect 9314 19012 9318 19068
rect 9254 19008 9318 19012
rect 9334 19068 9398 19072
rect 9334 19012 9338 19068
rect 9338 19012 9394 19068
rect 9394 19012 9398 19068
rect 9334 19008 9398 19012
rect 14522 19068 14586 19072
rect 14522 19012 14526 19068
rect 14526 19012 14582 19068
rect 14582 19012 14586 19068
rect 14522 19008 14586 19012
rect 14602 19068 14666 19072
rect 14602 19012 14606 19068
rect 14606 19012 14662 19068
rect 14662 19012 14666 19068
rect 14602 19008 14666 19012
rect 14682 19068 14746 19072
rect 14682 19012 14686 19068
rect 14686 19012 14742 19068
rect 14742 19012 14746 19068
rect 14682 19008 14746 19012
rect 14762 19068 14826 19072
rect 14762 19012 14766 19068
rect 14766 19012 14822 19068
rect 14822 19012 14826 19068
rect 14762 19008 14826 19012
rect 19950 19068 20014 19072
rect 19950 19012 19954 19068
rect 19954 19012 20010 19068
rect 20010 19012 20014 19068
rect 19950 19008 20014 19012
rect 20030 19068 20094 19072
rect 20030 19012 20034 19068
rect 20034 19012 20090 19068
rect 20090 19012 20094 19068
rect 20030 19008 20094 19012
rect 20110 19068 20174 19072
rect 20110 19012 20114 19068
rect 20114 19012 20170 19068
rect 20170 19012 20174 19068
rect 20110 19008 20174 19012
rect 20190 19068 20254 19072
rect 20190 19012 20194 19068
rect 20194 19012 20250 19068
rect 20250 19012 20254 19068
rect 20190 19008 20254 19012
rect 6380 18524 6444 18528
rect 6380 18468 6384 18524
rect 6384 18468 6440 18524
rect 6440 18468 6444 18524
rect 6380 18464 6444 18468
rect 6460 18524 6524 18528
rect 6460 18468 6464 18524
rect 6464 18468 6520 18524
rect 6520 18468 6524 18524
rect 6460 18464 6524 18468
rect 6540 18524 6604 18528
rect 6540 18468 6544 18524
rect 6544 18468 6600 18524
rect 6600 18468 6604 18524
rect 6540 18464 6604 18468
rect 6620 18524 6684 18528
rect 6620 18468 6624 18524
rect 6624 18468 6680 18524
rect 6680 18468 6684 18524
rect 6620 18464 6684 18468
rect 11808 18524 11872 18528
rect 11808 18468 11812 18524
rect 11812 18468 11868 18524
rect 11868 18468 11872 18524
rect 11808 18464 11872 18468
rect 11888 18524 11952 18528
rect 11888 18468 11892 18524
rect 11892 18468 11948 18524
rect 11948 18468 11952 18524
rect 11888 18464 11952 18468
rect 11968 18524 12032 18528
rect 11968 18468 11972 18524
rect 11972 18468 12028 18524
rect 12028 18468 12032 18524
rect 11968 18464 12032 18468
rect 12048 18524 12112 18528
rect 12048 18468 12052 18524
rect 12052 18468 12108 18524
rect 12108 18468 12112 18524
rect 12048 18464 12112 18468
rect 17236 18524 17300 18528
rect 17236 18468 17240 18524
rect 17240 18468 17296 18524
rect 17296 18468 17300 18524
rect 17236 18464 17300 18468
rect 17316 18524 17380 18528
rect 17316 18468 17320 18524
rect 17320 18468 17376 18524
rect 17376 18468 17380 18524
rect 17316 18464 17380 18468
rect 17396 18524 17460 18528
rect 17396 18468 17400 18524
rect 17400 18468 17456 18524
rect 17456 18468 17460 18524
rect 17396 18464 17460 18468
rect 17476 18524 17540 18528
rect 17476 18468 17480 18524
rect 17480 18468 17536 18524
rect 17536 18468 17540 18524
rect 17476 18464 17540 18468
rect 22664 18524 22728 18528
rect 22664 18468 22668 18524
rect 22668 18468 22724 18524
rect 22724 18468 22728 18524
rect 22664 18464 22728 18468
rect 22744 18524 22808 18528
rect 22744 18468 22748 18524
rect 22748 18468 22804 18524
rect 22804 18468 22808 18524
rect 22744 18464 22808 18468
rect 22824 18524 22888 18528
rect 22824 18468 22828 18524
rect 22828 18468 22884 18524
rect 22884 18468 22888 18524
rect 22824 18464 22888 18468
rect 22904 18524 22968 18528
rect 22904 18468 22908 18524
rect 22908 18468 22964 18524
rect 22964 18468 22968 18524
rect 22904 18464 22968 18468
rect 3666 17980 3730 17984
rect 3666 17924 3670 17980
rect 3670 17924 3726 17980
rect 3726 17924 3730 17980
rect 3666 17920 3730 17924
rect 3746 17980 3810 17984
rect 3746 17924 3750 17980
rect 3750 17924 3806 17980
rect 3806 17924 3810 17980
rect 3746 17920 3810 17924
rect 3826 17980 3890 17984
rect 3826 17924 3830 17980
rect 3830 17924 3886 17980
rect 3886 17924 3890 17980
rect 3826 17920 3890 17924
rect 3906 17980 3970 17984
rect 3906 17924 3910 17980
rect 3910 17924 3966 17980
rect 3966 17924 3970 17980
rect 3906 17920 3970 17924
rect 9094 17980 9158 17984
rect 9094 17924 9098 17980
rect 9098 17924 9154 17980
rect 9154 17924 9158 17980
rect 9094 17920 9158 17924
rect 9174 17980 9238 17984
rect 9174 17924 9178 17980
rect 9178 17924 9234 17980
rect 9234 17924 9238 17980
rect 9174 17920 9238 17924
rect 9254 17980 9318 17984
rect 9254 17924 9258 17980
rect 9258 17924 9314 17980
rect 9314 17924 9318 17980
rect 9254 17920 9318 17924
rect 9334 17980 9398 17984
rect 9334 17924 9338 17980
rect 9338 17924 9394 17980
rect 9394 17924 9398 17980
rect 9334 17920 9398 17924
rect 14522 17980 14586 17984
rect 14522 17924 14526 17980
rect 14526 17924 14582 17980
rect 14582 17924 14586 17980
rect 14522 17920 14586 17924
rect 14602 17980 14666 17984
rect 14602 17924 14606 17980
rect 14606 17924 14662 17980
rect 14662 17924 14666 17980
rect 14602 17920 14666 17924
rect 14682 17980 14746 17984
rect 14682 17924 14686 17980
rect 14686 17924 14742 17980
rect 14742 17924 14746 17980
rect 14682 17920 14746 17924
rect 14762 17980 14826 17984
rect 14762 17924 14766 17980
rect 14766 17924 14822 17980
rect 14822 17924 14826 17980
rect 14762 17920 14826 17924
rect 19950 17980 20014 17984
rect 19950 17924 19954 17980
rect 19954 17924 20010 17980
rect 20010 17924 20014 17980
rect 19950 17920 20014 17924
rect 20030 17980 20094 17984
rect 20030 17924 20034 17980
rect 20034 17924 20090 17980
rect 20090 17924 20094 17980
rect 20030 17920 20094 17924
rect 20110 17980 20174 17984
rect 20110 17924 20114 17980
rect 20114 17924 20170 17980
rect 20170 17924 20174 17980
rect 20110 17920 20174 17924
rect 20190 17980 20254 17984
rect 20190 17924 20194 17980
rect 20194 17924 20250 17980
rect 20250 17924 20254 17980
rect 20190 17920 20254 17924
rect 6380 17436 6444 17440
rect 6380 17380 6384 17436
rect 6384 17380 6440 17436
rect 6440 17380 6444 17436
rect 6380 17376 6444 17380
rect 6460 17436 6524 17440
rect 6460 17380 6464 17436
rect 6464 17380 6520 17436
rect 6520 17380 6524 17436
rect 6460 17376 6524 17380
rect 6540 17436 6604 17440
rect 6540 17380 6544 17436
rect 6544 17380 6600 17436
rect 6600 17380 6604 17436
rect 6540 17376 6604 17380
rect 6620 17436 6684 17440
rect 6620 17380 6624 17436
rect 6624 17380 6680 17436
rect 6680 17380 6684 17436
rect 6620 17376 6684 17380
rect 11808 17436 11872 17440
rect 11808 17380 11812 17436
rect 11812 17380 11868 17436
rect 11868 17380 11872 17436
rect 11808 17376 11872 17380
rect 11888 17436 11952 17440
rect 11888 17380 11892 17436
rect 11892 17380 11948 17436
rect 11948 17380 11952 17436
rect 11888 17376 11952 17380
rect 11968 17436 12032 17440
rect 11968 17380 11972 17436
rect 11972 17380 12028 17436
rect 12028 17380 12032 17436
rect 11968 17376 12032 17380
rect 12048 17436 12112 17440
rect 12048 17380 12052 17436
rect 12052 17380 12108 17436
rect 12108 17380 12112 17436
rect 12048 17376 12112 17380
rect 17236 17436 17300 17440
rect 17236 17380 17240 17436
rect 17240 17380 17296 17436
rect 17296 17380 17300 17436
rect 17236 17376 17300 17380
rect 17316 17436 17380 17440
rect 17316 17380 17320 17436
rect 17320 17380 17376 17436
rect 17376 17380 17380 17436
rect 17316 17376 17380 17380
rect 17396 17436 17460 17440
rect 17396 17380 17400 17436
rect 17400 17380 17456 17436
rect 17456 17380 17460 17436
rect 17396 17376 17460 17380
rect 17476 17436 17540 17440
rect 17476 17380 17480 17436
rect 17480 17380 17536 17436
rect 17536 17380 17540 17436
rect 17476 17376 17540 17380
rect 22664 17436 22728 17440
rect 22664 17380 22668 17436
rect 22668 17380 22724 17436
rect 22724 17380 22728 17436
rect 22664 17376 22728 17380
rect 22744 17436 22808 17440
rect 22744 17380 22748 17436
rect 22748 17380 22804 17436
rect 22804 17380 22808 17436
rect 22744 17376 22808 17380
rect 22824 17436 22888 17440
rect 22824 17380 22828 17436
rect 22828 17380 22884 17436
rect 22884 17380 22888 17436
rect 22824 17376 22888 17380
rect 22904 17436 22968 17440
rect 22904 17380 22908 17436
rect 22908 17380 22964 17436
rect 22964 17380 22968 17436
rect 22904 17376 22968 17380
rect 3666 16892 3730 16896
rect 3666 16836 3670 16892
rect 3670 16836 3726 16892
rect 3726 16836 3730 16892
rect 3666 16832 3730 16836
rect 3746 16892 3810 16896
rect 3746 16836 3750 16892
rect 3750 16836 3806 16892
rect 3806 16836 3810 16892
rect 3746 16832 3810 16836
rect 3826 16892 3890 16896
rect 3826 16836 3830 16892
rect 3830 16836 3886 16892
rect 3886 16836 3890 16892
rect 3826 16832 3890 16836
rect 3906 16892 3970 16896
rect 3906 16836 3910 16892
rect 3910 16836 3966 16892
rect 3966 16836 3970 16892
rect 3906 16832 3970 16836
rect 9094 16892 9158 16896
rect 9094 16836 9098 16892
rect 9098 16836 9154 16892
rect 9154 16836 9158 16892
rect 9094 16832 9158 16836
rect 9174 16892 9238 16896
rect 9174 16836 9178 16892
rect 9178 16836 9234 16892
rect 9234 16836 9238 16892
rect 9174 16832 9238 16836
rect 9254 16892 9318 16896
rect 9254 16836 9258 16892
rect 9258 16836 9314 16892
rect 9314 16836 9318 16892
rect 9254 16832 9318 16836
rect 9334 16892 9398 16896
rect 9334 16836 9338 16892
rect 9338 16836 9394 16892
rect 9394 16836 9398 16892
rect 9334 16832 9398 16836
rect 14522 16892 14586 16896
rect 14522 16836 14526 16892
rect 14526 16836 14582 16892
rect 14582 16836 14586 16892
rect 14522 16832 14586 16836
rect 14602 16892 14666 16896
rect 14602 16836 14606 16892
rect 14606 16836 14662 16892
rect 14662 16836 14666 16892
rect 14602 16832 14666 16836
rect 14682 16892 14746 16896
rect 14682 16836 14686 16892
rect 14686 16836 14742 16892
rect 14742 16836 14746 16892
rect 14682 16832 14746 16836
rect 14762 16892 14826 16896
rect 14762 16836 14766 16892
rect 14766 16836 14822 16892
rect 14822 16836 14826 16892
rect 14762 16832 14826 16836
rect 19950 16892 20014 16896
rect 19950 16836 19954 16892
rect 19954 16836 20010 16892
rect 20010 16836 20014 16892
rect 19950 16832 20014 16836
rect 20030 16892 20094 16896
rect 20030 16836 20034 16892
rect 20034 16836 20090 16892
rect 20090 16836 20094 16892
rect 20030 16832 20094 16836
rect 20110 16892 20174 16896
rect 20110 16836 20114 16892
rect 20114 16836 20170 16892
rect 20170 16836 20174 16892
rect 20110 16832 20174 16836
rect 20190 16892 20254 16896
rect 20190 16836 20194 16892
rect 20194 16836 20250 16892
rect 20250 16836 20254 16892
rect 20190 16832 20254 16836
rect 6380 16348 6444 16352
rect 6380 16292 6384 16348
rect 6384 16292 6440 16348
rect 6440 16292 6444 16348
rect 6380 16288 6444 16292
rect 6460 16348 6524 16352
rect 6460 16292 6464 16348
rect 6464 16292 6520 16348
rect 6520 16292 6524 16348
rect 6460 16288 6524 16292
rect 6540 16348 6604 16352
rect 6540 16292 6544 16348
rect 6544 16292 6600 16348
rect 6600 16292 6604 16348
rect 6540 16288 6604 16292
rect 6620 16348 6684 16352
rect 6620 16292 6624 16348
rect 6624 16292 6680 16348
rect 6680 16292 6684 16348
rect 6620 16288 6684 16292
rect 11808 16348 11872 16352
rect 11808 16292 11812 16348
rect 11812 16292 11868 16348
rect 11868 16292 11872 16348
rect 11808 16288 11872 16292
rect 11888 16348 11952 16352
rect 11888 16292 11892 16348
rect 11892 16292 11948 16348
rect 11948 16292 11952 16348
rect 11888 16288 11952 16292
rect 11968 16348 12032 16352
rect 11968 16292 11972 16348
rect 11972 16292 12028 16348
rect 12028 16292 12032 16348
rect 11968 16288 12032 16292
rect 12048 16348 12112 16352
rect 12048 16292 12052 16348
rect 12052 16292 12108 16348
rect 12108 16292 12112 16348
rect 12048 16288 12112 16292
rect 17236 16348 17300 16352
rect 17236 16292 17240 16348
rect 17240 16292 17296 16348
rect 17296 16292 17300 16348
rect 17236 16288 17300 16292
rect 17316 16348 17380 16352
rect 17316 16292 17320 16348
rect 17320 16292 17376 16348
rect 17376 16292 17380 16348
rect 17316 16288 17380 16292
rect 17396 16348 17460 16352
rect 17396 16292 17400 16348
rect 17400 16292 17456 16348
rect 17456 16292 17460 16348
rect 17396 16288 17460 16292
rect 17476 16348 17540 16352
rect 17476 16292 17480 16348
rect 17480 16292 17536 16348
rect 17536 16292 17540 16348
rect 17476 16288 17540 16292
rect 22664 16348 22728 16352
rect 22664 16292 22668 16348
rect 22668 16292 22724 16348
rect 22724 16292 22728 16348
rect 22664 16288 22728 16292
rect 22744 16348 22808 16352
rect 22744 16292 22748 16348
rect 22748 16292 22804 16348
rect 22804 16292 22808 16348
rect 22744 16288 22808 16292
rect 22824 16348 22888 16352
rect 22824 16292 22828 16348
rect 22828 16292 22884 16348
rect 22884 16292 22888 16348
rect 22824 16288 22888 16292
rect 22904 16348 22968 16352
rect 22904 16292 22908 16348
rect 22908 16292 22964 16348
rect 22964 16292 22968 16348
rect 22904 16288 22968 16292
rect 3666 15804 3730 15808
rect 3666 15748 3670 15804
rect 3670 15748 3726 15804
rect 3726 15748 3730 15804
rect 3666 15744 3730 15748
rect 3746 15804 3810 15808
rect 3746 15748 3750 15804
rect 3750 15748 3806 15804
rect 3806 15748 3810 15804
rect 3746 15744 3810 15748
rect 3826 15804 3890 15808
rect 3826 15748 3830 15804
rect 3830 15748 3886 15804
rect 3886 15748 3890 15804
rect 3826 15744 3890 15748
rect 3906 15804 3970 15808
rect 3906 15748 3910 15804
rect 3910 15748 3966 15804
rect 3966 15748 3970 15804
rect 3906 15744 3970 15748
rect 9094 15804 9158 15808
rect 9094 15748 9098 15804
rect 9098 15748 9154 15804
rect 9154 15748 9158 15804
rect 9094 15744 9158 15748
rect 9174 15804 9238 15808
rect 9174 15748 9178 15804
rect 9178 15748 9234 15804
rect 9234 15748 9238 15804
rect 9174 15744 9238 15748
rect 9254 15804 9318 15808
rect 9254 15748 9258 15804
rect 9258 15748 9314 15804
rect 9314 15748 9318 15804
rect 9254 15744 9318 15748
rect 9334 15804 9398 15808
rect 9334 15748 9338 15804
rect 9338 15748 9394 15804
rect 9394 15748 9398 15804
rect 9334 15744 9398 15748
rect 14522 15804 14586 15808
rect 14522 15748 14526 15804
rect 14526 15748 14582 15804
rect 14582 15748 14586 15804
rect 14522 15744 14586 15748
rect 14602 15804 14666 15808
rect 14602 15748 14606 15804
rect 14606 15748 14662 15804
rect 14662 15748 14666 15804
rect 14602 15744 14666 15748
rect 14682 15804 14746 15808
rect 14682 15748 14686 15804
rect 14686 15748 14742 15804
rect 14742 15748 14746 15804
rect 14682 15744 14746 15748
rect 14762 15804 14826 15808
rect 14762 15748 14766 15804
rect 14766 15748 14822 15804
rect 14822 15748 14826 15804
rect 14762 15744 14826 15748
rect 19950 15804 20014 15808
rect 19950 15748 19954 15804
rect 19954 15748 20010 15804
rect 20010 15748 20014 15804
rect 19950 15744 20014 15748
rect 20030 15804 20094 15808
rect 20030 15748 20034 15804
rect 20034 15748 20090 15804
rect 20090 15748 20094 15804
rect 20030 15744 20094 15748
rect 20110 15804 20174 15808
rect 20110 15748 20114 15804
rect 20114 15748 20170 15804
rect 20170 15748 20174 15804
rect 20110 15744 20174 15748
rect 20190 15804 20254 15808
rect 20190 15748 20194 15804
rect 20194 15748 20250 15804
rect 20250 15748 20254 15804
rect 20190 15744 20254 15748
rect 6380 15260 6444 15264
rect 6380 15204 6384 15260
rect 6384 15204 6440 15260
rect 6440 15204 6444 15260
rect 6380 15200 6444 15204
rect 6460 15260 6524 15264
rect 6460 15204 6464 15260
rect 6464 15204 6520 15260
rect 6520 15204 6524 15260
rect 6460 15200 6524 15204
rect 6540 15260 6604 15264
rect 6540 15204 6544 15260
rect 6544 15204 6600 15260
rect 6600 15204 6604 15260
rect 6540 15200 6604 15204
rect 6620 15260 6684 15264
rect 6620 15204 6624 15260
rect 6624 15204 6680 15260
rect 6680 15204 6684 15260
rect 6620 15200 6684 15204
rect 11808 15260 11872 15264
rect 11808 15204 11812 15260
rect 11812 15204 11868 15260
rect 11868 15204 11872 15260
rect 11808 15200 11872 15204
rect 11888 15260 11952 15264
rect 11888 15204 11892 15260
rect 11892 15204 11948 15260
rect 11948 15204 11952 15260
rect 11888 15200 11952 15204
rect 11968 15260 12032 15264
rect 11968 15204 11972 15260
rect 11972 15204 12028 15260
rect 12028 15204 12032 15260
rect 11968 15200 12032 15204
rect 12048 15260 12112 15264
rect 12048 15204 12052 15260
rect 12052 15204 12108 15260
rect 12108 15204 12112 15260
rect 12048 15200 12112 15204
rect 17236 15260 17300 15264
rect 17236 15204 17240 15260
rect 17240 15204 17296 15260
rect 17296 15204 17300 15260
rect 17236 15200 17300 15204
rect 17316 15260 17380 15264
rect 17316 15204 17320 15260
rect 17320 15204 17376 15260
rect 17376 15204 17380 15260
rect 17316 15200 17380 15204
rect 17396 15260 17460 15264
rect 17396 15204 17400 15260
rect 17400 15204 17456 15260
rect 17456 15204 17460 15260
rect 17396 15200 17460 15204
rect 17476 15260 17540 15264
rect 17476 15204 17480 15260
rect 17480 15204 17536 15260
rect 17536 15204 17540 15260
rect 17476 15200 17540 15204
rect 22664 15260 22728 15264
rect 22664 15204 22668 15260
rect 22668 15204 22724 15260
rect 22724 15204 22728 15260
rect 22664 15200 22728 15204
rect 22744 15260 22808 15264
rect 22744 15204 22748 15260
rect 22748 15204 22804 15260
rect 22804 15204 22808 15260
rect 22744 15200 22808 15204
rect 22824 15260 22888 15264
rect 22824 15204 22828 15260
rect 22828 15204 22884 15260
rect 22884 15204 22888 15260
rect 22824 15200 22888 15204
rect 22904 15260 22968 15264
rect 22904 15204 22908 15260
rect 22908 15204 22964 15260
rect 22964 15204 22968 15260
rect 22904 15200 22968 15204
rect 3666 14716 3730 14720
rect 3666 14660 3670 14716
rect 3670 14660 3726 14716
rect 3726 14660 3730 14716
rect 3666 14656 3730 14660
rect 3746 14716 3810 14720
rect 3746 14660 3750 14716
rect 3750 14660 3806 14716
rect 3806 14660 3810 14716
rect 3746 14656 3810 14660
rect 3826 14716 3890 14720
rect 3826 14660 3830 14716
rect 3830 14660 3886 14716
rect 3886 14660 3890 14716
rect 3826 14656 3890 14660
rect 3906 14716 3970 14720
rect 3906 14660 3910 14716
rect 3910 14660 3966 14716
rect 3966 14660 3970 14716
rect 3906 14656 3970 14660
rect 9094 14716 9158 14720
rect 9094 14660 9098 14716
rect 9098 14660 9154 14716
rect 9154 14660 9158 14716
rect 9094 14656 9158 14660
rect 9174 14716 9238 14720
rect 9174 14660 9178 14716
rect 9178 14660 9234 14716
rect 9234 14660 9238 14716
rect 9174 14656 9238 14660
rect 9254 14716 9318 14720
rect 9254 14660 9258 14716
rect 9258 14660 9314 14716
rect 9314 14660 9318 14716
rect 9254 14656 9318 14660
rect 9334 14716 9398 14720
rect 9334 14660 9338 14716
rect 9338 14660 9394 14716
rect 9394 14660 9398 14716
rect 9334 14656 9398 14660
rect 14522 14716 14586 14720
rect 14522 14660 14526 14716
rect 14526 14660 14582 14716
rect 14582 14660 14586 14716
rect 14522 14656 14586 14660
rect 14602 14716 14666 14720
rect 14602 14660 14606 14716
rect 14606 14660 14662 14716
rect 14662 14660 14666 14716
rect 14602 14656 14666 14660
rect 14682 14716 14746 14720
rect 14682 14660 14686 14716
rect 14686 14660 14742 14716
rect 14742 14660 14746 14716
rect 14682 14656 14746 14660
rect 14762 14716 14826 14720
rect 14762 14660 14766 14716
rect 14766 14660 14822 14716
rect 14822 14660 14826 14716
rect 14762 14656 14826 14660
rect 19950 14716 20014 14720
rect 19950 14660 19954 14716
rect 19954 14660 20010 14716
rect 20010 14660 20014 14716
rect 19950 14656 20014 14660
rect 20030 14716 20094 14720
rect 20030 14660 20034 14716
rect 20034 14660 20090 14716
rect 20090 14660 20094 14716
rect 20030 14656 20094 14660
rect 20110 14716 20174 14720
rect 20110 14660 20114 14716
rect 20114 14660 20170 14716
rect 20170 14660 20174 14716
rect 20110 14656 20174 14660
rect 20190 14716 20254 14720
rect 20190 14660 20194 14716
rect 20194 14660 20250 14716
rect 20250 14660 20254 14716
rect 20190 14656 20254 14660
rect 6380 14172 6444 14176
rect 6380 14116 6384 14172
rect 6384 14116 6440 14172
rect 6440 14116 6444 14172
rect 6380 14112 6444 14116
rect 6460 14172 6524 14176
rect 6460 14116 6464 14172
rect 6464 14116 6520 14172
rect 6520 14116 6524 14172
rect 6460 14112 6524 14116
rect 6540 14172 6604 14176
rect 6540 14116 6544 14172
rect 6544 14116 6600 14172
rect 6600 14116 6604 14172
rect 6540 14112 6604 14116
rect 6620 14172 6684 14176
rect 6620 14116 6624 14172
rect 6624 14116 6680 14172
rect 6680 14116 6684 14172
rect 6620 14112 6684 14116
rect 11808 14172 11872 14176
rect 11808 14116 11812 14172
rect 11812 14116 11868 14172
rect 11868 14116 11872 14172
rect 11808 14112 11872 14116
rect 11888 14172 11952 14176
rect 11888 14116 11892 14172
rect 11892 14116 11948 14172
rect 11948 14116 11952 14172
rect 11888 14112 11952 14116
rect 11968 14172 12032 14176
rect 11968 14116 11972 14172
rect 11972 14116 12028 14172
rect 12028 14116 12032 14172
rect 11968 14112 12032 14116
rect 12048 14172 12112 14176
rect 12048 14116 12052 14172
rect 12052 14116 12108 14172
rect 12108 14116 12112 14172
rect 12048 14112 12112 14116
rect 17236 14172 17300 14176
rect 17236 14116 17240 14172
rect 17240 14116 17296 14172
rect 17296 14116 17300 14172
rect 17236 14112 17300 14116
rect 17316 14172 17380 14176
rect 17316 14116 17320 14172
rect 17320 14116 17376 14172
rect 17376 14116 17380 14172
rect 17316 14112 17380 14116
rect 17396 14172 17460 14176
rect 17396 14116 17400 14172
rect 17400 14116 17456 14172
rect 17456 14116 17460 14172
rect 17396 14112 17460 14116
rect 17476 14172 17540 14176
rect 17476 14116 17480 14172
rect 17480 14116 17536 14172
rect 17536 14116 17540 14172
rect 17476 14112 17540 14116
rect 22664 14172 22728 14176
rect 22664 14116 22668 14172
rect 22668 14116 22724 14172
rect 22724 14116 22728 14172
rect 22664 14112 22728 14116
rect 22744 14172 22808 14176
rect 22744 14116 22748 14172
rect 22748 14116 22804 14172
rect 22804 14116 22808 14172
rect 22744 14112 22808 14116
rect 22824 14172 22888 14176
rect 22824 14116 22828 14172
rect 22828 14116 22884 14172
rect 22884 14116 22888 14172
rect 22824 14112 22888 14116
rect 22904 14172 22968 14176
rect 22904 14116 22908 14172
rect 22908 14116 22964 14172
rect 22964 14116 22968 14172
rect 22904 14112 22968 14116
rect 3666 13628 3730 13632
rect 3666 13572 3670 13628
rect 3670 13572 3726 13628
rect 3726 13572 3730 13628
rect 3666 13568 3730 13572
rect 3746 13628 3810 13632
rect 3746 13572 3750 13628
rect 3750 13572 3806 13628
rect 3806 13572 3810 13628
rect 3746 13568 3810 13572
rect 3826 13628 3890 13632
rect 3826 13572 3830 13628
rect 3830 13572 3886 13628
rect 3886 13572 3890 13628
rect 3826 13568 3890 13572
rect 3906 13628 3970 13632
rect 3906 13572 3910 13628
rect 3910 13572 3966 13628
rect 3966 13572 3970 13628
rect 3906 13568 3970 13572
rect 9094 13628 9158 13632
rect 9094 13572 9098 13628
rect 9098 13572 9154 13628
rect 9154 13572 9158 13628
rect 9094 13568 9158 13572
rect 9174 13628 9238 13632
rect 9174 13572 9178 13628
rect 9178 13572 9234 13628
rect 9234 13572 9238 13628
rect 9174 13568 9238 13572
rect 9254 13628 9318 13632
rect 9254 13572 9258 13628
rect 9258 13572 9314 13628
rect 9314 13572 9318 13628
rect 9254 13568 9318 13572
rect 9334 13628 9398 13632
rect 9334 13572 9338 13628
rect 9338 13572 9394 13628
rect 9394 13572 9398 13628
rect 9334 13568 9398 13572
rect 14522 13628 14586 13632
rect 14522 13572 14526 13628
rect 14526 13572 14582 13628
rect 14582 13572 14586 13628
rect 14522 13568 14586 13572
rect 14602 13628 14666 13632
rect 14602 13572 14606 13628
rect 14606 13572 14662 13628
rect 14662 13572 14666 13628
rect 14602 13568 14666 13572
rect 14682 13628 14746 13632
rect 14682 13572 14686 13628
rect 14686 13572 14742 13628
rect 14742 13572 14746 13628
rect 14682 13568 14746 13572
rect 14762 13628 14826 13632
rect 14762 13572 14766 13628
rect 14766 13572 14822 13628
rect 14822 13572 14826 13628
rect 14762 13568 14826 13572
rect 19950 13628 20014 13632
rect 19950 13572 19954 13628
rect 19954 13572 20010 13628
rect 20010 13572 20014 13628
rect 19950 13568 20014 13572
rect 20030 13628 20094 13632
rect 20030 13572 20034 13628
rect 20034 13572 20090 13628
rect 20090 13572 20094 13628
rect 20030 13568 20094 13572
rect 20110 13628 20174 13632
rect 20110 13572 20114 13628
rect 20114 13572 20170 13628
rect 20170 13572 20174 13628
rect 20110 13568 20174 13572
rect 20190 13628 20254 13632
rect 20190 13572 20194 13628
rect 20194 13572 20250 13628
rect 20250 13572 20254 13628
rect 20190 13568 20254 13572
rect 6380 13084 6444 13088
rect 6380 13028 6384 13084
rect 6384 13028 6440 13084
rect 6440 13028 6444 13084
rect 6380 13024 6444 13028
rect 6460 13084 6524 13088
rect 6460 13028 6464 13084
rect 6464 13028 6520 13084
rect 6520 13028 6524 13084
rect 6460 13024 6524 13028
rect 6540 13084 6604 13088
rect 6540 13028 6544 13084
rect 6544 13028 6600 13084
rect 6600 13028 6604 13084
rect 6540 13024 6604 13028
rect 6620 13084 6684 13088
rect 6620 13028 6624 13084
rect 6624 13028 6680 13084
rect 6680 13028 6684 13084
rect 6620 13024 6684 13028
rect 11808 13084 11872 13088
rect 11808 13028 11812 13084
rect 11812 13028 11868 13084
rect 11868 13028 11872 13084
rect 11808 13024 11872 13028
rect 11888 13084 11952 13088
rect 11888 13028 11892 13084
rect 11892 13028 11948 13084
rect 11948 13028 11952 13084
rect 11888 13024 11952 13028
rect 11968 13084 12032 13088
rect 11968 13028 11972 13084
rect 11972 13028 12028 13084
rect 12028 13028 12032 13084
rect 11968 13024 12032 13028
rect 12048 13084 12112 13088
rect 12048 13028 12052 13084
rect 12052 13028 12108 13084
rect 12108 13028 12112 13084
rect 12048 13024 12112 13028
rect 17236 13084 17300 13088
rect 17236 13028 17240 13084
rect 17240 13028 17296 13084
rect 17296 13028 17300 13084
rect 17236 13024 17300 13028
rect 17316 13084 17380 13088
rect 17316 13028 17320 13084
rect 17320 13028 17376 13084
rect 17376 13028 17380 13084
rect 17316 13024 17380 13028
rect 17396 13084 17460 13088
rect 17396 13028 17400 13084
rect 17400 13028 17456 13084
rect 17456 13028 17460 13084
rect 17396 13024 17460 13028
rect 17476 13084 17540 13088
rect 17476 13028 17480 13084
rect 17480 13028 17536 13084
rect 17536 13028 17540 13084
rect 17476 13024 17540 13028
rect 22664 13084 22728 13088
rect 22664 13028 22668 13084
rect 22668 13028 22724 13084
rect 22724 13028 22728 13084
rect 22664 13024 22728 13028
rect 22744 13084 22808 13088
rect 22744 13028 22748 13084
rect 22748 13028 22804 13084
rect 22804 13028 22808 13084
rect 22744 13024 22808 13028
rect 22824 13084 22888 13088
rect 22824 13028 22828 13084
rect 22828 13028 22884 13084
rect 22884 13028 22888 13084
rect 22824 13024 22888 13028
rect 22904 13084 22968 13088
rect 22904 13028 22908 13084
rect 22908 13028 22964 13084
rect 22964 13028 22968 13084
rect 22904 13024 22968 13028
rect 3666 12540 3730 12544
rect 3666 12484 3670 12540
rect 3670 12484 3726 12540
rect 3726 12484 3730 12540
rect 3666 12480 3730 12484
rect 3746 12540 3810 12544
rect 3746 12484 3750 12540
rect 3750 12484 3806 12540
rect 3806 12484 3810 12540
rect 3746 12480 3810 12484
rect 3826 12540 3890 12544
rect 3826 12484 3830 12540
rect 3830 12484 3886 12540
rect 3886 12484 3890 12540
rect 3826 12480 3890 12484
rect 3906 12540 3970 12544
rect 3906 12484 3910 12540
rect 3910 12484 3966 12540
rect 3966 12484 3970 12540
rect 3906 12480 3970 12484
rect 9094 12540 9158 12544
rect 9094 12484 9098 12540
rect 9098 12484 9154 12540
rect 9154 12484 9158 12540
rect 9094 12480 9158 12484
rect 9174 12540 9238 12544
rect 9174 12484 9178 12540
rect 9178 12484 9234 12540
rect 9234 12484 9238 12540
rect 9174 12480 9238 12484
rect 9254 12540 9318 12544
rect 9254 12484 9258 12540
rect 9258 12484 9314 12540
rect 9314 12484 9318 12540
rect 9254 12480 9318 12484
rect 9334 12540 9398 12544
rect 9334 12484 9338 12540
rect 9338 12484 9394 12540
rect 9394 12484 9398 12540
rect 9334 12480 9398 12484
rect 14522 12540 14586 12544
rect 14522 12484 14526 12540
rect 14526 12484 14582 12540
rect 14582 12484 14586 12540
rect 14522 12480 14586 12484
rect 14602 12540 14666 12544
rect 14602 12484 14606 12540
rect 14606 12484 14662 12540
rect 14662 12484 14666 12540
rect 14602 12480 14666 12484
rect 14682 12540 14746 12544
rect 14682 12484 14686 12540
rect 14686 12484 14742 12540
rect 14742 12484 14746 12540
rect 14682 12480 14746 12484
rect 14762 12540 14826 12544
rect 14762 12484 14766 12540
rect 14766 12484 14822 12540
rect 14822 12484 14826 12540
rect 14762 12480 14826 12484
rect 19950 12540 20014 12544
rect 19950 12484 19954 12540
rect 19954 12484 20010 12540
rect 20010 12484 20014 12540
rect 19950 12480 20014 12484
rect 20030 12540 20094 12544
rect 20030 12484 20034 12540
rect 20034 12484 20090 12540
rect 20090 12484 20094 12540
rect 20030 12480 20094 12484
rect 20110 12540 20174 12544
rect 20110 12484 20114 12540
rect 20114 12484 20170 12540
rect 20170 12484 20174 12540
rect 20110 12480 20174 12484
rect 20190 12540 20254 12544
rect 20190 12484 20194 12540
rect 20194 12484 20250 12540
rect 20250 12484 20254 12540
rect 20190 12480 20254 12484
rect 6380 11996 6444 12000
rect 6380 11940 6384 11996
rect 6384 11940 6440 11996
rect 6440 11940 6444 11996
rect 6380 11936 6444 11940
rect 6460 11996 6524 12000
rect 6460 11940 6464 11996
rect 6464 11940 6520 11996
rect 6520 11940 6524 11996
rect 6460 11936 6524 11940
rect 6540 11996 6604 12000
rect 6540 11940 6544 11996
rect 6544 11940 6600 11996
rect 6600 11940 6604 11996
rect 6540 11936 6604 11940
rect 6620 11996 6684 12000
rect 6620 11940 6624 11996
rect 6624 11940 6680 11996
rect 6680 11940 6684 11996
rect 6620 11936 6684 11940
rect 11808 11996 11872 12000
rect 11808 11940 11812 11996
rect 11812 11940 11868 11996
rect 11868 11940 11872 11996
rect 11808 11936 11872 11940
rect 11888 11996 11952 12000
rect 11888 11940 11892 11996
rect 11892 11940 11948 11996
rect 11948 11940 11952 11996
rect 11888 11936 11952 11940
rect 11968 11996 12032 12000
rect 11968 11940 11972 11996
rect 11972 11940 12028 11996
rect 12028 11940 12032 11996
rect 11968 11936 12032 11940
rect 12048 11996 12112 12000
rect 12048 11940 12052 11996
rect 12052 11940 12108 11996
rect 12108 11940 12112 11996
rect 12048 11936 12112 11940
rect 17236 11996 17300 12000
rect 17236 11940 17240 11996
rect 17240 11940 17296 11996
rect 17296 11940 17300 11996
rect 17236 11936 17300 11940
rect 17316 11996 17380 12000
rect 17316 11940 17320 11996
rect 17320 11940 17376 11996
rect 17376 11940 17380 11996
rect 17316 11936 17380 11940
rect 17396 11996 17460 12000
rect 17396 11940 17400 11996
rect 17400 11940 17456 11996
rect 17456 11940 17460 11996
rect 17396 11936 17460 11940
rect 17476 11996 17540 12000
rect 17476 11940 17480 11996
rect 17480 11940 17536 11996
rect 17536 11940 17540 11996
rect 17476 11936 17540 11940
rect 22664 11996 22728 12000
rect 22664 11940 22668 11996
rect 22668 11940 22724 11996
rect 22724 11940 22728 11996
rect 22664 11936 22728 11940
rect 22744 11996 22808 12000
rect 22744 11940 22748 11996
rect 22748 11940 22804 11996
rect 22804 11940 22808 11996
rect 22744 11936 22808 11940
rect 22824 11996 22888 12000
rect 22824 11940 22828 11996
rect 22828 11940 22884 11996
rect 22884 11940 22888 11996
rect 22824 11936 22888 11940
rect 22904 11996 22968 12000
rect 22904 11940 22908 11996
rect 22908 11940 22964 11996
rect 22964 11940 22968 11996
rect 22904 11936 22968 11940
rect 3666 11452 3730 11456
rect 3666 11396 3670 11452
rect 3670 11396 3726 11452
rect 3726 11396 3730 11452
rect 3666 11392 3730 11396
rect 3746 11452 3810 11456
rect 3746 11396 3750 11452
rect 3750 11396 3806 11452
rect 3806 11396 3810 11452
rect 3746 11392 3810 11396
rect 3826 11452 3890 11456
rect 3826 11396 3830 11452
rect 3830 11396 3886 11452
rect 3886 11396 3890 11452
rect 3826 11392 3890 11396
rect 3906 11452 3970 11456
rect 3906 11396 3910 11452
rect 3910 11396 3966 11452
rect 3966 11396 3970 11452
rect 3906 11392 3970 11396
rect 9094 11452 9158 11456
rect 9094 11396 9098 11452
rect 9098 11396 9154 11452
rect 9154 11396 9158 11452
rect 9094 11392 9158 11396
rect 9174 11452 9238 11456
rect 9174 11396 9178 11452
rect 9178 11396 9234 11452
rect 9234 11396 9238 11452
rect 9174 11392 9238 11396
rect 9254 11452 9318 11456
rect 9254 11396 9258 11452
rect 9258 11396 9314 11452
rect 9314 11396 9318 11452
rect 9254 11392 9318 11396
rect 9334 11452 9398 11456
rect 9334 11396 9338 11452
rect 9338 11396 9394 11452
rect 9394 11396 9398 11452
rect 9334 11392 9398 11396
rect 14522 11452 14586 11456
rect 14522 11396 14526 11452
rect 14526 11396 14582 11452
rect 14582 11396 14586 11452
rect 14522 11392 14586 11396
rect 14602 11452 14666 11456
rect 14602 11396 14606 11452
rect 14606 11396 14662 11452
rect 14662 11396 14666 11452
rect 14602 11392 14666 11396
rect 14682 11452 14746 11456
rect 14682 11396 14686 11452
rect 14686 11396 14742 11452
rect 14742 11396 14746 11452
rect 14682 11392 14746 11396
rect 14762 11452 14826 11456
rect 14762 11396 14766 11452
rect 14766 11396 14822 11452
rect 14822 11396 14826 11452
rect 14762 11392 14826 11396
rect 19950 11452 20014 11456
rect 19950 11396 19954 11452
rect 19954 11396 20010 11452
rect 20010 11396 20014 11452
rect 19950 11392 20014 11396
rect 20030 11452 20094 11456
rect 20030 11396 20034 11452
rect 20034 11396 20090 11452
rect 20090 11396 20094 11452
rect 20030 11392 20094 11396
rect 20110 11452 20174 11456
rect 20110 11396 20114 11452
rect 20114 11396 20170 11452
rect 20170 11396 20174 11452
rect 20110 11392 20174 11396
rect 20190 11452 20254 11456
rect 20190 11396 20194 11452
rect 20194 11396 20250 11452
rect 20250 11396 20254 11452
rect 20190 11392 20254 11396
rect 15148 11052 15212 11116
rect 6380 10908 6444 10912
rect 6380 10852 6384 10908
rect 6384 10852 6440 10908
rect 6440 10852 6444 10908
rect 6380 10848 6444 10852
rect 6460 10908 6524 10912
rect 6460 10852 6464 10908
rect 6464 10852 6520 10908
rect 6520 10852 6524 10908
rect 6460 10848 6524 10852
rect 6540 10908 6604 10912
rect 6540 10852 6544 10908
rect 6544 10852 6600 10908
rect 6600 10852 6604 10908
rect 6540 10848 6604 10852
rect 6620 10908 6684 10912
rect 6620 10852 6624 10908
rect 6624 10852 6680 10908
rect 6680 10852 6684 10908
rect 6620 10848 6684 10852
rect 11808 10908 11872 10912
rect 11808 10852 11812 10908
rect 11812 10852 11868 10908
rect 11868 10852 11872 10908
rect 11808 10848 11872 10852
rect 11888 10908 11952 10912
rect 11888 10852 11892 10908
rect 11892 10852 11948 10908
rect 11948 10852 11952 10908
rect 11888 10848 11952 10852
rect 11968 10908 12032 10912
rect 11968 10852 11972 10908
rect 11972 10852 12028 10908
rect 12028 10852 12032 10908
rect 11968 10848 12032 10852
rect 12048 10908 12112 10912
rect 12048 10852 12052 10908
rect 12052 10852 12108 10908
rect 12108 10852 12112 10908
rect 12048 10848 12112 10852
rect 17236 10908 17300 10912
rect 17236 10852 17240 10908
rect 17240 10852 17296 10908
rect 17296 10852 17300 10908
rect 17236 10848 17300 10852
rect 17316 10908 17380 10912
rect 17316 10852 17320 10908
rect 17320 10852 17376 10908
rect 17376 10852 17380 10908
rect 17316 10848 17380 10852
rect 17396 10908 17460 10912
rect 17396 10852 17400 10908
rect 17400 10852 17456 10908
rect 17456 10852 17460 10908
rect 17396 10848 17460 10852
rect 17476 10908 17540 10912
rect 17476 10852 17480 10908
rect 17480 10852 17536 10908
rect 17536 10852 17540 10908
rect 17476 10848 17540 10852
rect 22664 10908 22728 10912
rect 22664 10852 22668 10908
rect 22668 10852 22724 10908
rect 22724 10852 22728 10908
rect 22664 10848 22728 10852
rect 22744 10908 22808 10912
rect 22744 10852 22748 10908
rect 22748 10852 22804 10908
rect 22804 10852 22808 10908
rect 22744 10848 22808 10852
rect 22824 10908 22888 10912
rect 22824 10852 22828 10908
rect 22828 10852 22884 10908
rect 22884 10852 22888 10908
rect 22824 10848 22888 10852
rect 22904 10908 22968 10912
rect 22904 10852 22908 10908
rect 22908 10852 22964 10908
rect 22964 10852 22968 10908
rect 22904 10848 22968 10852
rect 3666 10364 3730 10368
rect 3666 10308 3670 10364
rect 3670 10308 3726 10364
rect 3726 10308 3730 10364
rect 3666 10304 3730 10308
rect 3746 10364 3810 10368
rect 3746 10308 3750 10364
rect 3750 10308 3806 10364
rect 3806 10308 3810 10364
rect 3746 10304 3810 10308
rect 3826 10364 3890 10368
rect 3826 10308 3830 10364
rect 3830 10308 3886 10364
rect 3886 10308 3890 10364
rect 3826 10304 3890 10308
rect 3906 10364 3970 10368
rect 3906 10308 3910 10364
rect 3910 10308 3966 10364
rect 3966 10308 3970 10364
rect 3906 10304 3970 10308
rect 9094 10364 9158 10368
rect 9094 10308 9098 10364
rect 9098 10308 9154 10364
rect 9154 10308 9158 10364
rect 9094 10304 9158 10308
rect 9174 10364 9238 10368
rect 9174 10308 9178 10364
rect 9178 10308 9234 10364
rect 9234 10308 9238 10364
rect 9174 10304 9238 10308
rect 9254 10364 9318 10368
rect 9254 10308 9258 10364
rect 9258 10308 9314 10364
rect 9314 10308 9318 10364
rect 9254 10304 9318 10308
rect 9334 10364 9398 10368
rect 9334 10308 9338 10364
rect 9338 10308 9394 10364
rect 9394 10308 9398 10364
rect 9334 10304 9398 10308
rect 14522 10364 14586 10368
rect 14522 10308 14526 10364
rect 14526 10308 14582 10364
rect 14582 10308 14586 10364
rect 14522 10304 14586 10308
rect 14602 10364 14666 10368
rect 14602 10308 14606 10364
rect 14606 10308 14662 10364
rect 14662 10308 14666 10364
rect 14602 10304 14666 10308
rect 14682 10364 14746 10368
rect 14682 10308 14686 10364
rect 14686 10308 14742 10364
rect 14742 10308 14746 10364
rect 14682 10304 14746 10308
rect 14762 10364 14826 10368
rect 14762 10308 14766 10364
rect 14766 10308 14822 10364
rect 14822 10308 14826 10364
rect 14762 10304 14826 10308
rect 19950 10364 20014 10368
rect 19950 10308 19954 10364
rect 19954 10308 20010 10364
rect 20010 10308 20014 10364
rect 19950 10304 20014 10308
rect 20030 10364 20094 10368
rect 20030 10308 20034 10364
rect 20034 10308 20090 10364
rect 20090 10308 20094 10364
rect 20030 10304 20094 10308
rect 20110 10364 20174 10368
rect 20110 10308 20114 10364
rect 20114 10308 20170 10364
rect 20170 10308 20174 10364
rect 20110 10304 20174 10308
rect 20190 10364 20254 10368
rect 20190 10308 20194 10364
rect 20194 10308 20250 10364
rect 20250 10308 20254 10364
rect 20190 10304 20254 10308
rect 6380 9820 6444 9824
rect 6380 9764 6384 9820
rect 6384 9764 6440 9820
rect 6440 9764 6444 9820
rect 6380 9760 6444 9764
rect 6460 9820 6524 9824
rect 6460 9764 6464 9820
rect 6464 9764 6520 9820
rect 6520 9764 6524 9820
rect 6460 9760 6524 9764
rect 6540 9820 6604 9824
rect 6540 9764 6544 9820
rect 6544 9764 6600 9820
rect 6600 9764 6604 9820
rect 6540 9760 6604 9764
rect 6620 9820 6684 9824
rect 6620 9764 6624 9820
rect 6624 9764 6680 9820
rect 6680 9764 6684 9820
rect 6620 9760 6684 9764
rect 11808 9820 11872 9824
rect 11808 9764 11812 9820
rect 11812 9764 11868 9820
rect 11868 9764 11872 9820
rect 11808 9760 11872 9764
rect 11888 9820 11952 9824
rect 11888 9764 11892 9820
rect 11892 9764 11948 9820
rect 11948 9764 11952 9820
rect 11888 9760 11952 9764
rect 11968 9820 12032 9824
rect 11968 9764 11972 9820
rect 11972 9764 12028 9820
rect 12028 9764 12032 9820
rect 11968 9760 12032 9764
rect 12048 9820 12112 9824
rect 12048 9764 12052 9820
rect 12052 9764 12108 9820
rect 12108 9764 12112 9820
rect 12048 9760 12112 9764
rect 17236 9820 17300 9824
rect 17236 9764 17240 9820
rect 17240 9764 17296 9820
rect 17296 9764 17300 9820
rect 17236 9760 17300 9764
rect 17316 9820 17380 9824
rect 17316 9764 17320 9820
rect 17320 9764 17376 9820
rect 17376 9764 17380 9820
rect 17316 9760 17380 9764
rect 17396 9820 17460 9824
rect 17396 9764 17400 9820
rect 17400 9764 17456 9820
rect 17456 9764 17460 9820
rect 17396 9760 17460 9764
rect 17476 9820 17540 9824
rect 17476 9764 17480 9820
rect 17480 9764 17536 9820
rect 17536 9764 17540 9820
rect 17476 9760 17540 9764
rect 22664 9820 22728 9824
rect 22664 9764 22668 9820
rect 22668 9764 22724 9820
rect 22724 9764 22728 9820
rect 22664 9760 22728 9764
rect 22744 9820 22808 9824
rect 22744 9764 22748 9820
rect 22748 9764 22804 9820
rect 22804 9764 22808 9820
rect 22744 9760 22808 9764
rect 22824 9820 22888 9824
rect 22824 9764 22828 9820
rect 22828 9764 22884 9820
rect 22884 9764 22888 9820
rect 22824 9760 22888 9764
rect 22904 9820 22968 9824
rect 22904 9764 22908 9820
rect 22908 9764 22964 9820
rect 22964 9764 22968 9820
rect 22904 9760 22968 9764
rect 3666 9276 3730 9280
rect 3666 9220 3670 9276
rect 3670 9220 3726 9276
rect 3726 9220 3730 9276
rect 3666 9216 3730 9220
rect 3746 9276 3810 9280
rect 3746 9220 3750 9276
rect 3750 9220 3806 9276
rect 3806 9220 3810 9276
rect 3746 9216 3810 9220
rect 3826 9276 3890 9280
rect 3826 9220 3830 9276
rect 3830 9220 3886 9276
rect 3886 9220 3890 9276
rect 3826 9216 3890 9220
rect 3906 9276 3970 9280
rect 3906 9220 3910 9276
rect 3910 9220 3966 9276
rect 3966 9220 3970 9276
rect 3906 9216 3970 9220
rect 9094 9276 9158 9280
rect 9094 9220 9098 9276
rect 9098 9220 9154 9276
rect 9154 9220 9158 9276
rect 9094 9216 9158 9220
rect 9174 9276 9238 9280
rect 9174 9220 9178 9276
rect 9178 9220 9234 9276
rect 9234 9220 9238 9276
rect 9174 9216 9238 9220
rect 9254 9276 9318 9280
rect 9254 9220 9258 9276
rect 9258 9220 9314 9276
rect 9314 9220 9318 9276
rect 9254 9216 9318 9220
rect 9334 9276 9398 9280
rect 9334 9220 9338 9276
rect 9338 9220 9394 9276
rect 9394 9220 9398 9276
rect 9334 9216 9398 9220
rect 14522 9276 14586 9280
rect 14522 9220 14526 9276
rect 14526 9220 14582 9276
rect 14582 9220 14586 9276
rect 14522 9216 14586 9220
rect 14602 9276 14666 9280
rect 14602 9220 14606 9276
rect 14606 9220 14662 9276
rect 14662 9220 14666 9276
rect 14602 9216 14666 9220
rect 14682 9276 14746 9280
rect 14682 9220 14686 9276
rect 14686 9220 14742 9276
rect 14742 9220 14746 9276
rect 14682 9216 14746 9220
rect 14762 9276 14826 9280
rect 14762 9220 14766 9276
rect 14766 9220 14822 9276
rect 14822 9220 14826 9276
rect 14762 9216 14826 9220
rect 19950 9276 20014 9280
rect 19950 9220 19954 9276
rect 19954 9220 20010 9276
rect 20010 9220 20014 9276
rect 19950 9216 20014 9220
rect 20030 9276 20094 9280
rect 20030 9220 20034 9276
rect 20034 9220 20090 9276
rect 20090 9220 20094 9276
rect 20030 9216 20094 9220
rect 20110 9276 20174 9280
rect 20110 9220 20114 9276
rect 20114 9220 20170 9276
rect 20170 9220 20174 9276
rect 20110 9216 20174 9220
rect 20190 9276 20254 9280
rect 20190 9220 20194 9276
rect 20194 9220 20250 9276
rect 20250 9220 20254 9276
rect 20190 9216 20254 9220
rect 6380 8732 6444 8736
rect 6380 8676 6384 8732
rect 6384 8676 6440 8732
rect 6440 8676 6444 8732
rect 6380 8672 6444 8676
rect 6460 8732 6524 8736
rect 6460 8676 6464 8732
rect 6464 8676 6520 8732
rect 6520 8676 6524 8732
rect 6460 8672 6524 8676
rect 6540 8732 6604 8736
rect 6540 8676 6544 8732
rect 6544 8676 6600 8732
rect 6600 8676 6604 8732
rect 6540 8672 6604 8676
rect 6620 8732 6684 8736
rect 6620 8676 6624 8732
rect 6624 8676 6680 8732
rect 6680 8676 6684 8732
rect 6620 8672 6684 8676
rect 11808 8732 11872 8736
rect 11808 8676 11812 8732
rect 11812 8676 11868 8732
rect 11868 8676 11872 8732
rect 11808 8672 11872 8676
rect 11888 8732 11952 8736
rect 11888 8676 11892 8732
rect 11892 8676 11948 8732
rect 11948 8676 11952 8732
rect 11888 8672 11952 8676
rect 11968 8732 12032 8736
rect 11968 8676 11972 8732
rect 11972 8676 12028 8732
rect 12028 8676 12032 8732
rect 11968 8672 12032 8676
rect 12048 8732 12112 8736
rect 12048 8676 12052 8732
rect 12052 8676 12108 8732
rect 12108 8676 12112 8732
rect 12048 8672 12112 8676
rect 17236 8732 17300 8736
rect 17236 8676 17240 8732
rect 17240 8676 17296 8732
rect 17296 8676 17300 8732
rect 17236 8672 17300 8676
rect 17316 8732 17380 8736
rect 17316 8676 17320 8732
rect 17320 8676 17376 8732
rect 17376 8676 17380 8732
rect 17316 8672 17380 8676
rect 17396 8732 17460 8736
rect 17396 8676 17400 8732
rect 17400 8676 17456 8732
rect 17456 8676 17460 8732
rect 17396 8672 17460 8676
rect 17476 8732 17540 8736
rect 17476 8676 17480 8732
rect 17480 8676 17536 8732
rect 17536 8676 17540 8732
rect 17476 8672 17540 8676
rect 22664 8732 22728 8736
rect 22664 8676 22668 8732
rect 22668 8676 22724 8732
rect 22724 8676 22728 8732
rect 22664 8672 22728 8676
rect 22744 8732 22808 8736
rect 22744 8676 22748 8732
rect 22748 8676 22804 8732
rect 22804 8676 22808 8732
rect 22744 8672 22808 8676
rect 22824 8732 22888 8736
rect 22824 8676 22828 8732
rect 22828 8676 22884 8732
rect 22884 8676 22888 8732
rect 22824 8672 22888 8676
rect 22904 8732 22968 8736
rect 22904 8676 22908 8732
rect 22908 8676 22964 8732
rect 22964 8676 22968 8732
rect 22904 8672 22968 8676
rect 3666 8188 3730 8192
rect 3666 8132 3670 8188
rect 3670 8132 3726 8188
rect 3726 8132 3730 8188
rect 3666 8128 3730 8132
rect 3746 8188 3810 8192
rect 3746 8132 3750 8188
rect 3750 8132 3806 8188
rect 3806 8132 3810 8188
rect 3746 8128 3810 8132
rect 3826 8188 3890 8192
rect 3826 8132 3830 8188
rect 3830 8132 3886 8188
rect 3886 8132 3890 8188
rect 3826 8128 3890 8132
rect 3906 8188 3970 8192
rect 3906 8132 3910 8188
rect 3910 8132 3966 8188
rect 3966 8132 3970 8188
rect 3906 8128 3970 8132
rect 9094 8188 9158 8192
rect 9094 8132 9098 8188
rect 9098 8132 9154 8188
rect 9154 8132 9158 8188
rect 9094 8128 9158 8132
rect 9174 8188 9238 8192
rect 9174 8132 9178 8188
rect 9178 8132 9234 8188
rect 9234 8132 9238 8188
rect 9174 8128 9238 8132
rect 9254 8188 9318 8192
rect 9254 8132 9258 8188
rect 9258 8132 9314 8188
rect 9314 8132 9318 8188
rect 9254 8128 9318 8132
rect 9334 8188 9398 8192
rect 9334 8132 9338 8188
rect 9338 8132 9394 8188
rect 9394 8132 9398 8188
rect 9334 8128 9398 8132
rect 14522 8188 14586 8192
rect 14522 8132 14526 8188
rect 14526 8132 14582 8188
rect 14582 8132 14586 8188
rect 14522 8128 14586 8132
rect 14602 8188 14666 8192
rect 14602 8132 14606 8188
rect 14606 8132 14662 8188
rect 14662 8132 14666 8188
rect 14602 8128 14666 8132
rect 14682 8188 14746 8192
rect 14682 8132 14686 8188
rect 14686 8132 14742 8188
rect 14742 8132 14746 8188
rect 14682 8128 14746 8132
rect 14762 8188 14826 8192
rect 14762 8132 14766 8188
rect 14766 8132 14822 8188
rect 14822 8132 14826 8188
rect 14762 8128 14826 8132
rect 19950 8188 20014 8192
rect 19950 8132 19954 8188
rect 19954 8132 20010 8188
rect 20010 8132 20014 8188
rect 19950 8128 20014 8132
rect 20030 8188 20094 8192
rect 20030 8132 20034 8188
rect 20034 8132 20090 8188
rect 20090 8132 20094 8188
rect 20030 8128 20094 8132
rect 20110 8188 20174 8192
rect 20110 8132 20114 8188
rect 20114 8132 20170 8188
rect 20170 8132 20174 8188
rect 20110 8128 20174 8132
rect 20190 8188 20254 8192
rect 20190 8132 20194 8188
rect 20194 8132 20250 8188
rect 20250 8132 20254 8188
rect 20190 8128 20254 8132
rect 6380 7644 6444 7648
rect 6380 7588 6384 7644
rect 6384 7588 6440 7644
rect 6440 7588 6444 7644
rect 6380 7584 6444 7588
rect 6460 7644 6524 7648
rect 6460 7588 6464 7644
rect 6464 7588 6520 7644
rect 6520 7588 6524 7644
rect 6460 7584 6524 7588
rect 6540 7644 6604 7648
rect 6540 7588 6544 7644
rect 6544 7588 6600 7644
rect 6600 7588 6604 7644
rect 6540 7584 6604 7588
rect 6620 7644 6684 7648
rect 6620 7588 6624 7644
rect 6624 7588 6680 7644
rect 6680 7588 6684 7644
rect 6620 7584 6684 7588
rect 11808 7644 11872 7648
rect 11808 7588 11812 7644
rect 11812 7588 11868 7644
rect 11868 7588 11872 7644
rect 11808 7584 11872 7588
rect 11888 7644 11952 7648
rect 11888 7588 11892 7644
rect 11892 7588 11948 7644
rect 11948 7588 11952 7644
rect 11888 7584 11952 7588
rect 11968 7644 12032 7648
rect 11968 7588 11972 7644
rect 11972 7588 12028 7644
rect 12028 7588 12032 7644
rect 11968 7584 12032 7588
rect 12048 7644 12112 7648
rect 12048 7588 12052 7644
rect 12052 7588 12108 7644
rect 12108 7588 12112 7644
rect 12048 7584 12112 7588
rect 17236 7644 17300 7648
rect 17236 7588 17240 7644
rect 17240 7588 17296 7644
rect 17296 7588 17300 7644
rect 17236 7584 17300 7588
rect 17316 7644 17380 7648
rect 17316 7588 17320 7644
rect 17320 7588 17376 7644
rect 17376 7588 17380 7644
rect 17316 7584 17380 7588
rect 17396 7644 17460 7648
rect 17396 7588 17400 7644
rect 17400 7588 17456 7644
rect 17456 7588 17460 7644
rect 17396 7584 17460 7588
rect 17476 7644 17540 7648
rect 17476 7588 17480 7644
rect 17480 7588 17536 7644
rect 17536 7588 17540 7644
rect 17476 7584 17540 7588
rect 22664 7644 22728 7648
rect 22664 7588 22668 7644
rect 22668 7588 22724 7644
rect 22724 7588 22728 7644
rect 22664 7584 22728 7588
rect 22744 7644 22808 7648
rect 22744 7588 22748 7644
rect 22748 7588 22804 7644
rect 22804 7588 22808 7644
rect 22744 7584 22808 7588
rect 22824 7644 22888 7648
rect 22824 7588 22828 7644
rect 22828 7588 22884 7644
rect 22884 7588 22888 7644
rect 22824 7584 22888 7588
rect 22904 7644 22968 7648
rect 22904 7588 22908 7644
rect 22908 7588 22964 7644
rect 22964 7588 22968 7644
rect 22904 7584 22968 7588
rect 15148 7380 15212 7444
rect 3666 7100 3730 7104
rect 3666 7044 3670 7100
rect 3670 7044 3726 7100
rect 3726 7044 3730 7100
rect 3666 7040 3730 7044
rect 3746 7100 3810 7104
rect 3746 7044 3750 7100
rect 3750 7044 3806 7100
rect 3806 7044 3810 7100
rect 3746 7040 3810 7044
rect 3826 7100 3890 7104
rect 3826 7044 3830 7100
rect 3830 7044 3886 7100
rect 3886 7044 3890 7100
rect 3826 7040 3890 7044
rect 3906 7100 3970 7104
rect 3906 7044 3910 7100
rect 3910 7044 3966 7100
rect 3966 7044 3970 7100
rect 3906 7040 3970 7044
rect 9094 7100 9158 7104
rect 9094 7044 9098 7100
rect 9098 7044 9154 7100
rect 9154 7044 9158 7100
rect 9094 7040 9158 7044
rect 9174 7100 9238 7104
rect 9174 7044 9178 7100
rect 9178 7044 9234 7100
rect 9234 7044 9238 7100
rect 9174 7040 9238 7044
rect 9254 7100 9318 7104
rect 9254 7044 9258 7100
rect 9258 7044 9314 7100
rect 9314 7044 9318 7100
rect 9254 7040 9318 7044
rect 9334 7100 9398 7104
rect 9334 7044 9338 7100
rect 9338 7044 9394 7100
rect 9394 7044 9398 7100
rect 9334 7040 9398 7044
rect 14522 7100 14586 7104
rect 14522 7044 14526 7100
rect 14526 7044 14582 7100
rect 14582 7044 14586 7100
rect 14522 7040 14586 7044
rect 14602 7100 14666 7104
rect 14602 7044 14606 7100
rect 14606 7044 14662 7100
rect 14662 7044 14666 7100
rect 14602 7040 14666 7044
rect 14682 7100 14746 7104
rect 14682 7044 14686 7100
rect 14686 7044 14742 7100
rect 14742 7044 14746 7100
rect 14682 7040 14746 7044
rect 14762 7100 14826 7104
rect 14762 7044 14766 7100
rect 14766 7044 14822 7100
rect 14822 7044 14826 7100
rect 14762 7040 14826 7044
rect 19950 7100 20014 7104
rect 19950 7044 19954 7100
rect 19954 7044 20010 7100
rect 20010 7044 20014 7100
rect 19950 7040 20014 7044
rect 20030 7100 20094 7104
rect 20030 7044 20034 7100
rect 20034 7044 20090 7100
rect 20090 7044 20094 7100
rect 20030 7040 20094 7044
rect 20110 7100 20174 7104
rect 20110 7044 20114 7100
rect 20114 7044 20170 7100
rect 20170 7044 20174 7100
rect 20110 7040 20174 7044
rect 20190 7100 20254 7104
rect 20190 7044 20194 7100
rect 20194 7044 20250 7100
rect 20250 7044 20254 7100
rect 20190 7040 20254 7044
rect 6380 6556 6444 6560
rect 6380 6500 6384 6556
rect 6384 6500 6440 6556
rect 6440 6500 6444 6556
rect 6380 6496 6444 6500
rect 6460 6556 6524 6560
rect 6460 6500 6464 6556
rect 6464 6500 6520 6556
rect 6520 6500 6524 6556
rect 6460 6496 6524 6500
rect 6540 6556 6604 6560
rect 6540 6500 6544 6556
rect 6544 6500 6600 6556
rect 6600 6500 6604 6556
rect 6540 6496 6604 6500
rect 6620 6556 6684 6560
rect 6620 6500 6624 6556
rect 6624 6500 6680 6556
rect 6680 6500 6684 6556
rect 6620 6496 6684 6500
rect 11808 6556 11872 6560
rect 11808 6500 11812 6556
rect 11812 6500 11868 6556
rect 11868 6500 11872 6556
rect 11808 6496 11872 6500
rect 11888 6556 11952 6560
rect 11888 6500 11892 6556
rect 11892 6500 11948 6556
rect 11948 6500 11952 6556
rect 11888 6496 11952 6500
rect 11968 6556 12032 6560
rect 11968 6500 11972 6556
rect 11972 6500 12028 6556
rect 12028 6500 12032 6556
rect 11968 6496 12032 6500
rect 12048 6556 12112 6560
rect 12048 6500 12052 6556
rect 12052 6500 12108 6556
rect 12108 6500 12112 6556
rect 12048 6496 12112 6500
rect 17236 6556 17300 6560
rect 17236 6500 17240 6556
rect 17240 6500 17296 6556
rect 17296 6500 17300 6556
rect 17236 6496 17300 6500
rect 17316 6556 17380 6560
rect 17316 6500 17320 6556
rect 17320 6500 17376 6556
rect 17376 6500 17380 6556
rect 17316 6496 17380 6500
rect 17396 6556 17460 6560
rect 17396 6500 17400 6556
rect 17400 6500 17456 6556
rect 17456 6500 17460 6556
rect 17396 6496 17460 6500
rect 17476 6556 17540 6560
rect 17476 6500 17480 6556
rect 17480 6500 17536 6556
rect 17536 6500 17540 6556
rect 17476 6496 17540 6500
rect 22664 6556 22728 6560
rect 22664 6500 22668 6556
rect 22668 6500 22724 6556
rect 22724 6500 22728 6556
rect 22664 6496 22728 6500
rect 22744 6556 22808 6560
rect 22744 6500 22748 6556
rect 22748 6500 22804 6556
rect 22804 6500 22808 6556
rect 22744 6496 22808 6500
rect 22824 6556 22888 6560
rect 22824 6500 22828 6556
rect 22828 6500 22884 6556
rect 22884 6500 22888 6556
rect 22824 6496 22888 6500
rect 22904 6556 22968 6560
rect 22904 6500 22908 6556
rect 22908 6500 22964 6556
rect 22964 6500 22968 6556
rect 22904 6496 22968 6500
rect 3666 6012 3730 6016
rect 3666 5956 3670 6012
rect 3670 5956 3726 6012
rect 3726 5956 3730 6012
rect 3666 5952 3730 5956
rect 3746 6012 3810 6016
rect 3746 5956 3750 6012
rect 3750 5956 3806 6012
rect 3806 5956 3810 6012
rect 3746 5952 3810 5956
rect 3826 6012 3890 6016
rect 3826 5956 3830 6012
rect 3830 5956 3886 6012
rect 3886 5956 3890 6012
rect 3826 5952 3890 5956
rect 3906 6012 3970 6016
rect 3906 5956 3910 6012
rect 3910 5956 3966 6012
rect 3966 5956 3970 6012
rect 3906 5952 3970 5956
rect 9094 6012 9158 6016
rect 9094 5956 9098 6012
rect 9098 5956 9154 6012
rect 9154 5956 9158 6012
rect 9094 5952 9158 5956
rect 9174 6012 9238 6016
rect 9174 5956 9178 6012
rect 9178 5956 9234 6012
rect 9234 5956 9238 6012
rect 9174 5952 9238 5956
rect 9254 6012 9318 6016
rect 9254 5956 9258 6012
rect 9258 5956 9314 6012
rect 9314 5956 9318 6012
rect 9254 5952 9318 5956
rect 9334 6012 9398 6016
rect 9334 5956 9338 6012
rect 9338 5956 9394 6012
rect 9394 5956 9398 6012
rect 9334 5952 9398 5956
rect 14522 6012 14586 6016
rect 14522 5956 14526 6012
rect 14526 5956 14582 6012
rect 14582 5956 14586 6012
rect 14522 5952 14586 5956
rect 14602 6012 14666 6016
rect 14602 5956 14606 6012
rect 14606 5956 14662 6012
rect 14662 5956 14666 6012
rect 14602 5952 14666 5956
rect 14682 6012 14746 6016
rect 14682 5956 14686 6012
rect 14686 5956 14742 6012
rect 14742 5956 14746 6012
rect 14682 5952 14746 5956
rect 14762 6012 14826 6016
rect 14762 5956 14766 6012
rect 14766 5956 14822 6012
rect 14822 5956 14826 6012
rect 14762 5952 14826 5956
rect 19950 6012 20014 6016
rect 19950 5956 19954 6012
rect 19954 5956 20010 6012
rect 20010 5956 20014 6012
rect 19950 5952 20014 5956
rect 20030 6012 20094 6016
rect 20030 5956 20034 6012
rect 20034 5956 20090 6012
rect 20090 5956 20094 6012
rect 20030 5952 20094 5956
rect 20110 6012 20174 6016
rect 20110 5956 20114 6012
rect 20114 5956 20170 6012
rect 20170 5956 20174 6012
rect 20110 5952 20174 5956
rect 20190 6012 20254 6016
rect 20190 5956 20194 6012
rect 20194 5956 20250 6012
rect 20250 5956 20254 6012
rect 20190 5952 20254 5956
rect 6380 5468 6444 5472
rect 6380 5412 6384 5468
rect 6384 5412 6440 5468
rect 6440 5412 6444 5468
rect 6380 5408 6444 5412
rect 6460 5468 6524 5472
rect 6460 5412 6464 5468
rect 6464 5412 6520 5468
rect 6520 5412 6524 5468
rect 6460 5408 6524 5412
rect 6540 5468 6604 5472
rect 6540 5412 6544 5468
rect 6544 5412 6600 5468
rect 6600 5412 6604 5468
rect 6540 5408 6604 5412
rect 6620 5468 6684 5472
rect 6620 5412 6624 5468
rect 6624 5412 6680 5468
rect 6680 5412 6684 5468
rect 6620 5408 6684 5412
rect 11808 5468 11872 5472
rect 11808 5412 11812 5468
rect 11812 5412 11868 5468
rect 11868 5412 11872 5468
rect 11808 5408 11872 5412
rect 11888 5468 11952 5472
rect 11888 5412 11892 5468
rect 11892 5412 11948 5468
rect 11948 5412 11952 5468
rect 11888 5408 11952 5412
rect 11968 5468 12032 5472
rect 11968 5412 11972 5468
rect 11972 5412 12028 5468
rect 12028 5412 12032 5468
rect 11968 5408 12032 5412
rect 12048 5468 12112 5472
rect 12048 5412 12052 5468
rect 12052 5412 12108 5468
rect 12108 5412 12112 5468
rect 12048 5408 12112 5412
rect 17236 5468 17300 5472
rect 17236 5412 17240 5468
rect 17240 5412 17296 5468
rect 17296 5412 17300 5468
rect 17236 5408 17300 5412
rect 17316 5468 17380 5472
rect 17316 5412 17320 5468
rect 17320 5412 17376 5468
rect 17376 5412 17380 5468
rect 17316 5408 17380 5412
rect 17396 5468 17460 5472
rect 17396 5412 17400 5468
rect 17400 5412 17456 5468
rect 17456 5412 17460 5468
rect 17396 5408 17460 5412
rect 17476 5468 17540 5472
rect 17476 5412 17480 5468
rect 17480 5412 17536 5468
rect 17536 5412 17540 5468
rect 17476 5408 17540 5412
rect 22664 5468 22728 5472
rect 22664 5412 22668 5468
rect 22668 5412 22724 5468
rect 22724 5412 22728 5468
rect 22664 5408 22728 5412
rect 22744 5468 22808 5472
rect 22744 5412 22748 5468
rect 22748 5412 22804 5468
rect 22804 5412 22808 5468
rect 22744 5408 22808 5412
rect 22824 5468 22888 5472
rect 22824 5412 22828 5468
rect 22828 5412 22884 5468
rect 22884 5412 22888 5468
rect 22824 5408 22888 5412
rect 22904 5468 22968 5472
rect 22904 5412 22908 5468
rect 22908 5412 22964 5468
rect 22964 5412 22968 5468
rect 22904 5408 22968 5412
rect 3666 4924 3730 4928
rect 3666 4868 3670 4924
rect 3670 4868 3726 4924
rect 3726 4868 3730 4924
rect 3666 4864 3730 4868
rect 3746 4924 3810 4928
rect 3746 4868 3750 4924
rect 3750 4868 3806 4924
rect 3806 4868 3810 4924
rect 3746 4864 3810 4868
rect 3826 4924 3890 4928
rect 3826 4868 3830 4924
rect 3830 4868 3886 4924
rect 3886 4868 3890 4924
rect 3826 4864 3890 4868
rect 3906 4924 3970 4928
rect 3906 4868 3910 4924
rect 3910 4868 3966 4924
rect 3966 4868 3970 4924
rect 3906 4864 3970 4868
rect 9094 4924 9158 4928
rect 9094 4868 9098 4924
rect 9098 4868 9154 4924
rect 9154 4868 9158 4924
rect 9094 4864 9158 4868
rect 9174 4924 9238 4928
rect 9174 4868 9178 4924
rect 9178 4868 9234 4924
rect 9234 4868 9238 4924
rect 9174 4864 9238 4868
rect 9254 4924 9318 4928
rect 9254 4868 9258 4924
rect 9258 4868 9314 4924
rect 9314 4868 9318 4924
rect 9254 4864 9318 4868
rect 9334 4924 9398 4928
rect 9334 4868 9338 4924
rect 9338 4868 9394 4924
rect 9394 4868 9398 4924
rect 9334 4864 9398 4868
rect 14522 4924 14586 4928
rect 14522 4868 14526 4924
rect 14526 4868 14582 4924
rect 14582 4868 14586 4924
rect 14522 4864 14586 4868
rect 14602 4924 14666 4928
rect 14602 4868 14606 4924
rect 14606 4868 14662 4924
rect 14662 4868 14666 4924
rect 14602 4864 14666 4868
rect 14682 4924 14746 4928
rect 14682 4868 14686 4924
rect 14686 4868 14742 4924
rect 14742 4868 14746 4924
rect 14682 4864 14746 4868
rect 14762 4924 14826 4928
rect 14762 4868 14766 4924
rect 14766 4868 14822 4924
rect 14822 4868 14826 4924
rect 14762 4864 14826 4868
rect 19950 4924 20014 4928
rect 19950 4868 19954 4924
rect 19954 4868 20010 4924
rect 20010 4868 20014 4924
rect 19950 4864 20014 4868
rect 20030 4924 20094 4928
rect 20030 4868 20034 4924
rect 20034 4868 20090 4924
rect 20090 4868 20094 4924
rect 20030 4864 20094 4868
rect 20110 4924 20174 4928
rect 20110 4868 20114 4924
rect 20114 4868 20170 4924
rect 20170 4868 20174 4924
rect 20110 4864 20174 4868
rect 20190 4924 20254 4928
rect 20190 4868 20194 4924
rect 20194 4868 20250 4924
rect 20250 4868 20254 4924
rect 20190 4864 20254 4868
rect 6380 4380 6444 4384
rect 6380 4324 6384 4380
rect 6384 4324 6440 4380
rect 6440 4324 6444 4380
rect 6380 4320 6444 4324
rect 6460 4380 6524 4384
rect 6460 4324 6464 4380
rect 6464 4324 6520 4380
rect 6520 4324 6524 4380
rect 6460 4320 6524 4324
rect 6540 4380 6604 4384
rect 6540 4324 6544 4380
rect 6544 4324 6600 4380
rect 6600 4324 6604 4380
rect 6540 4320 6604 4324
rect 6620 4380 6684 4384
rect 6620 4324 6624 4380
rect 6624 4324 6680 4380
rect 6680 4324 6684 4380
rect 6620 4320 6684 4324
rect 11808 4380 11872 4384
rect 11808 4324 11812 4380
rect 11812 4324 11868 4380
rect 11868 4324 11872 4380
rect 11808 4320 11872 4324
rect 11888 4380 11952 4384
rect 11888 4324 11892 4380
rect 11892 4324 11948 4380
rect 11948 4324 11952 4380
rect 11888 4320 11952 4324
rect 11968 4380 12032 4384
rect 11968 4324 11972 4380
rect 11972 4324 12028 4380
rect 12028 4324 12032 4380
rect 11968 4320 12032 4324
rect 12048 4380 12112 4384
rect 12048 4324 12052 4380
rect 12052 4324 12108 4380
rect 12108 4324 12112 4380
rect 12048 4320 12112 4324
rect 17236 4380 17300 4384
rect 17236 4324 17240 4380
rect 17240 4324 17296 4380
rect 17296 4324 17300 4380
rect 17236 4320 17300 4324
rect 17316 4380 17380 4384
rect 17316 4324 17320 4380
rect 17320 4324 17376 4380
rect 17376 4324 17380 4380
rect 17316 4320 17380 4324
rect 17396 4380 17460 4384
rect 17396 4324 17400 4380
rect 17400 4324 17456 4380
rect 17456 4324 17460 4380
rect 17396 4320 17460 4324
rect 17476 4380 17540 4384
rect 17476 4324 17480 4380
rect 17480 4324 17536 4380
rect 17536 4324 17540 4380
rect 17476 4320 17540 4324
rect 22664 4380 22728 4384
rect 22664 4324 22668 4380
rect 22668 4324 22724 4380
rect 22724 4324 22728 4380
rect 22664 4320 22728 4324
rect 22744 4380 22808 4384
rect 22744 4324 22748 4380
rect 22748 4324 22804 4380
rect 22804 4324 22808 4380
rect 22744 4320 22808 4324
rect 22824 4380 22888 4384
rect 22824 4324 22828 4380
rect 22828 4324 22884 4380
rect 22884 4324 22888 4380
rect 22824 4320 22888 4324
rect 22904 4380 22968 4384
rect 22904 4324 22908 4380
rect 22908 4324 22964 4380
rect 22964 4324 22968 4380
rect 22904 4320 22968 4324
rect 3666 3836 3730 3840
rect 3666 3780 3670 3836
rect 3670 3780 3726 3836
rect 3726 3780 3730 3836
rect 3666 3776 3730 3780
rect 3746 3836 3810 3840
rect 3746 3780 3750 3836
rect 3750 3780 3806 3836
rect 3806 3780 3810 3836
rect 3746 3776 3810 3780
rect 3826 3836 3890 3840
rect 3826 3780 3830 3836
rect 3830 3780 3886 3836
rect 3886 3780 3890 3836
rect 3826 3776 3890 3780
rect 3906 3836 3970 3840
rect 3906 3780 3910 3836
rect 3910 3780 3966 3836
rect 3966 3780 3970 3836
rect 3906 3776 3970 3780
rect 9094 3836 9158 3840
rect 9094 3780 9098 3836
rect 9098 3780 9154 3836
rect 9154 3780 9158 3836
rect 9094 3776 9158 3780
rect 9174 3836 9238 3840
rect 9174 3780 9178 3836
rect 9178 3780 9234 3836
rect 9234 3780 9238 3836
rect 9174 3776 9238 3780
rect 9254 3836 9318 3840
rect 9254 3780 9258 3836
rect 9258 3780 9314 3836
rect 9314 3780 9318 3836
rect 9254 3776 9318 3780
rect 9334 3836 9398 3840
rect 9334 3780 9338 3836
rect 9338 3780 9394 3836
rect 9394 3780 9398 3836
rect 9334 3776 9398 3780
rect 14522 3836 14586 3840
rect 14522 3780 14526 3836
rect 14526 3780 14582 3836
rect 14582 3780 14586 3836
rect 14522 3776 14586 3780
rect 14602 3836 14666 3840
rect 14602 3780 14606 3836
rect 14606 3780 14662 3836
rect 14662 3780 14666 3836
rect 14602 3776 14666 3780
rect 14682 3836 14746 3840
rect 14682 3780 14686 3836
rect 14686 3780 14742 3836
rect 14742 3780 14746 3836
rect 14682 3776 14746 3780
rect 14762 3836 14826 3840
rect 14762 3780 14766 3836
rect 14766 3780 14822 3836
rect 14822 3780 14826 3836
rect 14762 3776 14826 3780
rect 19950 3836 20014 3840
rect 19950 3780 19954 3836
rect 19954 3780 20010 3836
rect 20010 3780 20014 3836
rect 19950 3776 20014 3780
rect 20030 3836 20094 3840
rect 20030 3780 20034 3836
rect 20034 3780 20090 3836
rect 20090 3780 20094 3836
rect 20030 3776 20094 3780
rect 20110 3836 20174 3840
rect 20110 3780 20114 3836
rect 20114 3780 20170 3836
rect 20170 3780 20174 3836
rect 20110 3776 20174 3780
rect 20190 3836 20254 3840
rect 20190 3780 20194 3836
rect 20194 3780 20250 3836
rect 20250 3780 20254 3836
rect 20190 3776 20254 3780
rect 6380 3292 6444 3296
rect 6380 3236 6384 3292
rect 6384 3236 6440 3292
rect 6440 3236 6444 3292
rect 6380 3232 6444 3236
rect 6460 3292 6524 3296
rect 6460 3236 6464 3292
rect 6464 3236 6520 3292
rect 6520 3236 6524 3292
rect 6460 3232 6524 3236
rect 6540 3292 6604 3296
rect 6540 3236 6544 3292
rect 6544 3236 6600 3292
rect 6600 3236 6604 3292
rect 6540 3232 6604 3236
rect 6620 3292 6684 3296
rect 6620 3236 6624 3292
rect 6624 3236 6680 3292
rect 6680 3236 6684 3292
rect 6620 3232 6684 3236
rect 11808 3292 11872 3296
rect 11808 3236 11812 3292
rect 11812 3236 11868 3292
rect 11868 3236 11872 3292
rect 11808 3232 11872 3236
rect 11888 3292 11952 3296
rect 11888 3236 11892 3292
rect 11892 3236 11948 3292
rect 11948 3236 11952 3292
rect 11888 3232 11952 3236
rect 11968 3292 12032 3296
rect 11968 3236 11972 3292
rect 11972 3236 12028 3292
rect 12028 3236 12032 3292
rect 11968 3232 12032 3236
rect 12048 3292 12112 3296
rect 12048 3236 12052 3292
rect 12052 3236 12108 3292
rect 12108 3236 12112 3292
rect 12048 3232 12112 3236
rect 17236 3292 17300 3296
rect 17236 3236 17240 3292
rect 17240 3236 17296 3292
rect 17296 3236 17300 3292
rect 17236 3232 17300 3236
rect 17316 3292 17380 3296
rect 17316 3236 17320 3292
rect 17320 3236 17376 3292
rect 17376 3236 17380 3292
rect 17316 3232 17380 3236
rect 17396 3292 17460 3296
rect 17396 3236 17400 3292
rect 17400 3236 17456 3292
rect 17456 3236 17460 3292
rect 17396 3232 17460 3236
rect 17476 3292 17540 3296
rect 17476 3236 17480 3292
rect 17480 3236 17536 3292
rect 17536 3236 17540 3292
rect 17476 3232 17540 3236
rect 22664 3292 22728 3296
rect 22664 3236 22668 3292
rect 22668 3236 22724 3292
rect 22724 3236 22728 3292
rect 22664 3232 22728 3236
rect 22744 3292 22808 3296
rect 22744 3236 22748 3292
rect 22748 3236 22804 3292
rect 22804 3236 22808 3292
rect 22744 3232 22808 3236
rect 22824 3292 22888 3296
rect 22824 3236 22828 3292
rect 22828 3236 22884 3292
rect 22884 3236 22888 3292
rect 22824 3232 22888 3236
rect 22904 3292 22968 3296
rect 22904 3236 22908 3292
rect 22908 3236 22964 3292
rect 22964 3236 22968 3292
rect 22904 3232 22968 3236
rect 3666 2748 3730 2752
rect 3666 2692 3670 2748
rect 3670 2692 3726 2748
rect 3726 2692 3730 2748
rect 3666 2688 3730 2692
rect 3746 2748 3810 2752
rect 3746 2692 3750 2748
rect 3750 2692 3806 2748
rect 3806 2692 3810 2748
rect 3746 2688 3810 2692
rect 3826 2748 3890 2752
rect 3826 2692 3830 2748
rect 3830 2692 3886 2748
rect 3886 2692 3890 2748
rect 3826 2688 3890 2692
rect 3906 2748 3970 2752
rect 3906 2692 3910 2748
rect 3910 2692 3966 2748
rect 3966 2692 3970 2748
rect 3906 2688 3970 2692
rect 9094 2748 9158 2752
rect 9094 2692 9098 2748
rect 9098 2692 9154 2748
rect 9154 2692 9158 2748
rect 9094 2688 9158 2692
rect 9174 2748 9238 2752
rect 9174 2692 9178 2748
rect 9178 2692 9234 2748
rect 9234 2692 9238 2748
rect 9174 2688 9238 2692
rect 9254 2748 9318 2752
rect 9254 2692 9258 2748
rect 9258 2692 9314 2748
rect 9314 2692 9318 2748
rect 9254 2688 9318 2692
rect 9334 2748 9398 2752
rect 9334 2692 9338 2748
rect 9338 2692 9394 2748
rect 9394 2692 9398 2748
rect 9334 2688 9398 2692
rect 14522 2748 14586 2752
rect 14522 2692 14526 2748
rect 14526 2692 14582 2748
rect 14582 2692 14586 2748
rect 14522 2688 14586 2692
rect 14602 2748 14666 2752
rect 14602 2692 14606 2748
rect 14606 2692 14662 2748
rect 14662 2692 14666 2748
rect 14602 2688 14666 2692
rect 14682 2748 14746 2752
rect 14682 2692 14686 2748
rect 14686 2692 14742 2748
rect 14742 2692 14746 2748
rect 14682 2688 14746 2692
rect 14762 2748 14826 2752
rect 14762 2692 14766 2748
rect 14766 2692 14822 2748
rect 14822 2692 14826 2748
rect 14762 2688 14826 2692
rect 19950 2748 20014 2752
rect 19950 2692 19954 2748
rect 19954 2692 20010 2748
rect 20010 2692 20014 2748
rect 19950 2688 20014 2692
rect 20030 2748 20094 2752
rect 20030 2692 20034 2748
rect 20034 2692 20090 2748
rect 20090 2692 20094 2748
rect 20030 2688 20094 2692
rect 20110 2748 20174 2752
rect 20110 2692 20114 2748
rect 20114 2692 20170 2748
rect 20170 2692 20174 2748
rect 20110 2688 20174 2692
rect 20190 2748 20254 2752
rect 20190 2692 20194 2748
rect 20194 2692 20250 2748
rect 20250 2692 20254 2748
rect 20190 2688 20254 2692
rect 6380 2204 6444 2208
rect 6380 2148 6384 2204
rect 6384 2148 6440 2204
rect 6440 2148 6444 2204
rect 6380 2144 6444 2148
rect 6460 2204 6524 2208
rect 6460 2148 6464 2204
rect 6464 2148 6520 2204
rect 6520 2148 6524 2204
rect 6460 2144 6524 2148
rect 6540 2204 6604 2208
rect 6540 2148 6544 2204
rect 6544 2148 6600 2204
rect 6600 2148 6604 2204
rect 6540 2144 6604 2148
rect 6620 2204 6684 2208
rect 6620 2148 6624 2204
rect 6624 2148 6680 2204
rect 6680 2148 6684 2204
rect 6620 2144 6684 2148
rect 11808 2204 11872 2208
rect 11808 2148 11812 2204
rect 11812 2148 11868 2204
rect 11868 2148 11872 2204
rect 11808 2144 11872 2148
rect 11888 2204 11952 2208
rect 11888 2148 11892 2204
rect 11892 2148 11948 2204
rect 11948 2148 11952 2204
rect 11888 2144 11952 2148
rect 11968 2204 12032 2208
rect 11968 2148 11972 2204
rect 11972 2148 12028 2204
rect 12028 2148 12032 2204
rect 11968 2144 12032 2148
rect 12048 2204 12112 2208
rect 12048 2148 12052 2204
rect 12052 2148 12108 2204
rect 12108 2148 12112 2204
rect 12048 2144 12112 2148
rect 17236 2204 17300 2208
rect 17236 2148 17240 2204
rect 17240 2148 17296 2204
rect 17296 2148 17300 2204
rect 17236 2144 17300 2148
rect 17316 2204 17380 2208
rect 17316 2148 17320 2204
rect 17320 2148 17376 2204
rect 17376 2148 17380 2204
rect 17316 2144 17380 2148
rect 17396 2204 17460 2208
rect 17396 2148 17400 2204
rect 17400 2148 17456 2204
rect 17456 2148 17460 2204
rect 17396 2144 17460 2148
rect 17476 2204 17540 2208
rect 17476 2148 17480 2204
rect 17480 2148 17536 2204
rect 17536 2148 17540 2204
rect 17476 2144 17540 2148
rect 22664 2204 22728 2208
rect 22664 2148 22668 2204
rect 22668 2148 22724 2204
rect 22724 2148 22728 2204
rect 22664 2144 22728 2148
rect 22744 2204 22808 2208
rect 22744 2148 22748 2204
rect 22748 2148 22804 2204
rect 22804 2148 22808 2204
rect 22744 2144 22808 2148
rect 22824 2204 22888 2208
rect 22824 2148 22828 2204
rect 22828 2148 22884 2204
rect 22884 2148 22888 2204
rect 22824 2144 22888 2148
rect 22904 2204 22968 2208
rect 22904 2148 22908 2204
rect 22908 2148 22964 2204
rect 22964 2148 22968 2204
rect 22904 2144 22968 2148
<< metal4 >>
rect 3658 21248 3978 21808
rect 3658 21184 3666 21248
rect 3730 21184 3746 21248
rect 3810 21184 3826 21248
rect 3890 21184 3906 21248
rect 3970 21184 3978 21248
rect 3658 20160 3978 21184
rect 3658 20096 3666 20160
rect 3730 20096 3746 20160
rect 3810 20096 3826 20160
rect 3890 20096 3906 20160
rect 3970 20096 3978 20160
rect 3658 19072 3978 20096
rect 3658 19008 3666 19072
rect 3730 19008 3746 19072
rect 3810 19008 3826 19072
rect 3890 19008 3906 19072
rect 3970 19008 3978 19072
rect 3658 17984 3978 19008
rect 3658 17920 3666 17984
rect 3730 17920 3746 17984
rect 3810 17920 3826 17984
rect 3890 17920 3906 17984
rect 3970 17920 3978 17984
rect 3658 16896 3978 17920
rect 3658 16832 3666 16896
rect 3730 16832 3746 16896
rect 3810 16832 3826 16896
rect 3890 16832 3906 16896
rect 3970 16832 3978 16896
rect 3658 15808 3978 16832
rect 3658 15744 3666 15808
rect 3730 15744 3746 15808
rect 3810 15744 3826 15808
rect 3890 15744 3906 15808
rect 3970 15744 3978 15808
rect 3658 14720 3978 15744
rect 3658 14656 3666 14720
rect 3730 14656 3746 14720
rect 3810 14656 3826 14720
rect 3890 14656 3906 14720
rect 3970 14656 3978 14720
rect 3658 13632 3978 14656
rect 3658 13568 3666 13632
rect 3730 13568 3746 13632
rect 3810 13568 3826 13632
rect 3890 13568 3906 13632
rect 3970 13568 3978 13632
rect 3658 12544 3978 13568
rect 3658 12480 3666 12544
rect 3730 12480 3746 12544
rect 3810 12480 3826 12544
rect 3890 12480 3906 12544
rect 3970 12480 3978 12544
rect 3658 11456 3978 12480
rect 3658 11392 3666 11456
rect 3730 11392 3746 11456
rect 3810 11392 3826 11456
rect 3890 11392 3906 11456
rect 3970 11392 3978 11456
rect 3658 10368 3978 11392
rect 3658 10304 3666 10368
rect 3730 10304 3746 10368
rect 3810 10304 3826 10368
rect 3890 10304 3906 10368
rect 3970 10304 3978 10368
rect 3658 9280 3978 10304
rect 3658 9216 3666 9280
rect 3730 9216 3746 9280
rect 3810 9216 3826 9280
rect 3890 9216 3906 9280
rect 3970 9216 3978 9280
rect 3658 8192 3978 9216
rect 3658 8128 3666 8192
rect 3730 8128 3746 8192
rect 3810 8128 3826 8192
rect 3890 8128 3906 8192
rect 3970 8128 3978 8192
rect 3658 7104 3978 8128
rect 3658 7040 3666 7104
rect 3730 7040 3746 7104
rect 3810 7040 3826 7104
rect 3890 7040 3906 7104
rect 3970 7040 3978 7104
rect 3658 6016 3978 7040
rect 3658 5952 3666 6016
rect 3730 5952 3746 6016
rect 3810 5952 3826 6016
rect 3890 5952 3906 6016
rect 3970 5952 3978 6016
rect 3658 4928 3978 5952
rect 3658 4864 3666 4928
rect 3730 4864 3746 4928
rect 3810 4864 3826 4928
rect 3890 4864 3906 4928
rect 3970 4864 3978 4928
rect 3658 3840 3978 4864
rect 3658 3776 3666 3840
rect 3730 3776 3746 3840
rect 3810 3776 3826 3840
rect 3890 3776 3906 3840
rect 3970 3776 3978 3840
rect 3658 2752 3978 3776
rect 3658 2688 3666 2752
rect 3730 2688 3746 2752
rect 3810 2688 3826 2752
rect 3890 2688 3906 2752
rect 3970 2688 3978 2752
rect 3658 2128 3978 2688
rect 6372 21792 6692 21808
rect 6372 21728 6380 21792
rect 6444 21728 6460 21792
rect 6524 21728 6540 21792
rect 6604 21728 6620 21792
rect 6684 21728 6692 21792
rect 6372 20704 6692 21728
rect 6372 20640 6380 20704
rect 6444 20640 6460 20704
rect 6524 20640 6540 20704
rect 6604 20640 6620 20704
rect 6684 20640 6692 20704
rect 6372 19616 6692 20640
rect 6372 19552 6380 19616
rect 6444 19552 6460 19616
rect 6524 19552 6540 19616
rect 6604 19552 6620 19616
rect 6684 19552 6692 19616
rect 6372 18528 6692 19552
rect 6372 18464 6380 18528
rect 6444 18464 6460 18528
rect 6524 18464 6540 18528
rect 6604 18464 6620 18528
rect 6684 18464 6692 18528
rect 6372 17440 6692 18464
rect 6372 17376 6380 17440
rect 6444 17376 6460 17440
rect 6524 17376 6540 17440
rect 6604 17376 6620 17440
rect 6684 17376 6692 17440
rect 6372 16352 6692 17376
rect 6372 16288 6380 16352
rect 6444 16288 6460 16352
rect 6524 16288 6540 16352
rect 6604 16288 6620 16352
rect 6684 16288 6692 16352
rect 6372 15264 6692 16288
rect 6372 15200 6380 15264
rect 6444 15200 6460 15264
rect 6524 15200 6540 15264
rect 6604 15200 6620 15264
rect 6684 15200 6692 15264
rect 6372 14176 6692 15200
rect 6372 14112 6380 14176
rect 6444 14112 6460 14176
rect 6524 14112 6540 14176
rect 6604 14112 6620 14176
rect 6684 14112 6692 14176
rect 6372 13088 6692 14112
rect 6372 13024 6380 13088
rect 6444 13024 6460 13088
rect 6524 13024 6540 13088
rect 6604 13024 6620 13088
rect 6684 13024 6692 13088
rect 6372 12000 6692 13024
rect 6372 11936 6380 12000
rect 6444 11936 6460 12000
rect 6524 11936 6540 12000
rect 6604 11936 6620 12000
rect 6684 11936 6692 12000
rect 6372 10912 6692 11936
rect 6372 10848 6380 10912
rect 6444 10848 6460 10912
rect 6524 10848 6540 10912
rect 6604 10848 6620 10912
rect 6684 10848 6692 10912
rect 6372 9824 6692 10848
rect 6372 9760 6380 9824
rect 6444 9760 6460 9824
rect 6524 9760 6540 9824
rect 6604 9760 6620 9824
rect 6684 9760 6692 9824
rect 6372 8736 6692 9760
rect 6372 8672 6380 8736
rect 6444 8672 6460 8736
rect 6524 8672 6540 8736
rect 6604 8672 6620 8736
rect 6684 8672 6692 8736
rect 6372 7648 6692 8672
rect 6372 7584 6380 7648
rect 6444 7584 6460 7648
rect 6524 7584 6540 7648
rect 6604 7584 6620 7648
rect 6684 7584 6692 7648
rect 6372 6560 6692 7584
rect 6372 6496 6380 6560
rect 6444 6496 6460 6560
rect 6524 6496 6540 6560
rect 6604 6496 6620 6560
rect 6684 6496 6692 6560
rect 6372 5472 6692 6496
rect 6372 5408 6380 5472
rect 6444 5408 6460 5472
rect 6524 5408 6540 5472
rect 6604 5408 6620 5472
rect 6684 5408 6692 5472
rect 6372 4384 6692 5408
rect 6372 4320 6380 4384
rect 6444 4320 6460 4384
rect 6524 4320 6540 4384
rect 6604 4320 6620 4384
rect 6684 4320 6692 4384
rect 6372 3296 6692 4320
rect 6372 3232 6380 3296
rect 6444 3232 6460 3296
rect 6524 3232 6540 3296
rect 6604 3232 6620 3296
rect 6684 3232 6692 3296
rect 6372 2208 6692 3232
rect 6372 2144 6380 2208
rect 6444 2144 6460 2208
rect 6524 2144 6540 2208
rect 6604 2144 6620 2208
rect 6684 2144 6692 2208
rect 6372 2128 6692 2144
rect 9086 21248 9406 21808
rect 9086 21184 9094 21248
rect 9158 21184 9174 21248
rect 9238 21184 9254 21248
rect 9318 21184 9334 21248
rect 9398 21184 9406 21248
rect 9086 20160 9406 21184
rect 9086 20096 9094 20160
rect 9158 20096 9174 20160
rect 9238 20096 9254 20160
rect 9318 20096 9334 20160
rect 9398 20096 9406 20160
rect 9086 19072 9406 20096
rect 9086 19008 9094 19072
rect 9158 19008 9174 19072
rect 9238 19008 9254 19072
rect 9318 19008 9334 19072
rect 9398 19008 9406 19072
rect 9086 17984 9406 19008
rect 9086 17920 9094 17984
rect 9158 17920 9174 17984
rect 9238 17920 9254 17984
rect 9318 17920 9334 17984
rect 9398 17920 9406 17984
rect 9086 16896 9406 17920
rect 9086 16832 9094 16896
rect 9158 16832 9174 16896
rect 9238 16832 9254 16896
rect 9318 16832 9334 16896
rect 9398 16832 9406 16896
rect 9086 15808 9406 16832
rect 9086 15744 9094 15808
rect 9158 15744 9174 15808
rect 9238 15744 9254 15808
rect 9318 15744 9334 15808
rect 9398 15744 9406 15808
rect 9086 14720 9406 15744
rect 9086 14656 9094 14720
rect 9158 14656 9174 14720
rect 9238 14656 9254 14720
rect 9318 14656 9334 14720
rect 9398 14656 9406 14720
rect 9086 13632 9406 14656
rect 9086 13568 9094 13632
rect 9158 13568 9174 13632
rect 9238 13568 9254 13632
rect 9318 13568 9334 13632
rect 9398 13568 9406 13632
rect 9086 12544 9406 13568
rect 9086 12480 9094 12544
rect 9158 12480 9174 12544
rect 9238 12480 9254 12544
rect 9318 12480 9334 12544
rect 9398 12480 9406 12544
rect 9086 11456 9406 12480
rect 9086 11392 9094 11456
rect 9158 11392 9174 11456
rect 9238 11392 9254 11456
rect 9318 11392 9334 11456
rect 9398 11392 9406 11456
rect 9086 10368 9406 11392
rect 9086 10304 9094 10368
rect 9158 10304 9174 10368
rect 9238 10304 9254 10368
rect 9318 10304 9334 10368
rect 9398 10304 9406 10368
rect 9086 9280 9406 10304
rect 9086 9216 9094 9280
rect 9158 9216 9174 9280
rect 9238 9216 9254 9280
rect 9318 9216 9334 9280
rect 9398 9216 9406 9280
rect 9086 8192 9406 9216
rect 9086 8128 9094 8192
rect 9158 8128 9174 8192
rect 9238 8128 9254 8192
rect 9318 8128 9334 8192
rect 9398 8128 9406 8192
rect 9086 7104 9406 8128
rect 9086 7040 9094 7104
rect 9158 7040 9174 7104
rect 9238 7040 9254 7104
rect 9318 7040 9334 7104
rect 9398 7040 9406 7104
rect 9086 6016 9406 7040
rect 9086 5952 9094 6016
rect 9158 5952 9174 6016
rect 9238 5952 9254 6016
rect 9318 5952 9334 6016
rect 9398 5952 9406 6016
rect 9086 4928 9406 5952
rect 9086 4864 9094 4928
rect 9158 4864 9174 4928
rect 9238 4864 9254 4928
rect 9318 4864 9334 4928
rect 9398 4864 9406 4928
rect 9086 3840 9406 4864
rect 9086 3776 9094 3840
rect 9158 3776 9174 3840
rect 9238 3776 9254 3840
rect 9318 3776 9334 3840
rect 9398 3776 9406 3840
rect 9086 2752 9406 3776
rect 9086 2688 9094 2752
rect 9158 2688 9174 2752
rect 9238 2688 9254 2752
rect 9318 2688 9334 2752
rect 9398 2688 9406 2752
rect 9086 2128 9406 2688
rect 11800 21792 12120 21808
rect 11800 21728 11808 21792
rect 11872 21728 11888 21792
rect 11952 21728 11968 21792
rect 12032 21728 12048 21792
rect 12112 21728 12120 21792
rect 11800 20704 12120 21728
rect 11800 20640 11808 20704
rect 11872 20640 11888 20704
rect 11952 20640 11968 20704
rect 12032 20640 12048 20704
rect 12112 20640 12120 20704
rect 11800 19616 12120 20640
rect 11800 19552 11808 19616
rect 11872 19552 11888 19616
rect 11952 19552 11968 19616
rect 12032 19552 12048 19616
rect 12112 19552 12120 19616
rect 11800 18528 12120 19552
rect 11800 18464 11808 18528
rect 11872 18464 11888 18528
rect 11952 18464 11968 18528
rect 12032 18464 12048 18528
rect 12112 18464 12120 18528
rect 11800 17440 12120 18464
rect 11800 17376 11808 17440
rect 11872 17376 11888 17440
rect 11952 17376 11968 17440
rect 12032 17376 12048 17440
rect 12112 17376 12120 17440
rect 11800 16352 12120 17376
rect 11800 16288 11808 16352
rect 11872 16288 11888 16352
rect 11952 16288 11968 16352
rect 12032 16288 12048 16352
rect 12112 16288 12120 16352
rect 11800 15264 12120 16288
rect 11800 15200 11808 15264
rect 11872 15200 11888 15264
rect 11952 15200 11968 15264
rect 12032 15200 12048 15264
rect 12112 15200 12120 15264
rect 11800 14176 12120 15200
rect 11800 14112 11808 14176
rect 11872 14112 11888 14176
rect 11952 14112 11968 14176
rect 12032 14112 12048 14176
rect 12112 14112 12120 14176
rect 11800 13088 12120 14112
rect 11800 13024 11808 13088
rect 11872 13024 11888 13088
rect 11952 13024 11968 13088
rect 12032 13024 12048 13088
rect 12112 13024 12120 13088
rect 11800 12000 12120 13024
rect 11800 11936 11808 12000
rect 11872 11936 11888 12000
rect 11952 11936 11968 12000
rect 12032 11936 12048 12000
rect 12112 11936 12120 12000
rect 11800 10912 12120 11936
rect 11800 10848 11808 10912
rect 11872 10848 11888 10912
rect 11952 10848 11968 10912
rect 12032 10848 12048 10912
rect 12112 10848 12120 10912
rect 11800 9824 12120 10848
rect 11800 9760 11808 9824
rect 11872 9760 11888 9824
rect 11952 9760 11968 9824
rect 12032 9760 12048 9824
rect 12112 9760 12120 9824
rect 11800 8736 12120 9760
rect 11800 8672 11808 8736
rect 11872 8672 11888 8736
rect 11952 8672 11968 8736
rect 12032 8672 12048 8736
rect 12112 8672 12120 8736
rect 11800 7648 12120 8672
rect 11800 7584 11808 7648
rect 11872 7584 11888 7648
rect 11952 7584 11968 7648
rect 12032 7584 12048 7648
rect 12112 7584 12120 7648
rect 11800 6560 12120 7584
rect 11800 6496 11808 6560
rect 11872 6496 11888 6560
rect 11952 6496 11968 6560
rect 12032 6496 12048 6560
rect 12112 6496 12120 6560
rect 11800 5472 12120 6496
rect 11800 5408 11808 5472
rect 11872 5408 11888 5472
rect 11952 5408 11968 5472
rect 12032 5408 12048 5472
rect 12112 5408 12120 5472
rect 11800 4384 12120 5408
rect 11800 4320 11808 4384
rect 11872 4320 11888 4384
rect 11952 4320 11968 4384
rect 12032 4320 12048 4384
rect 12112 4320 12120 4384
rect 11800 3296 12120 4320
rect 11800 3232 11808 3296
rect 11872 3232 11888 3296
rect 11952 3232 11968 3296
rect 12032 3232 12048 3296
rect 12112 3232 12120 3296
rect 11800 2208 12120 3232
rect 11800 2144 11808 2208
rect 11872 2144 11888 2208
rect 11952 2144 11968 2208
rect 12032 2144 12048 2208
rect 12112 2144 12120 2208
rect 11800 2128 12120 2144
rect 14514 21248 14834 21808
rect 14514 21184 14522 21248
rect 14586 21184 14602 21248
rect 14666 21184 14682 21248
rect 14746 21184 14762 21248
rect 14826 21184 14834 21248
rect 14514 20160 14834 21184
rect 14514 20096 14522 20160
rect 14586 20096 14602 20160
rect 14666 20096 14682 20160
rect 14746 20096 14762 20160
rect 14826 20096 14834 20160
rect 14514 19072 14834 20096
rect 14514 19008 14522 19072
rect 14586 19008 14602 19072
rect 14666 19008 14682 19072
rect 14746 19008 14762 19072
rect 14826 19008 14834 19072
rect 14514 17984 14834 19008
rect 14514 17920 14522 17984
rect 14586 17920 14602 17984
rect 14666 17920 14682 17984
rect 14746 17920 14762 17984
rect 14826 17920 14834 17984
rect 14514 16896 14834 17920
rect 14514 16832 14522 16896
rect 14586 16832 14602 16896
rect 14666 16832 14682 16896
rect 14746 16832 14762 16896
rect 14826 16832 14834 16896
rect 14514 15808 14834 16832
rect 14514 15744 14522 15808
rect 14586 15744 14602 15808
rect 14666 15744 14682 15808
rect 14746 15744 14762 15808
rect 14826 15744 14834 15808
rect 14514 14720 14834 15744
rect 14514 14656 14522 14720
rect 14586 14656 14602 14720
rect 14666 14656 14682 14720
rect 14746 14656 14762 14720
rect 14826 14656 14834 14720
rect 14514 13632 14834 14656
rect 14514 13568 14522 13632
rect 14586 13568 14602 13632
rect 14666 13568 14682 13632
rect 14746 13568 14762 13632
rect 14826 13568 14834 13632
rect 14514 12544 14834 13568
rect 14514 12480 14522 12544
rect 14586 12480 14602 12544
rect 14666 12480 14682 12544
rect 14746 12480 14762 12544
rect 14826 12480 14834 12544
rect 14514 11456 14834 12480
rect 14514 11392 14522 11456
rect 14586 11392 14602 11456
rect 14666 11392 14682 11456
rect 14746 11392 14762 11456
rect 14826 11392 14834 11456
rect 14514 10368 14834 11392
rect 17228 21792 17548 21808
rect 17228 21728 17236 21792
rect 17300 21728 17316 21792
rect 17380 21728 17396 21792
rect 17460 21728 17476 21792
rect 17540 21728 17548 21792
rect 17228 20704 17548 21728
rect 17228 20640 17236 20704
rect 17300 20640 17316 20704
rect 17380 20640 17396 20704
rect 17460 20640 17476 20704
rect 17540 20640 17548 20704
rect 17228 19616 17548 20640
rect 17228 19552 17236 19616
rect 17300 19552 17316 19616
rect 17380 19552 17396 19616
rect 17460 19552 17476 19616
rect 17540 19552 17548 19616
rect 17228 18528 17548 19552
rect 17228 18464 17236 18528
rect 17300 18464 17316 18528
rect 17380 18464 17396 18528
rect 17460 18464 17476 18528
rect 17540 18464 17548 18528
rect 17228 17440 17548 18464
rect 17228 17376 17236 17440
rect 17300 17376 17316 17440
rect 17380 17376 17396 17440
rect 17460 17376 17476 17440
rect 17540 17376 17548 17440
rect 17228 16352 17548 17376
rect 17228 16288 17236 16352
rect 17300 16288 17316 16352
rect 17380 16288 17396 16352
rect 17460 16288 17476 16352
rect 17540 16288 17548 16352
rect 17228 15264 17548 16288
rect 17228 15200 17236 15264
rect 17300 15200 17316 15264
rect 17380 15200 17396 15264
rect 17460 15200 17476 15264
rect 17540 15200 17548 15264
rect 17228 14176 17548 15200
rect 17228 14112 17236 14176
rect 17300 14112 17316 14176
rect 17380 14112 17396 14176
rect 17460 14112 17476 14176
rect 17540 14112 17548 14176
rect 17228 13088 17548 14112
rect 17228 13024 17236 13088
rect 17300 13024 17316 13088
rect 17380 13024 17396 13088
rect 17460 13024 17476 13088
rect 17540 13024 17548 13088
rect 17228 12000 17548 13024
rect 17228 11936 17236 12000
rect 17300 11936 17316 12000
rect 17380 11936 17396 12000
rect 17460 11936 17476 12000
rect 17540 11936 17548 12000
rect 15147 11116 15213 11117
rect 15147 11052 15148 11116
rect 15212 11052 15213 11116
rect 15147 11051 15213 11052
rect 14514 10304 14522 10368
rect 14586 10304 14602 10368
rect 14666 10304 14682 10368
rect 14746 10304 14762 10368
rect 14826 10304 14834 10368
rect 14514 9280 14834 10304
rect 14514 9216 14522 9280
rect 14586 9216 14602 9280
rect 14666 9216 14682 9280
rect 14746 9216 14762 9280
rect 14826 9216 14834 9280
rect 14514 8192 14834 9216
rect 14514 8128 14522 8192
rect 14586 8128 14602 8192
rect 14666 8128 14682 8192
rect 14746 8128 14762 8192
rect 14826 8128 14834 8192
rect 14514 7104 14834 8128
rect 15150 7445 15210 11051
rect 17228 10912 17548 11936
rect 17228 10848 17236 10912
rect 17300 10848 17316 10912
rect 17380 10848 17396 10912
rect 17460 10848 17476 10912
rect 17540 10848 17548 10912
rect 17228 9824 17548 10848
rect 17228 9760 17236 9824
rect 17300 9760 17316 9824
rect 17380 9760 17396 9824
rect 17460 9760 17476 9824
rect 17540 9760 17548 9824
rect 17228 8736 17548 9760
rect 17228 8672 17236 8736
rect 17300 8672 17316 8736
rect 17380 8672 17396 8736
rect 17460 8672 17476 8736
rect 17540 8672 17548 8736
rect 17228 7648 17548 8672
rect 17228 7584 17236 7648
rect 17300 7584 17316 7648
rect 17380 7584 17396 7648
rect 17460 7584 17476 7648
rect 17540 7584 17548 7648
rect 15147 7444 15213 7445
rect 15147 7380 15148 7444
rect 15212 7380 15213 7444
rect 15147 7379 15213 7380
rect 14514 7040 14522 7104
rect 14586 7040 14602 7104
rect 14666 7040 14682 7104
rect 14746 7040 14762 7104
rect 14826 7040 14834 7104
rect 14514 6016 14834 7040
rect 14514 5952 14522 6016
rect 14586 5952 14602 6016
rect 14666 5952 14682 6016
rect 14746 5952 14762 6016
rect 14826 5952 14834 6016
rect 14514 4928 14834 5952
rect 14514 4864 14522 4928
rect 14586 4864 14602 4928
rect 14666 4864 14682 4928
rect 14746 4864 14762 4928
rect 14826 4864 14834 4928
rect 14514 3840 14834 4864
rect 14514 3776 14522 3840
rect 14586 3776 14602 3840
rect 14666 3776 14682 3840
rect 14746 3776 14762 3840
rect 14826 3776 14834 3840
rect 14514 2752 14834 3776
rect 14514 2688 14522 2752
rect 14586 2688 14602 2752
rect 14666 2688 14682 2752
rect 14746 2688 14762 2752
rect 14826 2688 14834 2752
rect 14514 2128 14834 2688
rect 17228 6560 17548 7584
rect 17228 6496 17236 6560
rect 17300 6496 17316 6560
rect 17380 6496 17396 6560
rect 17460 6496 17476 6560
rect 17540 6496 17548 6560
rect 17228 5472 17548 6496
rect 17228 5408 17236 5472
rect 17300 5408 17316 5472
rect 17380 5408 17396 5472
rect 17460 5408 17476 5472
rect 17540 5408 17548 5472
rect 17228 4384 17548 5408
rect 17228 4320 17236 4384
rect 17300 4320 17316 4384
rect 17380 4320 17396 4384
rect 17460 4320 17476 4384
rect 17540 4320 17548 4384
rect 17228 3296 17548 4320
rect 17228 3232 17236 3296
rect 17300 3232 17316 3296
rect 17380 3232 17396 3296
rect 17460 3232 17476 3296
rect 17540 3232 17548 3296
rect 17228 2208 17548 3232
rect 17228 2144 17236 2208
rect 17300 2144 17316 2208
rect 17380 2144 17396 2208
rect 17460 2144 17476 2208
rect 17540 2144 17548 2208
rect 17228 2128 17548 2144
rect 19942 21248 20262 21808
rect 19942 21184 19950 21248
rect 20014 21184 20030 21248
rect 20094 21184 20110 21248
rect 20174 21184 20190 21248
rect 20254 21184 20262 21248
rect 19942 20160 20262 21184
rect 19942 20096 19950 20160
rect 20014 20096 20030 20160
rect 20094 20096 20110 20160
rect 20174 20096 20190 20160
rect 20254 20096 20262 20160
rect 19942 19072 20262 20096
rect 19942 19008 19950 19072
rect 20014 19008 20030 19072
rect 20094 19008 20110 19072
rect 20174 19008 20190 19072
rect 20254 19008 20262 19072
rect 19942 17984 20262 19008
rect 19942 17920 19950 17984
rect 20014 17920 20030 17984
rect 20094 17920 20110 17984
rect 20174 17920 20190 17984
rect 20254 17920 20262 17984
rect 19942 16896 20262 17920
rect 19942 16832 19950 16896
rect 20014 16832 20030 16896
rect 20094 16832 20110 16896
rect 20174 16832 20190 16896
rect 20254 16832 20262 16896
rect 19942 15808 20262 16832
rect 19942 15744 19950 15808
rect 20014 15744 20030 15808
rect 20094 15744 20110 15808
rect 20174 15744 20190 15808
rect 20254 15744 20262 15808
rect 19942 14720 20262 15744
rect 19942 14656 19950 14720
rect 20014 14656 20030 14720
rect 20094 14656 20110 14720
rect 20174 14656 20190 14720
rect 20254 14656 20262 14720
rect 19942 13632 20262 14656
rect 19942 13568 19950 13632
rect 20014 13568 20030 13632
rect 20094 13568 20110 13632
rect 20174 13568 20190 13632
rect 20254 13568 20262 13632
rect 19942 12544 20262 13568
rect 19942 12480 19950 12544
rect 20014 12480 20030 12544
rect 20094 12480 20110 12544
rect 20174 12480 20190 12544
rect 20254 12480 20262 12544
rect 19942 11456 20262 12480
rect 19942 11392 19950 11456
rect 20014 11392 20030 11456
rect 20094 11392 20110 11456
rect 20174 11392 20190 11456
rect 20254 11392 20262 11456
rect 19942 10368 20262 11392
rect 19942 10304 19950 10368
rect 20014 10304 20030 10368
rect 20094 10304 20110 10368
rect 20174 10304 20190 10368
rect 20254 10304 20262 10368
rect 19942 9280 20262 10304
rect 19942 9216 19950 9280
rect 20014 9216 20030 9280
rect 20094 9216 20110 9280
rect 20174 9216 20190 9280
rect 20254 9216 20262 9280
rect 19942 8192 20262 9216
rect 19942 8128 19950 8192
rect 20014 8128 20030 8192
rect 20094 8128 20110 8192
rect 20174 8128 20190 8192
rect 20254 8128 20262 8192
rect 19942 7104 20262 8128
rect 19942 7040 19950 7104
rect 20014 7040 20030 7104
rect 20094 7040 20110 7104
rect 20174 7040 20190 7104
rect 20254 7040 20262 7104
rect 19942 6016 20262 7040
rect 19942 5952 19950 6016
rect 20014 5952 20030 6016
rect 20094 5952 20110 6016
rect 20174 5952 20190 6016
rect 20254 5952 20262 6016
rect 19942 4928 20262 5952
rect 19942 4864 19950 4928
rect 20014 4864 20030 4928
rect 20094 4864 20110 4928
rect 20174 4864 20190 4928
rect 20254 4864 20262 4928
rect 19942 3840 20262 4864
rect 19942 3776 19950 3840
rect 20014 3776 20030 3840
rect 20094 3776 20110 3840
rect 20174 3776 20190 3840
rect 20254 3776 20262 3840
rect 19942 2752 20262 3776
rect 19942 2688 19950 2752
rect 20014 2688 20030 2752
rect 20094 2688 20110 2752
rect 20174 2688 20190 2752
rect 20254 2688 20262 2752
rect 19942 2128 20262 2688
rect 22656 21792 22976 21808
rect 22656 21728 22664 21792
rect 22728 21728 22744 21792
rect 22808 21728 22824 21792
rect 22888 21728 22904 21792
rect 22968 21728 22976 21792
rect 22656 20704 22976 21728
rect 22656 20640 22664 20704
rect 22728 20640 22744 20704
rect 22808 20640 22824 20704
rect 22888 20640 22904 20704
rect 22968 20640 22976 20704
rect 22656 19616 22976 20640
rect 22656 19552 22664 19616
rect 22728 19552 22744 19616
rect 22808 19552 22824 19616
rect 22888 19552 22904 19616
rect 22968 19552 22976 19616
rect 22656 18528 22976 19552
rect 22656 18464 22664 18528
rect 22728 18464 22744 18528
rect 22808 18464 22824 18528
rect 22888 18464 22904 18528
rect 22968 18464 22976 18528
rect 22656 17440 22976 18464
rect 22656 17376 22664 17440
rect 22728 17376 22744 17440
rect 22808 17376 22824 17440
rect 22888 17376 22904 17440
rect 22968 17376 22976 17440
rect 22656 16352 22976 17376
rect 22656 16288 22664 16352
rect 22728 16288 22744 16352
rect 22808 16288 22824 16352
rect 22888 16288 22904 16352
rect 22968 16288 22976 16352
rect 22656 15264 22976 16288
rect 22656 15200 22664 15264
rect 22728 15200 22744 15264
rect 22808 15200 22824 15264
rect 22888 15200 22904 15264
rect 22968 15200 22976 15264
rect 22656 14176 22976 15200
rect 22656 14112 22664 14176
rect 22728 14112 22744 14176
rect 22808 14112 22824 14176
rect 22888 14112 22904 14176
rect 22968 14112 22976 14176
rect 22656 13088 22976 14112
rect 22656 13024 22664 13088
rect 22728 13024 22744 13088
rect 22808 13024 22824 13088
rect 22888 13024 22904 13088
rect 22968 13024 22976 13088
rect 22656 12000 22976 13024
rect 22656 11936 22664 12000
rect 22728 11936 22744 12000
rect 22808 11936 22824 12000
rect 22888 11936 22904 12000
rect 22968 11936 22976 12000
rect 22656 10912 22976 11936
rect 22656 10848 22664 10912
rect 22728 10848 22744 10912
rect 22808 10848 22824 10912
rect 22888 10848 22904 10912
rect 22968 10848 22976 10912
rect 22656 9824 22976 10848
rect 22656 9760 22664 9824
rect 22728 9760 22744 9824
rect 22808 9760 22824 9824
rect 22888 9760 22904 9824
rect 22968 9760 22976 9824
rect 22656 8736 22976 9760
rect 22656 8672 22664 8736
rect 22728 8672 22744 8736
rect 22808 8672 22824 8736
rect 22888 8672 22904 8736
rect 22968 8672 22976 8736
rect 22656 7648 22976 8672
rect 22656 7584 22664 7648
rect 22728 7584 22744 7648
rect 22808 7584 22824 7648
rect 22888 7584 22904 7648
rect 22968 7584 22976 7648
rect 22656 6560 22976 7584
rect 22656 6496 22664 6560
rect 22728 6496 22744 6560
rect 22808 6496 22824 6560
rect 22888 6496 22904 6560
rect 22968 6496 22976 6560
rect 22656 5472 22976 6496
rect 22656 5408 22664 5472
rect 22728 5408 22744 5472
rect 22808 5408 22824 5472
rect 22888 5408 22904 5472
rect 22968 5408 22976 5472
rect 22656 4384 22976 5408
rect 22656 4320 22664 4384
rect 22728 4320 22744 4384
rect 22808 4320 22824 4384
rect 22888 4320 22904 4384
rect 22968 4320 22976 4384
rect 22656 3296 22976 4320
rect 22656 3232 22664 3296
rect 22728 3232 22744 3296
rect 22808 3232 22824 3296
rect 22888 3232 22904 3296
rect 22968 3232 22976 3296
rect 22656 2208 22976 3232
rect 22656 2144 22664 2208
rect 22728 2144 22744 2208
rect 22808 2144 22824 2208
rect 22888 2144 22904 2208
rect 22968 2144 22976 2208
rect 22656 2128 22976 2144
use sky130_fd_sc_hd__decap_8  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20
timestamp 1676037725
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1676037725
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65
timestamp 1676037725
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75
timestamp 1676037725
transform 1 0 8004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1676037725
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9384 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_102 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_121
timestamp 1676037725
transform 1 0 12236 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_126
timestamp 1676037725
transform 1 0 12696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1676037725
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_22
timestamp 1676037725
transform 1 0 3128 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_30
timestamp 1676037725
transform 1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_36
timestamp 1676037725
transform 1 0 4416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_80
timestamp 1676037725
transform 1 0 8464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_90
timestamp 1676037725
transform 1 0 9384 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_96
timestamp 1676037725
transform 1 0 9936 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_124
timestamp 1676037725
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_136
timestamp 1676037725
transform 1 0 13616 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_156
timestamp 1676037725
transform 1 0 15456 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_9
timestamp 1676037725
transform 1 0 1932 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_17
timestamp 1676037725
transform 1 0 2668 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_25
timestamp 1676037725
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_37
timestamp 1676037725
transform 1 0 4508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_48
timestamp 1676037725
transform 1 0 5520 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_55
timestamp 1676037725
transform 1 0 6164 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_67
timestamp 1676037725
transform 1 0 7268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_107
timestamp 1676037725
transform 1 0 10948 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_115
timestamp 1676037725
transform 1 0 11684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_127
timestamp 1676037725
transform 1 0 12788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp 1676037725
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1676037725
transform 1 0 14720 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_155
timestamp 1676037725
transform 1 0 15364 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_167
timestamp 1676037725
transform 1 0 16468 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_179
timestamp 1676037725
transform 1 0 17572 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1676037725
transform 1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_22
timestamp 1676037725
transform 1 0 3128 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_50
timestamp 1676037725
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp 1676037725
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_130
timestamp 1676037725
transform 1 0 13064 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_142
timestamp 1676037725
transform 1 0 14168 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_156
timestamp 1676037725
transform 1 0 15456 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1676037725
transform 1 0 1748 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1676037725
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_60
timestamp 1676037725
transform 1 0 6624 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1676037725
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1676037725
transform 1 0 9476 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_108
timestamp 1676037725
transform 1 0 11040 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_120
timestamp 1676037725
transform 1 0 12144 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_124
timestamp 1676037725
transform 1 0 12512 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_132
timestamp 1676037725
transform 1 0 13248 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_161
timestamp 1676037725
transform 1 0 15916 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_169
timestamp 1676037725
transform 1 0 16652 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_36
timestamp 1676037725
transform 1 0 4416 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_48
timestamp 1676037725
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_133
timestamp 1676037725
transform 1 0 13340 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_138
timestamp 1676037725
transform 1 0 13800 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_151
timestamp 1676037725
transform 1 0 14996 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_163
timestamp 1676037725
transform 1 0 16100 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_186
timestamp 1676037725
transform 1 0 18216 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_198
timestamp 1676037725
transform 1 0 19320 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_210
timestamp 1676037725
transform 1 0 20424 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1676037725
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1676037725
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_51
timestamp 1676037725
transform 1 0 5796 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_63
timestamp 1676037725
transform 1 0 6900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_75
timestamp 1676037725
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_89
timestamp 1676037725
transform 1 0 9292 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_125
timestamp 1676037725
transform 1 0 12604 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1676037725
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_152
timestamp 1676037725
transform 1 0 15088 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_158
timestamp 1676037725
transform 1 0 15640 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_164
timestamp 1676037725
transform 1 0 16192 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_176
timestamp 1676037725
transform 1 0 17296 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_188
timestamp 1676037725
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_23
timestamp 1676037725
transform 1 0 3220 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1676037725
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_75
timestamp 1676037725
transform 1 0 8004 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_87
timestamp 1676037725
transform 1 0 9108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1676037725
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_133
timestamp 1676037725
transform 1 0 13340 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_142
timestamp 1676037725
transform 1 0 14168 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_154
timestamp 1676037725
transform 1 0 15272 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp 1676037725
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_190
timestamp 1676037725
transform 1 0 18584 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_204
timestamp 1676037725
transform 1 0 19872 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_216
timestamp 1676037725
transform 1 0 20976 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1676037725
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_51
timestamp 1676037725
transform 1 0 5796 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp 1676037725
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_108
timestamp 1676037725
transform 1 0 11040 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_128
timestamp 1676037725
transform 1 0 12880 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1676037725
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_156
timestamp 1676037725
transform 1 0 15456 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_171
timestamp 1676037725
transform 1 0 16836 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_184
timestamp 1676037725
transform 1 0 18032 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1676037725
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_206
timestamp 1676037725
transform 1 0 20056 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_218
timestamp 1676037725
transform 1 0 21160 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_230
timestamp 1676037725
transform 1 0 22264 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_36
timestamp 1676037725
transform 1 0 4416 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_48
timestamp 1676037725
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_121
timestamp 1676037725
transform 1 0 12236 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_131
timestamp 1676037725
transform 1 0 13156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_143
timestamp 1676037725
transform 1 0 14260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_151
timestamp 1676037725
transform 1 0 14996 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_155
timestamp 1676037725
transform 1 0 15364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_175
timestamp 1676037725
transform 1 0 17204 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_183
timestamp 1676037725
transform 1 0 17940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_195
timestamp 1676037725
transform 1 0 19044 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_201
timestamp 1676037725
transform 1 0 19596 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_212
timestamp 1676037725
transform 1 0 20608 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_11
timestamp 1676037725
transform 1 0 2116 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_16
timestamp 1676037725
transform 1 0 2576 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_49
timestamp 1676037725
transform 1 0 5612 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_70
timestamp 1676037725
transform 1 0 7544 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1676037725
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1676037725
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_108
timestamp 1676037725
transform 1 0 11040 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_120
timestamp 1676037725
transform 1 0 12144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_124
timestamp 1676037725
transform 1 0 12512 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_134
timestamp 1676037725
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_155
timestamp 1676037725
transform 1 0 15364 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_167
timestamp 1676037725
transform 1 0 16468 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_180
timestamp 1676037725
transform 1 0 17664 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1676037725
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_207
timestamp 1676037725
transform 1 0 20148 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_214
timestamp 1676037725
transform 1 0 20792 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_226
timestamp 1676037725
transform 1 0 21896 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_232
timestamp 1676037725
transform 1 0 22448 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_76
timestamp 1676037725
transform 1 0 8096 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_88
timestamp 1676037725
transform 1 0 9200 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1676037725
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_129
timestamp 1676037725
transform 1 0 12972 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_141
timestamp 1676037725
transform 1 0 14076 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_154
timestamp 1676037725
transform 1 0 15272 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_163
timestamp 1676037725
transform 1 0 16100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_174
timestamp 1676037725
transform 1 0 17112 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_184
timestamp 1676037725
transform 1 0 18032 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_192
timestamp 1676037725
transform 1 0 18768 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_201
timestamp 1676037725
transform 1 0 19596 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_209
timestamp 1676037725
transform 1 0 20332 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_215
timestamp 1676037725
transform 1 0 20884 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_9
timestamp 1676037725
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1676037725
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_107
timestamp 1676037725
transform 1 0 10948 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_119
timestamp 1676037725
transform 1 0 12052 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_127
timestamp 1676037725
transform 1 0 12788 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_132
timestamp 1676037725
transform 1 0 13248 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_145
timestamp 1676037725
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_152
timestamp 1676037725
transform 1 0 15088 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_160
timestamp 1676037725
transform 1 0 15824 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_170
timestamp 1676037725
transform 1 0 16744 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_174
timestamp 1676037725
transform 1 0 17112 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_180
timestamp 1676037725
transform 1 0 17664 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_191
timestamp 1676037725
transform 1 0 18676 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1676037725
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_220
timestamp 1676037725
transform 1 0 21344 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_232
timestamp 1676037725
transform 1 0 22448 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_23
timestamp 1676037725
transform 1 0 3220 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_31
timestamp 1676037725
transform 1 0 3956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_50
timestamp 1676037725
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_89
timestamp 1676037725
transform 1 0 9292 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1676037725
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_157
timestamp 1676037725
transform 1 0 15548 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_162
timestamp 1676037725
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_175
timestamp 1676037725
transform 1 0 17204 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_185
timestamp 1676037725
transform 1 0 18124 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_205
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_213
timestamp 1676037725
transform 1 0 20700 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_230
timestamp 1676037725
transform 1 0 22264 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_22
timestamp 1676037725
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_50
timestamp 1676037725
transform 1 0 5704 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_62
timestamp 1676037725
transform 1 0 6808 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1676037725
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_108
timestamp 1676037725
transform 1 0 11040 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_120
timestamp 1676037725
transform 1 0 12144 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1676037725
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_157
timestamp 1676037725
transform 1 0 15548 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_167
timestamp 1676037725
transform 1 0 16468 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_174
timestamp 1676037725
transform 1 0 17112 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_186
timestamp 1676037725
transform 1 0 18216 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_206
timestamp 1676037725
transform 1 0 20056 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_215
timestamp 1676037725
transform 1 0 20884 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_227
timestamp 1676037725
transform 1 0 21988 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_22
timestamp 1676037725
transform 1 0 3128 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_34
timestamp 1676037725
transform 1 0 4232 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1676037725
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_65
timestamp 1676037725
transform 1 0 7084 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_82
timestamp 1676037725
transform 1 0 8648 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_90
timestamp 1676037725
transform 1 0 9384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_107
timestamp 1676037725
transform 1 0 10948 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_117
timestamp 1676037725
transform 1 0 11868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_122
timestamp 1676037725
transform 1 0 12328 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_134
timestamp 1676037725
transform 1 0 13432 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_142
timestamp 1676037725
transform 1 0 14168 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_148
timestamp 1676037725
transform 1 0 14720 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_158
timestamp 1676037725
transform 1 0 15640 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_179
timestamp 1676037725
transform 1 0 17572 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_185
timestamp 1676037725
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_193
timestamp 1676037725
transform 1 0 18860 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_204
timestamp 1676037725
transform 1 0 19872 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_230
timestamp 1676037725
transform 1 0 22264 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_9
timestamp 1676037725
transform 1 0 1932 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_21
timestamp 1676037725
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_59
timestamp 1676037725
transform 1 0 6532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_79
timestamp 1676037725
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_129
timestamp 1676037725
transform 1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1676037725
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_150
timestamp 1676037725
transform 1 0 14904 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_161
timestamp 1676037725
transform 1 0 15916 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_171
timestamp 1676037725
transform 1 0 16836 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_179
timestamp 1676037725
transform 1 0 17572 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_187
timestamp 1676037725
transform 1 0 18308 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_206
timestamp 1676037725
transform 1 0 20056 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_223
timestamp 1676037725
transform 1 0 21620 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_231
timestamp 1676037725
transform 1 0 22356 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_41
timestamp 1676037725
transform 1 0 4876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1676037725
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_149
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_158
timestamp 1676037725
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_173
timestamp 1676037725
transform 1 0 17020 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_182
timestamp 1676037725
transform 1 0 17848 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_194
timestamp 1676037725
transform 1 0 18952 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_198
timestamp 1676037725
transform 1 0 19320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_207
timestamp 1676037725
transform 1 0 20148 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_215
timestamp 1676037725
transform 1 0 20884 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 1676037725
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1676037725
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_40
timestamp 1676037725
transform 1 0 4784 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_46
timestamp 1676037725
transform 1 0 5336 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_71
timestamp 1676037725
transform 1 0 7636 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_108
timestamp 1676037725
transform 1 0 11040 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_129
timestamp 1676037725
transform 1 0 12972 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp 1676037725
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_149
timestamp 1676037725
transform 1 0 14812 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_160
timestamp 1676037725
transform 1 0 15824 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_169
timestamp 1676037725
transform 1 0 16652 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_176
timestamp 1676037725
transform 1 0 17296 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_183
timestamp 1676037725
transform 1 0 17940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1676037725
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_205
timestamp 1676037725
transform 1 0 19964 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_213
timestamp 1676037725
transform 1 0 20700 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_221
timestamp 1676037725
transform 1 0 21436 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_225
timestamp 1676037725
transform 1 0 21804 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_11
timestamp 1676037725
transform 1 0 2116 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_18
timestamp 1676037725
transform 1 0 2760 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_22
timestamp 1676037725
transform 1 0 3128 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_28
timestamp 1676037725
transform 1 0 3680 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_36
timestamp 1676037725
transform 1 0 4416 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_41
timestamp 1676037725
transform 1 0 4876 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_47
timestamp 1676037725
transform 1 0 5428 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1676037725
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_63
timestamp 1676037725
transform 1 0 6900 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_73
timestamp 1676037725
transform 1 0 7820 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_83
timestamp 1676037725
transform 1 0 8740 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_92
timestamp 1676037725
transform 1 0 9568 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1676037725
transform 1 0 11960 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_131
timestamp 1676037725
transform 1 0 13156 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_140
timestamp 1676037725
transform 1 0 13984 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp 1676037725
transform 1 0 15732 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1676037725
transform 1 0 17480 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_190
timestamp 1676037725
transform 1 0 18584 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_202
timestamp 1676037725
transform 1 0 19688 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_214
timestamp 1676037725
transform 1 0 20792 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_230
timestamp 1676037725
transform 1 0 22264 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_11
timestamp 1676037725
transform 1 0 2116 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_18
timestamp 1676037725
transform 1 0 2760 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1676037725
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_90
timestamp 1676037725
transform 1 0 9384 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_110
timestamp 1676037725
transform 1 0 11224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_128
timestamp 1676037725
transform 1 0 12880 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1676037725
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_150
timestamp 1676037725
transform 1 0 14904 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1676037725
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_172
timestamp 1676037725
transform 1 0 16928 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_176
timestamp 1676037725
transform 1 0 17296 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_186
timestamp 1676037725
transform 1 0 18216 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_206
timestamp 1676037725
transform 1 0 20056 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_218
timestamp 1676037725
transform 1 0 21160 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_230
timestamp 1676037725
transform 1 0 22264 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_9
timestamp 1676037725
transform 1 0 1932 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_14
timestamp 1676037725
transform 1 0 2392 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_22
timestamp 1676037725
transform 1 0 3128 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_29
timestamp 1676037725
transform 1 0 3772 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_37
timestamp 1676037725
transform 1 0 4508 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_46
timestamp 1676037725
transform 1 0 5336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1676037725
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_67
timestamp 1676037725
transform 1 0 7268 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_75
timestamp 1676037725
transform 1 0 8004 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_84
timestamp 1676037725
transform 1 0 8832 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_94
timestamp 1676037725
transform 1 0 9752 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1676037725
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_129
timestamp 1676037725
transform 1 0 12972 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_149
timestamp 1676037725
transform 1 0 14812 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_159
timestamp 1676037725
transform 1 0 15732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1676037725
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1676037725
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1676037725
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1676037725
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1676037725
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1676037725
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_12
timestamp 1676037725
transform 1 0 2208 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_25
timestamp 1676037725
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_37
timestamp 1676037725
transform 1 0 4508 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_49
timestamp 1676037725
transform 1 0 5612 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_66
timestamp 1676037725
transform 1 0 7176 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_78
timestamp 1676037725
transform 1 0 8280 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_93
timestamp 1676037725
transform 1 0 9660 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_101
timestamp 1676037725
transform 1 0 10396 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_113
timestamp 1676037725
transform 1 0 11500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_125
timestamp 1676037725
transform 1 0 12604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 1676037725
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1676037725
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1676037725
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1676037725
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1676037725
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_12
timestamp 1676037725
transform 1 0 2208 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_23
timestamp 1676037725
transform 1 0 3220 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_35
timestamp 1676037725
transform 1 0 4324 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_44
timestamp 1676037725
transform 1 0 5152 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_68
timestamp 1676037725
transform 1 0 7360 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_78
timestamp 1676037725
transform 1 0 8280 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_90
timestamp 1676037725
transform 1 0 9384 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_102
timestamp 1676037725
transform 1 0 10488 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1676037725
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1676037725
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1676037725
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1676037725
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1676037725
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1676037725
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1676037725
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_44
timestamp 1676037725
transform 1 0 5152 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_56
timestamp 1676037725
transform 1 0 6256 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_67
timestamp 1676037725
transform 1 0 7268 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_79
timestamp 1676037725
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_90
timestamp 1676037725
transform 1 0 9384 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_103
timestamp 1676037725
transform 1 0 10580 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_112
timestamp 1676037725
transform 1 0 11408 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_124
timestamp 1676037725
transform 1 0 12512 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1676037725
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1676037725
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1676037725
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1676037725
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1676037725
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_20
timestamp 1676037725
transform 1 0 2944 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_32
timestamp 1676037725
transform 1 0 4048 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1676037725
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1676037725
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_75
timestamp 1676037725
transform 1 0 8004 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_83
timestamp 1676037725
transform 1 0 8740 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_118
timestamp 1676037725
transform 1 0 11960 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_130
timestamp 1676037725
transform 1 0 13064 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_142
timestamp 1676037725
transform 1 0 14168 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_154
timestamp 1676037725
transform 1 0 15272 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1676037725
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1676037725
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1676037725
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1676037725
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_25
timestamp 1676037725
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_58
timestamp 1676037725
transform 1 0 6440 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_70
timestamp 1676037725
transform 1 0 7544 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp 1676037725
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_91
timestamp 1676037725
transform 1 0 9476 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_107
timestamp 1676037725
transform 1 0 10948 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_119
timestamp 1676037725
transform 1 0 12052 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_131
timestamp 1676037725
transform 1 0 13156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1676037725
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1676037725
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1676037725
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1676037725
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1676037725
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1676037725
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_26
timestamp 1676037725
transform 1 0 3496 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_38
timestamp 1676037725
transform 1 0 4600 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_49
timestamp 1676037725
transform 1 0 5612 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_70
timestamp 1676037725
transform 1 0 7544 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_79
timestamp 1676037725
transform 1 0 8372 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_87
timestamp 1676037725
transform 1 0 9108 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_97
timestamp 1676037725
transform 1 0 10028 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_106
timestamp 1676037725
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1676037725
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1676037725
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1676037725
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1676037725
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1676037725
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1676037725
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_37
timestamp 1676037725
transform 1 0 4508 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_48
timestamp 1676037725
transform 1 0 5520 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_60
timestamp 1676037725
transform 1 0 6624 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_68
timestamp 1676037725
transform 1 0 7360 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_74
timestamp 1676037725
transform 1 0 7912 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_79
timestamp 1676037725
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_92
timestamp 1676037725
transform 1 0 9568 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_100
timestamp 1676037725
transform 1 0 10304 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_105
timestamp 1676037725
transform 1 0 10764 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_117
timestamp 1676037725
transform 1 0 11868 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_129
timestamp 1676037725
transform 1 0 12972 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1676037725
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1676037725
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1676037725
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1676037725
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1676037725
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1676037725
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1676037725
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1676037725
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_87
timestamp 1676037725
transform 1 0 9108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_99
timestamp 1676037725
transform 1 0 10212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1676037725
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1676037725
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1676037725
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1676037725
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1676037725
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1676037725
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1676037725
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1676037725
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1676037725
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1676037725
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1676037725
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1676037725
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1676037725
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1676037725
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1676037725
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1676037725
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1676037725
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1676037725
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_11
timestamp 1676037725
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1676037725
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1676037725
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1676037725
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1676037725
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1676037725
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1676037725
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1676037725
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1676037725
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1676037725
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1676037725
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1676037725
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1676037725
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1676037725
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1676037725
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1676037725
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1676037725
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1676037725
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1676037725
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1676037725
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1676037725
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1676037725
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1676037725
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1676037725
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1676037725
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1676037725
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1676037725
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1676037725
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1676037725
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1676037725
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1676037725
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1676037725
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1676037725
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1676037725
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_29
timestamp 1676037725
transform 1 0 3772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_41
timestamp 1676037725
transform 1 0 4876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1676037725
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_85
timestamp 1676037725
transform 1 0 8924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_97
timestamp 1676037725
transform 1 0 10028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_109
timestamp 1676037725
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_137
timestamp 1676037725
transform 1 0 13708 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_141
timestamp 1676037725
transform 1 0 14076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_153
timestamp 1676037725
transform 1 0 15180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1676037725
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_193
timestamp 1676037725
transform 1 0 18860 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_197
timestamp 1676037725
transform 1 0 19228 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_209
timestamp 1676037725
transform 1 0 20332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp 1676037725
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 22816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 22816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 22816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 22816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 22816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 22816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 22816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 22816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 22816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 22816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 22816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 22816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 22816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 22816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 22816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 22816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 22816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 22816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 22816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 22816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 22816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 22816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 22816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 22816 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 22816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 22816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 22816 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 22816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 22816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 22816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 22816 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 22816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 22816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 22816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 3680 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 8832 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 13984 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 19136 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _200_
timestamp 1676037725
transform -1 0 22264 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _201_
timestamp 1676037725
transform 1 0 12696 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _204_
timestamp 1676037725
transform 1 0 12328 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _205_
timestamp 1676037725
transform -1 0 10948 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _206_
timestamp 1676037725
transform -1 0 9384 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3220 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and4_4  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7268 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8188 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _211_
timestamp 1676037725
transform -1 0 9568 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11040 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_2  _213_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10304 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_4  _214_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12880 0 1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_2  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14168 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _216_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11224 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13064 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1676037725
transform 1 0 15180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13800 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14812 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_4  _221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4784 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1676037725
transform 1 0 15088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _223_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14444 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_4  _225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14444 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__xnor2_2  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15456 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_4  _227_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17940 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1676037725
transform 1 0 19688 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _229_
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17480 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15456 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_4  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__and2_2  _234_
timestamp 1676037725
transform 1 0 14536 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _235_
timestamp 1676037725
transform 1 0 21988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _236_
timestamp 1676037725
transform 1 0 15732 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _237_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13248 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _238_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15088 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _239_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1676037725
transform -1 0 17296 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _241_
timestamp 1676037725
transform -1 0 15364 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _242_
timestamp 1676037725
transform -1 0 16100 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15640 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _244_
timestamp 1676037725
transform -1 0 16836 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _245_
timestamp 1676037725
transform -1 0 15732 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _246_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16468 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16100 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1676037725
transform -1 0 17112 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _249_
timestamp 1676037725
transform 1 0 15732 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _250_
timestamp 1676037725
transform -1 0 20884 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _251_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13248 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _252_
timestamp 1676037725
transform 1 0 13064 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _253_
timestamp 1676037725
transform 1 0 13064 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  _254_
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _255_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16928 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1676037725
transform 1 0 15088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _257_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _258_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20792 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20608 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _260_
timestamp 1676037725
transform 1 0 18400 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _261_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17204 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _262_
timestamp 1676037725
transform -1 0 18676 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _263_
timestamp 1676037725
transform -1 0 17112 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16192 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17020 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _266_
timestamp 1676037725
transform -1 0 17204 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18124 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _268_
timestamp 1676037725
transform 1 0 20332 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _269_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19320 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _270_
timestamp 1676037725
transform 1 0 19412 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15824 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12604 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15640 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _274_
timestamp 1676037725
transform -1 0 17664 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _275_
timestamp 1676037725
transform -1 0 16652 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _276_
timestamp 1676037725
transform 1 0 21528 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14996 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15272 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12512 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _280_
timestamp 1676037725
transform -1 0 17940 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _281_
timestamp 1676037725
transform 1 0 20516 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20056 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _283_
timestamp 1676037725
transform 1 0 18492 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _284_
timestamp 1676037725
transform 1 0 18584 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18216 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17848 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _287_
timestamp 1676037725
transform 1 0 19780 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _288_
timestamp 1676037725
transform -1 0 20884 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _289_
timestamp 1676037725
transform 1 0 19228 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _290_
timestamp 1676037725
transform 1 0 18676 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _291_
timestamp 1676037725
transform 1 0 17112 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _292_
timestamp 1676037725
transform 1 0 17664 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _293_
timestamp 1676037725
transform -1 0 21528 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _294_
timestamp 1676037725
transform 1 0 19320 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _295_
timestamp 1676037725
transform 1 0 20056 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _296_
timestamp 1676037725
transform -1 0 19596 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _297_
timestamp 1676037725
transform -1 0 18860 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _300_
timestamp 1676037725
transform 1 0 21160 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _301_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20792 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _302_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20056 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14628 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _304_
timestamp 1676037725
transform 1 0 13156 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _305_
timestamp 1676037725
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _306_
timestamp 1676037725
transform 1 0 15640 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _307_
timestamp 1676037725
transform -1 0 14168 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _308_
timestamp 1676037725
transform 1 0 14260 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _309_
timestamp 1676037725
transform 1 0 12696 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _310_
timestamp 1676037725
transform 1 0 13340 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _311_
timestamp 1676037725
transform -1 0 13248 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _312_
timestamp 1676037725
transform -1 0 17572 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _313_
timestamp 1676037725
transform 1 0 12880 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _314_
timestamp 1676037725
transform -1 0 2208 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _315_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12696 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _316_
timestamp 1676037725
transform -1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _317_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8832 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _318_
timestamp 1676037725
transform 1 0 7176 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _319_
timestamp 1676037725
transform 1 0 12420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _320_
timestamp 1676037725
transform 1 0 13064 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _321_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12880 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _322_
timestamp 1676037725
transform 1 0 11684 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _323_
timestamp 1676037725
transform -1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _324_
timestamp 1676037725
transform 1 0 12604 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _325_
timestamp 1676037725
transform 1 0 12236 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _326_
timestamp 1676037725
transform -1 0 11684 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _327_
timestamp 1676037725
transform 1 0 10028 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _328_
timestamp 1676037725
transform 1 0 7636 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _329_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _330_
timestamp 1676037725
transform 1 0 13248 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _331_
timestamp 1676037725
transform 1 0 2944 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_2  _332_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_4  _333_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__o21ai_1  _334_
timestamp 1676037725
transform 1 0 2024 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _335_
timestamp 1676037725
transform 1 0 1840 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _336_
timestamp 1676037725
transform 1 0 11684 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _337_
timestamp 1676037725
transform 1 0 10396 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _338_
timestamp 1676037725
transform -1 0 10580 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _339_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11408 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _340_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10948 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1676037725
transform 1 0 2668 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _342_
timestamp 1676037725
transform 1 0 2116 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _343_
timestamp 1676037725
transform -1 0 9568 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _344_
timestamp 1676037725
transform -1 0 10856 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _345_
timestamp 1676037725
transform -1 0 9476 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _346_
timestamp 1676037725
transform -1 0 8372 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _347_
timestamp 1676037725
transform 1 0 6808 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _348_
timestamp 1676037725
transform 1 0 2576 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _349_
timestamp 1676037725
transform -1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _350_
timestamp 1676037725
transform 1 0 9292 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _351_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10488 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1676037725
transform 1 0 6532 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1676037725
transform -1 0 7176 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _354_
timestamp 1676037725
transform -1 0 8372 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _355_
timestamp 1676037725
transform -1 0 9108 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _356_
timestamp 1676037725
transform -1 0 7544 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _357_
timestamp 1676037725
transform 1 0 4784 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1676037725
transform 1 0 4416 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _359_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 9384 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _360_
timestamp 1676037725
transform 1 0 9384 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _361_
timestamp 1676037725
transform -1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _362_
timestamp 1676037725
transform 1 0 4692 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _363_
timestamp 1676037725
transform 1 0 4324 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _364_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10764 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _365_
timestamp 1676037725
transform 1 0 8096 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _366_
timestamp 1676037725
transform -1 0 7268 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _367_
timestamp 1676037725
transform 1 0 3956 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _368_
timestamp 1676037725
transform 1 0 4508 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _369_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 7360 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _370_
timestamp 1676037725
transform 1 0 2944 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _371_
timestamp 1676037725
transform -1 0 3772 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _372_
timestamp 1676037725
transform -1 0 7268 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _373_
timestamp 1676037725
transform -1 0 5336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1676037725
transform 1 0 11408 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _375_
timestamp 1676037725
transform 1 0 2300 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _376_
timestamp 1676037725
transform 1 0 2116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _377_
timestamp 1676037725
transform 1 0 1932 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _378_
timestamp 1676037725
transform -1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _379_
timestamp 1676037725
transform 1 0 3128 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _380_
timestamp 1676037725
transform 1 0 4600 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _381_
timestamp 1676037725
transform -1 0 4876 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _382_
timestamp 1676037725
transform 1 0 5520 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _383_
timestamp 1676037725
transform 1 0 5428 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _384_
timestamp 1676037725
transform -1 0 7084 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _385_
timestamp 1676037725
transform -1 0 6900 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _386_
timestamp 1676037725
transform 1 0 9108 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _387_
timestamp 1676037725
transform 1 0 8188 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _388_
timestamp 1676037725
transform 1 0 9200 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _389_
timestamp 1676037725
transform 1 0 8096 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _390_
timestamp 1676037725
transform -1 0 11224 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _391_
timestamp 1676037725
transform -1 0 14996 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _392_
timestamp 1676037725
transform -1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _393_
timestamp 1676037725
transform 1 0 2300 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _394_
timestamp 1676037725
transform -1 0 4416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _395_
timestamp 1676037725
transform 1 0 4324 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _396_
timestamp 1676037725
transform 1 0 4784 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _397_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2024 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _398_
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _399_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10948 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _400_
timestamp 1676037725
transform 1 0 6532 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _401_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9476 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _402_
timestamp 1676037725
transform 1 0 9476 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _403_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9476 0 -1 8704
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _404_
timestamp 1676037725
transform 1 0 6900 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _405_
timestamp 1676037725
transform 1 0 5152 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _406_
timestamp 1676037725
transform 1 0 7084 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _407_
timestamp 1676037725
transform 1 0 9568 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _408_
timestamp 1676037725
transform 1 0 6992 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _409_
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _410_
timestamp 1676037725
transform 1 0 9292 0 -1 6528
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _411_
timestamp 1676037725
transform 1 0 9384 0 1 5440
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _412_
timestamp 1676037725
transform 1 0 11408 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _413_
timestamp 1676037725
transform 1 0 9476 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _414_
timestamp 1676037725
transform 1 0 9568 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _415_
timestamp 1676037725
transform -1 0 5796 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _416_
timestamp 1676037725
transform 1 0 1656 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _417_
timestamp 1676037725
transform 1 0 1748 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _418_
timestamp 1676037725
transform 1 0 2024 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _419_
timestamp 1676037725
transform 1 0 6624 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _420_
timestamp 1676037725
transform 1 0 4232 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _421_
timestamp 1676037725
transform 1 0 4140 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _422_
timestamp 1676037725
transform -1 0 5980 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _423_
timestamp 1676037725
transform -1 0 5796 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _424_
timestamp 1676037725
transform 1 0 9568 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _425_
timestamp 1676037725
transform 1 0 1656 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _426_
timestamp 1676037725
transform 1 0 1656 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _427_
timestamp 1676037725
transform 1 0 1748 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _428_
timestamp 1676037725
transform -1 0 5796 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _429_
timestamp 1676037725
transform 1 0 5060 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _430_
timestamp 1676037725
transform 1 0 6900 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _431_
timestamp 1676037725
transform 1 0 7176 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _432_
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _433_
timestamp 1676037725
transform 1 0 9476 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _434_
timestamp 1676037725
transform 1 0 1656 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _435_
timestamp 1676037725
transform -1 0 3220 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _436_
timestamp 1676037725
transform 1 0 4232 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _437_
timestamp 1676037725
transform 1 0 1840 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _438_
timestamp 1676037725
transform 1 0 3956 0 -1 6528
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5704 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1676037725
transform -1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1676037725
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1676037725
transform 1 0 7820 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1676037725
transform 1 0 7820 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15640 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout4
timestamp 1676037725
transform -1 0 16836 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16376 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8280 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout7
timestamp 1676037725
transform -1 0 2760 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11500 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout9
timestamp 1676037725
transform 1 0 2208 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1676037725
transform 1 0 1564 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output2
timestamp 1676037725
transform -1 0 2116 0 1 19584
box -38 -48 590 592
<< labels >>
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 OP
port 0 nsew signal tristate
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 clk
port 1 nsew signal input
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 rst
port 2 nsew signal input
flabel metal4 s 3658 2128 3978 21808 0 FreeSans 1920 90 0 0 vccd1
port 3 nsew power bidirectional
flabel metal4 s 9086 2128 9406 21808 0 FreeSans 1920 90 0 0 vccd1
port 3 nsew power bidirectional
flabel metal4 s 14514 2128 14834 21808 0 FreeSans 1920 90 0 0 vccd1
port 3 nsew power bidirectional
flabel metal4 s 19942 2128 20262 21808 0 FreeSans 1920 90 0 0 vccd1
port 3 nsew power bidirectional
flabel metal4 s 6372 2128 6692 21808 0 FreeSans 1920 90 0 0 vssd1
port 4 nsew ground bidirectional
flabel metal4 s 11800 2128 12120 21808 0 FreeSans 1920 90 0 0 vssd1
port 4 nsew ground bidirectional
flabel metal4 s 17228 2128 17548 21808 0 FreeSans 1920 90 0 0 vssd1
port 4 nsew ground bidirectional
flabel metal4 s 22656 2128 22976 21808 0 FreeSans 1920 90 0 0 vssd1
port 4 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 24000 24000
<< end >>
