// This is the unpowered netlist.
module wrapped_vgatest (clk,
    io_in,
    rst,
    io_out);
 input clk;
 input io_in;
 input rst;
 output [9:0] io_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \vgatest.bitmap.res[0] ;
 wire \vgatest.bitmap.res[1] ;
 wire \vgatest.bitmap.res[2] ;
 wire \vgatest.bitmap.res[3] ;
 wire \vgatest.bitmapColAddr[10] ;
 wire \vgatest.bitmapColAddr[11] ;
 wire \vgatest.bitmapColAddr[12] ;
 wire \vgatest.bitmapColAddr[13] ;
 wire \vgatest.bitmapColAddr[14] ;
 wire \vgatest.bitmapColAddr[2] ;
 wire \vgatest.bitmapColAddr[3] ;
 wire \vgatest.bitmapColAddr[4] ;
 wire \vgatest.bitmapColAddr[5] ;
 wire \vgatest.bitmapColAddr[6] ;
 wire \vgatest.bitmapColAddr[7] ;
 wire \vgatest.bitmapColAddr[8] ;
 wire \vgatest.bitmapColAddr[9] ;
 wire \vgatest.framecounter[0] ;
 wire \vgatest.framecounter[1] ;
 wire \vgatest.framecounter[2] ;
 wire \vgatest.framecounter[3] ;
 wire \vgatest.framecounter[4] ;
 wire \vgatest.framecounter[5] ;
 wire \vgatest.hcounter[0] ;
 wire \vgatest.hcounter[1] ;
 wire \vgatest.hcounter[2] ;
 wire \vgatest.hcounter[3] ;
 wire \vgatest.hcounter[4] ;
 wire \vgatest.hcounter[5] ;
 wire \vgatest.hcounter[6] ;
 wire \vgatest.hcounter[7] ;
 wire \vgatest.hcounter[8] ;
 wire \vgatest.hcounter[9] ;
 wire \vgatest.vcounter[0] ;
 wire \vgatest.vcounter[1] ;
 wire \vgatest.vcounter[2] ;
 wire \vgatest.vcounter[3] ;
 wire \vgatest.vcounter[4] ;
 wire \vgatest.vcounter[5] ;
 wire \vgatest.vcounter[6] ;
 wire \vgatest.vcounter[7] ;
 wire \vgatest.vcounter[8] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0107_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(_1639_));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(_1639_));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(_1660_));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(_1677_));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(_1677_));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(_1677_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(_1709_));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(_1722_));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(_1722_));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(_1722_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(_1755_));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(_1760_));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(_1768_));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(_1890_));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(_1915_));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(_1921_));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(_1921_));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(_1951_));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(_1951_));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(_1951_));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(_1951_));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(_1992_));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(_1992_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(_2014_));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(_0086_));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_0499_));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(_0260_));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(_0309_));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(_0497_));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(_0505_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_0509_));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(_0530_));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0107_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_0593_));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(_1115_));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(_1267_));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(_1267_));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(_1285_));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(_1293_));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(_1294_));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(_1305_));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(_1305_));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(_1397_));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(_1408_));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(_1420_));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(_1440_));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(_1532_));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(_1649_));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(_1651_));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_0757_));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(_1812_));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(_1812_));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(_1890_));
 sky130_fd_sc_hd__diode_2 ANTENNA_268 (.DIODE(_1921_));
 sky130_fd_sc_hd__diode_2 ANTENNA_269 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA_270 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA_271 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA_272 (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA_273 (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA_274 (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA_275 (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA_276 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_277 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_278 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_279 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA_280 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_281 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_282 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_283 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_284 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_285 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_286 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_287 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_288 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_289 (.DIODE(_0086_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA_290 (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA_291 (.DIODE(_0499_));
 sky130_fd_sc_hd__diode_2 ANTENNA_292 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA_293 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA_294 (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA_295 (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA_296 (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA_297 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA_298 (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA_299 (.DIODE(_1395_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0139_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA_300 (.DIODE(_1440_));
 sky130_fd_sc_hd__diode_2 ANTENNA_301 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA_302 (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA_303 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA_304 (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA_305 (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA_306 (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA_307 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA_308 (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_309 (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA_310 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA_311 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA_312 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA_313 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA_314 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA_315 (.DIODE(_1890_));
 sky130_fd_sc_hd__diode_2 ANTENNA_316 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA_317 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_318 (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA_319 (.DIODE(_1395_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA_320 (.DIODE(_1440_));
 sky130_fd_sc_hd__diode_2 ANTENNA_321 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_322 (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA_323 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_1288_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_1290_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_1292_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_1342_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_1366_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_0263_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(_1421_));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(_1440_));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(_1507_));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(_1550_));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(_1577_));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(_1583_));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(_1631_));
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _2038_ (.A(\vgatest.bitmapColAddr[14] ),
    .Y(_2026_));
 sky130_fd_sc_hd__inv_2 _2039_ (.A(\vgatest.bitmapColAddr[13] ),
    .Y(_2037_));
 sky130_fd_sc_hd__inv_2 _2040_ (.A(\vgatest.bitmapColAddr[12] ),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _2041_ (.A(\vgatest.bitmapColAddr[9] ),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _2042_ (.A(\vgatest.vcounter[6] ),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _2043_ (.A(\vgatest.vcounter[1] ),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _2044_ (.A(\vgatest.hcounter[5] ),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _2045_ (.A(net278),
    .Y(_0116_));
 sky130_fd_sc_hd__clkinv_2 _2046_ (.A(net1),
    .Y(_0127_));
 sky130_fd_sc_hd__nor2_1 _2047_ (.A(\vgatest.vcounter[1] ),
    .B(\vgatest.vcounter[0] ),
    .Y(_0138_));
 sky130_fd_sc_hd__and4_1 _2048_ (.A(\vgatest.vcounter[8] ),
    .B(\vgatest.vcounter[7] ),
    .C(_0083_),
    .D(\vgatest.vcounter[4] ),
    .X(_0149_));
 sky130_fd_sc_hd__xnor2_1 _2049_ (.A(\vgatest.vcounter[2] ),
    .B(_0138_),
    .Y(_0160_));
 sky130_fd_sc_hd__or4bb_4 _2050_ (.A(\vgatest.vcounter[5] ),
    .B(\vgatest.vcounter[3] ),
    .C_N(_0149_),
    .D_N(_0160_),
    .X(net12));
 sky130_fd_sc_hd__and4b_1 _2051_ (.A_N(\vgatest.hcounter[8] ),
    .B(\vgatest.hcounter[9] ),
    .C(\vgatest.hcounter[6] ),
    .D(\vgatest.hcounter[7] ),
    .X(_0181_));
 sky130_fd_sc_hd__o21a_1 _2052_ (.A1(\vgatest.hcounter[4] ),
    .A2(\vgatest.hcounter[5] ),
    .B1(_0181_),
    .X(_0191_));
 sky130_fd_sc_hd__nand2_1 _2053_ (.A(\vgatest.hcounter[8] ),
    .B(\vgatest.hcounter[9] ),
    .Y(_0202_));
 sky130_fd_sc_hd__o2111ai_2 _2054_ (.A1(\vgatest.hcounter[3] ),
    .A2(\vgatest.hcounter[2] ),
    .B1(\vgatest.hcounter[4] ),
    .C1(\vgatest.hcounter[5] ),
    .D1(_0191_),
    .Y(_0213_));
 sky130_fd_sc_hd__a41o_1 _2055_ (.A1(\vgatest.hcounter[3] ),
    .A2(\vgatest.hcounter[2] ),
    .A3(\vgatest.hcounter[4] ),
    .A4(\vgatest.hcounter[5] ),
    .B1(_0202_),
    .X(_0224_));
 sky130_fd_sc_hd__o31a_1 _2056_ (.A1(\vgatest.hcounter[6] ),
    .A2(\vgatest.hcounter[7] ),
    .A3(_0224_),
    .B1(_0213_),
    .X(net11));
 sky130_fd_sc_hd__and2_1 _2057_ (.A(\vgatest.bitmapColAddr[3] ),
    .B(\vgatest.hcounter[5] ),
    .X(_0244_));
 sky130_fd_sc_hd__xor2_4 _2058_ (.A(\vgatest.bitmapColAddr[3] ),
    .B(\vgatest.hcounter[5] ),
    .X(_0255_));
 sky130_fd_sc_hd__and2_4 _2059_ (.A(\vgatest.bitmapColAddr[2] ),
    .B(\vgatest.hcounter[4] ),
    .X(_0266_));
 sky130_fd_sc_hd__nand2_2 _2060_ (.A(_0255_),
    .B(_0266_),
    .Y(_0277_));
 sky130_fd_sc_hd__a21o_4 _2061_ (.A1(_0255_),
    .A2(_0266_),
    .B1(_0244_),
    .X(_0288_));
 sky130_fd_sc_hd__and2_1 _2062_ (.A(\vgatest.bitmapColAddr[4] ),
    .B(\vgatest.hcounter[6] ),
    .X(_0299_));
 sky130_fd_sc_hd__xor2_4 _2063_ (.A(\vgatest.bitmapColAddr[4] ),
    .B(\vgatest.hcounter[6] ),
    .X(_0310_));
 sky130_fd_sc_hd__or2_2 _2064_ (.A(\vgatest.bitmapColAddr[5] ),
    .B(\vgatest.hcounter[7] ),
    .X(_0321_));
 sky130_fd_sc_hd__xor2_4 _2065_ (.A(\vgatest.bitmapColAddr[5] ),
    .B(\vgatest.hcounter[7] ),
    .X(_0332_));
 sky130_fd_sc_hd__and2_2 _2066_ (.A(_0310_),
    .B(_0332_),
    .X(_0343_));
 sky130_fd_sc_hd__xor2_4 _2067_ (.A(\vgatest.bitmapColAddr[7] ),
    .B(\vgatest.hcounter[9] ),
    .X(_0353_));
 sky130_fd_sc_hd__nand2_1 _2068_ (.A(\vgatest.bitmapColAddr[6] ),
    .B(\vgatest.hcounter[8] ),
    .Y(_0364_));
 sky130_fd_sc_hd__nor2_1 _2069_ (.A(\vgatest.bitmapColAddr[6] ),
    .B(\vgatest.hcounter[8] ),
    .Y(_0375_));
 sky130_fd_sc_hd__xor2_4 _2070_ (.A(\vgatest.bitmapColAddr[6] ),
    .B(\vgatest.hcounter[8] ),
    .X(_0386_));
 sky130_fd_sc_hd__nand4_4 _2071_ (.A(_0288_),
    .B(_0343_),
    .C(_0353_),
    .D(_0386_),
    .Y(_0397_));
 sky130_fd_sc_hd__a22o_2 _2072_ (.A1(\vgatest.bitmapColAddr[4] ),
    .A2(\vgatest.hcounter[6] ),
    .B1(\vgatest.hcounter[7] ),
    .B2(\vgatest.bitmapColAddr[5] ),
    .X(_0408_));
 sky130_fd_sc_hd__a22o_1 _2073_ (.A1(\vgatest.bitmapColAddr[6] ),
    .A2(\vgatest.hcounter[8] ),
    .B1(\vgatest.hcounter[9] ),
    .B2(\vgatest.bitmapColAddr[7] ),
    .X(_0418_));
 sky130_fd_sc_hd__a31o_1 _2074_ (.A1(_0321_),
    .A2(_0386_),
    .A3(_0408_),
    .B1(_0418_),
    .X(_0429_));
 sky130_fd_sc_hd__o21ai_4 _2075_ (.A1(\vgatest.bitmapColAddr[7] ),
    .A2(\vgatest.hcounter[9] ),
    .B1(_0429_),
    .Y(_0440_));
 sky130_fd_sc_hd__a21boi_4 _2076_ (.A1(_0397_),
    .A2(_0440_),
    .B1_N(\vgatest.bitmapColAddr[8] ),
    .Y(_0451_));
 sky130_fd_sc_hd__a21bo_2 _2077_ (.A1(_0397_),
    .A2(_0440_),
    .B1_N(\vgatest.bitmapColAddr[8] ),
    .X(_0462_));
 sky130_fd_sc_hd__nand2_4 _2078_ (.A(\vgatest.bitmapColAddr[9] ),
    .B(\vgatest.bitmapColAddr[8] ),
    .Y(_0473_));
 sky130_fd_sc_hd__a21oi_4 _2079_ (.A1(_0397_),
    .A2(_0440_),
    .B1(_0473_),
    .Y(_0484_));
 sky130_fd_sc_hd__nand2_1 _2080_ (.A(net276),
    .B(\vgatest.bitmapColAddr[10] ),
    .Y(_0495_));
 sky130_fd_sc_hd__and3_1 _2081_ (.A(net276),
    .B(\vgatest.bitmapColAddr[10] ),
    .C(_0484_),
    .X(_0506_));
 sky130_fd_sc_hd__a211o_4 _2082_ (.A1(_0397_),
    .A2(_0440_),
    .B1(_0473_),
    .C1(_0495_),
    .X(_0517_));
 sky130_fd_sc_hd__a2111o_4 _2083_ (.A1(_0397_),
    .A2(_0440_),
    .B1(_0473_),
    .C1(_0495_),
    .D1(_0061_),
    .X(_0528_));
 sky130_fd_sc_hd__xnor2_4 _2084_ (.A(\vgatest.bitmapColAddr[12] ),
    .B(_0517_),
    .Y(_0539_));
 sky130_fd_sc_hd__or2_4 _2085_ (.A(_2037_),
    .B(_0528_),
    .X(_0550_));
 sky130_fd_sc_hd__xnor2_4 _2086_ (.A(_2037_),
    .B(_0528_),
    .Y(_0561_));
 sky130_fd_sc_hd__nor2_2 _2087_ (.A(_0539_),
    .B(_0561_),
    .Y(_0572_));
 sky130_fd_sc_hd__or2_2 _2088_ (.A(_0539_),
    .B(_0561_),
    .X(_0583_));
 sky130_fd_sc_hd__xnor2_4 _2089_ (.A(_2026_),
    .B(_0550_),
    .Y(_0594_));
 sky130_fd_sc_hd__xnor2_4 _2090_ (.A(\vgatest.bitmapColAddr[14] ),
    .B(_0550_),
    .Y(_0605_));
 sky130_fd_sc_hd__xor2_4 _2091_ (.A(\vgatest.bitmapColAddr[10] ),
    .B(_0484_),
    .X(_0616_));
 sky130_fd_sc_hd__and4_2 _2092_ (.A(net276),
    .B(_0572_),
    .C(_0594_),
    .D(_0616_),
    .X(_0627_));
 sky130_fd_sc_hd__nor2_8 _2093_ (.A(\vgatest.bitmapColAddr[2] ),
    .B(\vgatest.hcounter[4] ),
    .Y(_0638_));
 sky130_fd_sc_hd__nor2_8 _2094_ (.A(_0266_),
    .B(_0638_),
    .Y(_0649_));
 sky130_fd_sc_hd__or2_4 _2095_ (.A(_0255_),
    .B(_0266_),
    .X(_0660_));
 sky130_fd_sc_hd__nand2_2 _2096_ (.A(_0277_),
    .B(_0660_),
    .Y(_0671_));
 sky130_fd_sc_hd__nor2_4 _2097_ (.A(_0649_),
    .B(_0671_),
    .Y(_0682_));
 sky130_fd_sc_hd__or2_1 _2098_ (.A(_0649_),
    .B(_0671_),
    .X(_0693_));
 sky130_fd_sc_hd__xor2_4 _2099_ (.A(_0288_),
    .B(_0310_),
    .X(_0704_));
 sky130_fd_sc_hd__xnor2_1 _2100_ (.A(_0288_),
    .B(_0310_),
    .Y(_0715_));
 sky130_fd_sc_hd__a21oi_4 _2101_ (.A1(_0288_),
    .A2(_0310_),
    .B1(_0299_),
    .Y(_0726_));
 sky130_fd_sc_hd__xor2_2 _2102_ (.A(_0332_),
    .B(_0726_),
    .X(_0737_));
 sky130_fd_sc_hd__xnor2_4 _2103_ (.A(_0332_),
    .B(_0726_),
    .Y(_0748_));
 sky130_fd_sc_hd__and3_2 _2104_ (.A(_0682_),
    .B(net272),
    .C(net267),
    .X(_0759_));
 sky130_fd_sc_hd__or3_4 _2105_ (.A(_0693_),
    .B(net270),
    .C(net265),
    .X(_0770_));
 sky130_fd_sc_hd__and3b_2 _2106_ (.A_N(\vgatest.bitmapColAddr[8] ),
    .B(_0397_),
    .C(_0440_),
    .X(_0781_));
 sky130_fd_sc_hd__nand3b_4 _2107_ (.A_N(\vgatest.bitmapColAddr[8] ),
    .B(_0397_),
    .C(_0440_),
    .Y(_0792_));
 sky130_fd_sc_hd__nor2_4 _2108_ (.A(_0451_),
    .B(_0781_),
    .Y(_0803_));
 sky130_fd_sc_hd__nand2_4 _2109_ (.A(_0462_),
    .B(_0792_),
    .Y(_0814_));
 sky130_fd_sc_hd__xnor2_4 _2110_ (.A(_0072_),
    .B(_0451_),
    .Y(_0825_));
 sky130_fd_sc_hd__xnor2_4 _2111_ (.A(\vgatest.bitmapColAddr[9] ),
    .B(_0451_),
    .Y(_0836_));
 sky130_fd_sc_hd__a22oi_4 _2112_ (.A1(_0288_),
    .A2(_0343_),
    .B1(_0408_),
    .B2(_0321_),
    .Y(_0847_));
 sky130_fd_sc_hd__xnor2_4 _2113_ (.A(_0386_),
    .B(_0847_),
    .Y(_0858_));
 sky130_fd_sc_hd__xor2_2 _2114_ (.A(_0386_),
    .B(_0847_),
    .X(_0869_));
 sky130_fd_sc_hd__o21a_4 _2115_ (.A1(_0375_),
    .A2(_0847_),
    .B1(_0364_),
    .X(_0880_));
 sky130_fd_sc_hd__xor2_4 _2116_ (.A(_0353_),
    .B(_0880_),
    .X(_0891_));
 sky130_fd_sc_hd__xnor2_1 _2117_ (.A(_0353_),
    .B(_0880_),
    .Y(_0902_));
 sky130_fd_sc_hd__and4_4 _2118_ (.A(_0814_),
    .B(_0825_),
    .C(net262),
    .D(net228),
    .X(_0913_));
 sky130_fd_sc_hd__or4_2 _2119_ (.A(_0803_),
    .B(_0836_),
    .C(net253),
    .D(net237),
    .X(_0924_));
 sky130_fd_sc_hd__nor2_8 _2120_ (.A(net241),
    .B(net126),
    .Y(_0935_));
 sky130_fd_sc_hd__and3_4 _2121_ (.A(\vgatest.bitmapColAddr[9] ),
    .B(_0462_),
    .C(_0792_),
    .X(_0946_));
 sky130_fd_sc_hd__and3_4 _2122_ (.A(net249),
    .B(net224),
    .C(net216),
    .X(_0957_));
 sky130_fd_sc_hd__or3b_4 _2123_ (.A(net262),
    .B(net237),
    .C_N(_0946_),
    .X(_0968_));
 sky130_fd_sc_hd__nor2_8 _2124_ (.A(net241),
    .B(_0968_),
    .Y(_0979_));
 sky130_fd_sc_hd__and3_4 _2125_ (.A(_0682_),
    .B(net272),
    .C(net264),
    .X(_0990_));
 sky130_fd_sc_hd__or3_4 _2126_ (.A(_0693_),
    .B(net270),
    .C(net266),
    .X(_1001_));
 sky130_fd_sc_hd__and4_4 _2127_ (.A(_0814_),
    .B(_0825_),
    .C(net253),
    .D(net228),
    .X(_1012_));
 sky130_fd_sc_hd__or4_4 _2128_ (.A(_0803_),
    .B(_0836_),
    .C(net262),
    .D(net237),
    .X(_1023_));
 sky130_fd_sc_hd__nor2_8 _2129_ (.A(net206),
    .B(net122),
    .Y(_1034_));
 sky130_fd_sc_hd__nor2_8 _2130_ (.A(_0638_),
    .B(_0660_),
    .Y(_1045_));
 sky130_fd_sc_hd__or2_1 _2131_ (.A(_0638_),
    .B(_0660_),
    .X(_1056_));
 sky130_fd_sc_hd__and3_4 _2132_ (.A(net270),
    .B(net264),
    .C(_1045_),
    .X(_1067_));
 sky130_fd_sc_hd__or3_4 _2133_ (.A(net273),
    .B(net266),
    .C(_1056_),
    .X(_1078_));
 sky130_fd_sc_hd__and4_4 _2134_ (.A(_0814_),
    .B(_0825_),
    .C(net253),
    .D(net237),
    .X(_1089_));
 sky130_fd_sc_hd__or4_4 _2135_ (.A(_0803_),
    .B(_0836_),
    .C(net262),
    .D(net228),
    .X(_1100_));
 sky130_fd_sc_hd__nor2_2 _2136_ (.A(net201),
    .B(net116),
    .Y(_1111_));
 sky130_fd_sc_hd__and2_4 _2137_ (.A(_0255_),
    .B(_0649_),
    .X(_1121_));
 sky130_fd_sc_hd__nand2_1 _2138_ (.A(_0255_),
    .B(_0649_),
    .Y(_1131_));
 sky130_fd_sc_hd__nor2_8 _2139_ (.A(net272),
    .B(net264),
    .Y(_1138_));
 sky130_fd_sc_hd__and3_4 _2140_ (.A(net271),
    .B(net267),
    .C(_1121_),
    .X(_1146_));
 sky130_fd_sc_hd__nand2_2 _2141_ (.A(_1121_),
    .B(_1138_),
    .Y(_1155_));
 sky130_fd_sc_hd__nor2_8 _2142_ (.A(_0968_),
    .B(net115),
    .Y(_1163_));
 sky130_fd_sc_hd__a21oi_4 _2143_ (.A1(_0277_),
    .A2(_0660_),
    .B1(_0649_),
    .Y(_1172_));
 sky130_fd_sc_hd__a21o_1 _2144_ (.A1(_0277_),
    .A2(_0660_),
    .B1(_0649_),
    .X(_1181_));
 sky130_fd_sc_hd__and3_2 _2145_ (.A(net270),
    .B(net264),
    .C(_1172_),
    .X(_1191_));
 sky130_fd_sc_hd__or3_4 _2146_ (.A(net273),
    .B(net266),
    .C(_1181_),
    .X(_1197_));
 sky130_fd_sc_hd__and4_4 _2147_ (.A(_0814_),
    .B(_0836_),
    .C(net253),
    .D(net228),
    .X(_1205_));
 sky130_fd_sc_hd__or4_2 _2148_ (.A(_0803_),
    .B(_0825_),
    .C(net262),
    .D(net237),
    .X(_1213_));
 sky130_fd_sc_hd__nor2_8 _2149_ (.A(net191),
    .B(net109),
    .Y(_1222_));
 sky130_fd_sc_hd__and3_4 _2150_ (.A(net272),
    .B(net267),
    .C(_1121_),
    .X(_1230_));
 sky130_fd_sc_hd__or3_4 _2151_ (.A(net271),
    .B(net265),
    .C(_1131_),
    .X(_1236_));
 sky130_fd_sc_hd__nor2_8 _2152_ (.A(net109),
    .B(net185),
    .Y(_1243_));
 sky130_fd_sc_hd__a21oi_2 _2153_ (.A1(net190),
    .A2(net185),
    .B1(net110),
    .Y(_1249_));
 sky130_fd_sc_hd__and3_2 _2154_ (.A(net270),
    .B(_0737_),
    .C(_1045_),
    .X(_1250_));
 sky130_fd_sc_hd__nand2_4 _2155_ (.A(_1045_),
    .B(_1138_),
    .Y(_1251_));
 sky130_fd_sc_hd__and4_4 _2156_ (.A(_0814_),
    .B(_0836_),
    .C(net253),
    .D(net237),
    .X(_1252_));
 sky130_fd_sc_hd__or4_4 _2157_ (.A(_0803_),
    .B(_0825_),
    .C(net262),
    .D(net228),
    .X(_1253_));
 sky130_fd_sc_hd__nor2_8 _2158_ (.A(net107),
    .B(net102),
    .Y(_1254_));
 sky130_fd_sc_hd__and3_4 _2159_ (.A(net270),
    .B(net266),
    .C(_1172_),
    .X(_1255_));
 sky130_fd_sc_hd__nand2_1 _2160_ (.A(_1138_),
    .B(_1172_),
    .Y(_1256_));
 sky130_fd_sc_hd__nor2_8 _2161_ (.A(net104),
    .B(net100),
    .Y(_1257_));
 sky130_fd_sc_hd__a21oi_4 _2162_ (.A1(net106),
    .A2(net100),
    .B1(net103),
    .Y(_1258_));
 sky130_fd_sc_hd__or4_1 _2163_ (.A(_1111_),
    .B(_1163_),
    .C(_1249_),
    .D(_1258_),
    .X(_1259_));
 sky130_fd_sc_hd__o41a_1 _2164_ (.A1(_0935_),
    .A2(_0979_),
    .A3(_1034_),
    .A4(_1259_),
    .B1(net66),
    .X(_1260_));
 sky130_fd_sc_hd__and2_1 _2165_ (.A(\vgatest.bitmapColAddr[13] ),
    .B(_0539_),
    .X(_1261_));
 sky130_fd_sc_hd__nand2_4 _2166_ (.A(\vgatest.bitmapColAddr[13] ),
    .B(_0539_),
    .Y(_1262_));
 sky130_fd_sc_hd__and4_4 _2167_ (.A(net276),
    .B(_0594_),
    .C(_0616_),
    .D(_1261_),
    .X(_1263_));
 sky130_fd_sc_hd__nor2_1 _2168_ (.A(net208),
    .B(net116),
    .Y(_1264_));
 sky130_fd_sc_hd__and3_4 _2169_ (.A(net272),
    .B(net264),
    .C(_1045_),
    .X(_1265_));
 sky130_fd_sc_hd__or3_4 _2170_ (.A(net271),
    .B(net266),
    .C(_1056_),
    .X(_1266_));
 sky130_fd_sc_hd__nor2_8 _2171_ (.A(net116),
    .B(net176),
    .Y(_1267_));
 sky130_fd_sc_hd__a21oi_4 _2172_ (.A1(net207),
    .A2(net174),
    .B1(net118),
    .Y(_1268_));
 sky130_fd_sc_hd__and3_4 _2173_ (.A(net272),
    .B(net264),
    .C(_1121_),
    .X(_1269_));
 sky130_fd_sc_hd__or3_2 _2174_ (.A(net271),
    .B(net266),
    .C(_1131_),
    .X(_1270_));
 sky130_fd_sc_hd__nor2_1 _2175_ (.A(net116),
    .B(net171),
    .Y(_1271_));
 sky130_fd_sc_hd__and4_4 _2176_ (.A(_0814_),
    .B(_0825_),
    .C(net262),
    .D(net237),
    .X(_1272_));
 sky130_fd_sc_hd__or4_4 _2177_ (.A(_0803_),
    .B(_0836_),
    .C(net253),
    .D(net228),
    .X(_1273_));
 sky130_fd_sc_hd__nor2_4 _2178_ (.A(net101),
    .B(net95),
    .Y(_1274_));
 sky130_fd_sc_hd__a22o_1 _2179_ (.A1(net120),
    .A2(net173),
    .B1(net98),
    .B2(net181),
    .X(_1275_));
 sky130_fd_sc_hd__or2_4 _2180_ (.A(_1268_),
    .B(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__and3_4 _2181_ (.A(_0682_),
    .B(net270),
    .C(net264),
    .X(_1277_));
 sky130_fd_sc_hd__or3_4 _2182_ (.A(_0693_),
    .B(net273),
    .C(net266),
    .X(_1278_));
 sky130_fd_sc_hd__nor2_1 _2183_ (.A(net102),
    .B(net165),
    .Y(_1279_));
 sky130_fd_sc_hd__nor2_8 _2184_ (.A(net201),
    .B(net102),
    .Y(_1280_));
 sky130_fd_sc_hd__a21oi_4 _2185_ (.A1(net199),
    .A2(net166),
    .B1(net104),
    .Y(_1281_));
 sky130_fd_sc_hd__nor2_1 _2186_ (.A(net186),
    .B(net102),
    .Y(_1282_));
 sky130_fd_sc_hd__nor2_8 _2187_ (.A(net192),
    .B(net102),
    .Y(_1283_));
 sky130_fd_sc_hd__a21oi_2 _2188_ (.A1(net190),
    .A2(net185),
    .B1(net104),
    .Y(_1284_));
 sky130_fd_sc_hd__or2_4 _2189_ (.A(_1281_),
    .B(_1284_),
    .X(_1285_));
 sky130_fd_sc_hd__and3_4 _2190_ (.A(_0072_),
    .B(_0462_),
    .C(_0792_),
    .X(_1286_));
 sky130_fd_sc_hd__or3_4 _2191_ (.A(\vgatest.bitmapColAddr[9] ),
    .B(_0451_),
    .C(_0781_),
    .X(_1287_));
 sky130_fd_sc_hd__and3_4 _2192_ (.A(net245),
    .B(net221),
    .C(net157),
    .X(_1288_));
 sky130_fd_sc_hd__or3_4 _2193_ (.A(net263),
    .B(net239),
    .C(_1287_),
    .X(_1289_));
 sky130_fd_sc_hd__and4_4 _2194_ (.A(net248),
    .B(net223),
    .C(net180),
    .D(net159),
    .X(_1290_));
 sky130_fd_sc_hd__and4_4 _2195_ (.A(net247),
    .B(net222),
    .C(net196),
    .D(net157),
    .X(_1291_));
 sky130_fd_sc_hd__or2_4 _2196_ (.A(_1290_),
    .B(_1291_),
    .X(_1292_));
 sky130_fd_sc_hd__and4_4 _2197_ (.A(net248),
    .B(net225),
    .C(net182),
    .D(net158),
    .X(_1293_));
 sky130_fd_sc_hd__and3_4 _2198_ (.A(_0682_),
    .B(net270),
    .C(net267),
    .X(_1294_));
 sky130_fd_sc_hd__nand2_2 _2199_ (.A(_0682_),
    .B(_1138_),
    .Y(_1295_));
 sky130_fd_sc_hd__and4_4 _2200_ (.A(net250),
    .B(net226),
    .C(net162),
    .D(net155),
    .X(_1296_));
 sky130_fd_sc_hd__or2_2 _2201_ (.A(net94),
    .B(_1296_),
    .X(_1297_));
 sky130_fd_sc_hd__or2_1 _2202_ (.A(_1292_),
    .B(_1297_),
    .X(_1298_));
 sky130_fd_sc_hd__and4_2 _2203_ (.A(_0814_),
    .B(_0836_),
    .C(net262),
    .D(net228),
    .X(_1299_));
 sky130_fd_sc_hd__or4_2 _2204_ (.A(_0803_),
    .B(_0825_),
    .C(net254),
    .D(net237),
    .X(_1300_));
 sky130_fd_sc_hd__nor2_4 _2205_ (.A(net185),
    .B(net85),
    .Y(_1301_));
 sky130_fd_sc_hd__and3_2 _2206_ (.A(net272),
    .B(net267),
    .C(_1172_),
    .X(_1302_));
 sky130_fd_sc_hd__or3_4 _2207_ (.A(net271),
    .B(net265),
    .C(_1181_),
    .X(_1303_));
 sky130_fd_sc_hd__nor2_1 _2208_ (.A(net87),
    .B(net150),
    .Y(_1304_));
 sky130_fd_sc_hd__a21oi_4 _2209_ (.A1(_1236_),
    .A2(net148),
    .B1(net86),
    .Y(_1305_));
 sky130_fd_sc_hd__and3_2 _2210_ (.A(net273),
    .B(net266),
    .C(_1045_),
    .X(_1306_));
 sky130_fd_sc_hd__or3_4 _2211_ (.A(net271),
    .B(net265),
    .C(_1056_),
    .X(_1307_));
 sky130_fd_sc_hd__nor2_8 _2212_ (.A(net87),
    .B(net142),
    .Y(_1308_));
 sky130_fd_sc_hd__nor2_4 _2213_ (.A(net241),
    .B(net87),
    .Y(_1309_));
 sky130_fd_sc_hd__o41a_2 _2214_ (.A1(net243),
    .A2(net189),
    .A3(net153),
    .A4(net146),
    .B1(net89),
    .X(_1310_));
 sky130_fd_sc_hd__or4_2 _2215_ (.A(_1276_),
    .B(_1285_),
    .C(_1298_),
    .D(_1310_),
    .X(_1311_));
 sky130_fd_sc_hd__a21o_1 _2216_ (.A1(\vgatest.bitmapColAddr[10] ),
    .A2(_0484_),
    .B1(net276),
    .X(_1312_));
 sky130_fd_sc_hd__a21o_4 _2217_ (.A1(_0517_),
    .A2(_1312_),
    .B1(_0616_),
    .X(_1313_));
 sky130_fd_sc_hd__nor3_2 _2218_ (.A(_0605_),
    .B(_1262_),
    .C(_1313_),
    .Y(_1314_));
 sky130_fd_sc_hd__nor2_2 _2219_ (.A(net107),
    .B(net95),
    .Y(_1315_));
 sky130_fd_sc_hd__nor2_2 _2220_ (.A(net97),
    .B(net150),
    .Y(_1316_));
 sky130_fd_sc_hd__and3_2 _2221_ (.A(net257),
    .B(net221),
    .C(net214),
    .X(_1317_));
 sky130_fd_sc_hd__or3b_4 _2222_ (.A(net250),
    .B(net236),
    .C_N(net219),
    .X(_1318_));
 sky130_fd_sc_hd__and4_4 _2223_ (.A(net261),
    .B(net226),
    .C(net219),
    .D(net154),
    .X(_1319_));
 sky130_fd_sc_hd__nor2_4 _2224_ (.A(net107),
    .B(_1318_),
    .Y(_1320_));
 sky130_fd_sc_hd__o2111a_4 _2225_ (.A1(net183),
    .A2(net154),
    .B1(net260),
    .C1(net225),
    .D1(net217),
    .X(_1321_));
 sky130_fd_sc_hd__nor2_8 _2226_ (.A(net186),
    .B(net95),
    .Y(_1322_));
 sky130_fd_sc_hd__nor2_4 _2227_ (.A(net115),
    .B(_1318_),
    .Y(_1323_));
 sky130_fd_sc_hd__and4_4 _2228_ (.A(net257),
    .B(net221),
    .C(net213),
    .D(net180),
    .X(_1324_));
 sky130_fd_sc_hd__a21oi_2 _2229_ (.A1(net115),
    .A2(net101),
    .B1(_1318_),
    .Y(_1325_));
 sky130_fd_sc_hd__and3_4 _2230_ (.A(net273),
    .B(net265),
    .C(_1172_),
    .X(_1326_));
 sky130_fd_sc_hd__or3_4 _2231_ (.A(net271),
    .B(net266),
    .C(_1181_),
    .X(_1327_));
 sky130_fd_sc_hd__and4_4 _2232_ (.A(net249),
    .B(net224),
    .C(net216),
    .D(net138),
    .X(_1328_));
 sky130_fd_sc_hd__and3_4 _2233_ (.A(net270),
    .B(net265),
    .C(_1121_),
    .X(_1329_));
 sky130_fd_sc_hd__or3_4 _2234_ (.A(net273),
    .B(net266),
    .C(_1131_),
    .X(_1330_));
 sky130_fd_sc_hd__and4_4 _2235_ (.A(net249),
    .B(net224),
    .C(net217),
    .D(net133),
    .X(_1331_));
 sky130_fd_sc_hd__or4_4 _2236_ (.A(_1308_),
    .B(_1315_),
    .C(_1322_),
    .D(_1325_),
    .X(_1332_));
 sky130_fd_sc_hd__or3_1 _2237_ (.A(_1316_),
    .B(net82),
    .C(_1331_),
    .X(_1333_));
 sky130_fd_sc_hd__or4_1 _2238_ (.A(_1271_),
    .B(_1321_),
    .C(_1332_),
    .D(_1333_),
    .X(_1334_));
 sky130_fd_sc_hd__a221o_1 _2239_ (.A1(net63),
    .A2(_1311_),
    .B1(net59),
    .B2(_1334_),
    .C1(_1260_),
    .X(_1335_));
 sky130_fd_sc_hd__or4b_4 _2240_ (.A(\vgatest.bitmapColAddr[14] ),
    .B(_0506_),
    .C(_0616_),
    .D_N(_1312_),
    .X(_1336_));
 sky130_fd_sc_hd__and2_1 _2241_ (.A(_2037_),
    .B(_0539_),
    .X(_1337_));
 sky130_fd_sc_hd__and2b_1 _2242_ (.A_N(_1336_),
    .B(_1337_),
    .X(_1338_));
 sky130_fd_sc_hd__and4_4 _2243_ (.A(net257),
    .B(net221),
    .C(net213),
    .D(net151),
    .X(_1339_));
 sky130_fd_sc_hd__and3_4 _2244_ (.A(net245),
    .B(net232),
    .C(net214),
    .X(_1340_));
 sky130_fd_sc_hd__and2_2 _2245_ (.A(net242),
    .B(_1340_),
    .X(_1341_));
 sky130_fd_sc_hd__and4_4 _2246_ (.A(net245),
    .B(net232),
    .C(net213),
    .D(net187),
    .X(_1342_));
 sky130_fd_sc_hd__o2111a_4 _2247_ (.A1(net243),
    .A2(net189),
    .B1(net220),
    .C1(net238),
    .D1(net251),
    .X(_1343_));
 sky130_fd_sc_hd__a211o_2 _2248_ (.A1(net196),
    .A2(net83),
    .B1(_1339_),
    .C1(_1343_),
    .X(_1344_));
 sky130_fd_sc_hd__nor2_8 _2249_ (.A(net201),
    .B(_1318_),
    .Y(_1345_));
 sky130_fd_sc_hd__o2111a_1 _2250_ (.A1(net202),
    .A2(net193),
    .B1(net260),
    .C1(net225),
    .D1(net217),
    .X(_1346_));
 sky130_fd_sc_hd__and4_4 _2251_ (.A(net256),
    .B(net222),
    .C(net212),
    .D(net144),
    .X(_1347_));
 sky130_fd_sc_hd__a211o_1 _2252_ (.A1(net105),
    .A2(net138),
    .B1(_1346_),
    .C1(_1347_),
    .X(_1348_));
 sky130_fd_sc_hd__nor2_4 _2253_ (.A(_0968_),
    .B(net176),
    .Y(_1349_));
 sky130_fd_sc_hd__nor2_2 _2254_ (.A(_1253_),
    .B(net176),
    .Y(_1350_));
 sky130_fd_sc_hd__or4_4 _2255_ (.A(_1319_),
    .B(net82),
    .C(_1349_),
    .D(_1350_),
    .X(_1351_));
 sky130_fd_sc_hd__o31a_1 _2256_ (.A1(_1344_),
    .A2(_1348_),
    .A3(_1351_),
    .B1(net54),
    .X(_1352_));
 sky130_fd_sc_hd__nor2_2 _2257_ (.A(_0583_),
    .B(_1336_),
    .Y(_1353_));
 sky130_fd_sc_hd__and4_4 _2258_ (.A(net257),
    .B(net221),
    .C(net214),
    .D(net172),
    .X(_1354_));
 sky130_fd_sc_hd__a21o_1 _2259_ (.A1(net210),
    .A2(net83),
    .B1(_1354_),
    .X(_1355_));
 sky130_fd_sc_hd__nor2_4 _2260_ (.A(net165),
    .B(_1318_),
    .Y(_1356_));
 sky130_fd_sc_hd__and4_4 _2261_ (.A(net257),
    .B(net223),
    .C(net215),
    .D(net133),
    .X(_1357_));
 sky130_fd_sc_hd__or3_1 _2262_ (.A(_1355_),
    .B(_1356_),
    .C(_1357_),
    .X(_1358_));
 sky130_fd_sc_hd__or3b_4 _2263_ (.A(net252),
    .B(net227),
    .C_N(net220),
    .X(_1359_));
 sky130_fd_sc_hd__and4_4 _2264_ (.A(net257),
    .B(net232),
    .C(net215),
    .D(net151),
    .X(_1360_));
 sky130_fd_sc_hd__a21o_2 _2265_ (.A1(net123),
    .A2(net187),
    .B1(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__nor2_8 _2266_ (.A(net241),
    .B(net121),
    .Y(_1362_));
 sky130_fd_sc_hd__and4_4 _2267_ (.A(net255),
    .B(net230),
    .C(net212),
    .D(net196),
    .X(_1363_));
 sky130_fd_sc_hd__or3_4 _2268_ (.A(_1361_),
    .B(_1362_),
    .C(_1363_),
    .X(_1364_));
 sky130_fd_sc_hd__and4_4 _2269_ (.A(net260),
    .B(net235),
    .C(net216),
    .D(net182),
    .X(_1365_));
 sky130_fd_sc_hd__and4_4 _2270_ (.A(net256),
    .B(net231),
    .C(net212),
    .D(net154),
    .X(_1366_));
 sky130_fd_sc_hd__and4_4 _2271_ (.A(net247),
    .B(net231),
    .C(net212),
    .D(net209),
    .X(_1367_));
 sky130_fd_sc_hd__and4_4 _2272_ (.A(net250),
    .B(net236),
    .C(net216),
    .D(net172),
    .X(_1368_));
 sky130_fd_sc_hd__or2_4 _2273_ (.A(_1367_),
    .B(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__or3_1 _2274_ (.A(_1365_),
    .B(_1366_),
    .C(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__o31a_1 _2275_ (.A1(_1358_),
    .A2(_1364_),
    .A3(_1370_),
    .B1(net52),
    .X(_1371_));
 sky130_fd_sc_hd__and4_4 _2276_ (.A(net276),
    .B(_0594_),
    .C(_0616_),
    .D(_1337_),
    .X(_1372_));
 sky130_fd_sc_hd__nor2_8 _2277_ (.A(net122),
    .B(net175),
    .Y(_1373_));
 sky130_fd_sc_hd__and4_4 _2278_ (.A(net261),
    .B(net235),
    .C(net217),
    .D(net169),
    .X(_1374_));
 sky130_fd_sc_hd__a21o_4 _2279_ (.A1(net124),
    .A2(net179),
    .B1(_1374_),
    .X(_1375_));
 sky130_fd_sc_hd__nor2_8 _2280_ (.A(_1023_),
    .B(net137),
    .Y(_1376_));
 sky130_fd_sc_hd__and4_4 _2281_ (.A(net257),
    .B(net232),
    .C(net214),
    .D(net202),
    .X(_1377_));
 sky130_fd_sc_hd__a21oi_4 _2282_ (.A1(net174),
    .A2(net137),
    .B1(net122),
    .Y(_1378_));
 sky130_fd_sc_hd__o2111a_4 _2283_ (.A1(net204),
    .A2(net168),
    .B1(net263),
    .C1(net238),
    .D1(net220),
    .X(_1379_));
 sky130_fd_sc_hd__nor2_2 _2284_ (.A(net121),
    .B(net143),
    .Y(_1380_));
 sky130_fd_sc_hd__nor2_2 _2285_ (.A(net121),
    .B(net192),
    .Y(_1381_));
 sky130_fd_sc_hd__a21oi_4 _2286_ (.A1(net190),
    .A2(net185),
    .B1(net121),
    .Y(_1382_));
 sky130_fd_sc_hd__or2_4 _2287_ (.A(_1360_),
    .B(_1363_),
    .X(_1383_));
 sky130_fd_sc_hd__or4_1 _2288_ (.A(_1378_),
    .B(_1379_),
    .C(_1382_),
    .D(_1383_),
    .X(_1384_));
 sky130_fd_sc_hd__o31a_1 _2289_ (.A1(_1362_),
    .A2(_1380_),
    .A3(_1384_),
    .B1(net49),
    .X(_1385_));
 sky130_fd_sc_hd__and2b_2 _2290_ (.A_N(net276),
    .B(_0616_),
    .X(_1386_));
 sky130_fd_sc_hd__and3_2 _2291_ (.A(_0594_),
    .B(_1261_),
    .C(_1386_),
    .X(_1387_));
 sky130_fd_sc_hd__and4_4 _2292_ (.A(net242),
    .B(net256),
    .C(net222),
    .D(net212),
    .X(_1388_));
 sky130_fd_sc_hd__or3_4 _2293_ (.A(net254),
    .B(net237),
    .C(_1287_),
    .X(_1389_));
 sky130_fd_sc_hd__and4_4 _2294_ (.A(net261),
    .B(net224),
    .C(net161),
    .D(net144),
    .X(_1390_));
 sky130_fd_sc_hd__and4_4 _2295_ (.A(net255),
    .B(net222),
    .C(net156),
    .D(net154),
    .X(_1391_));
 sky130_fd_sc_hd__a221o_1 _2296_ (.A1(net187),
    .A2(net99),
    .B1(net83),
    .B2(net193),
    .C1(_1354_),
    .X(_1392_));
 sky130_fd_sc_hd__or4_1 _2297_ (.A(_1388_),
    .B(_1390_),
    .C(_1391_),
    .D(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__and4_4 _2298_ (.A(net259),
    .B(net223),
    .C(net218),
    .D(net179),
    .X(_1394_));
 sky130_fd_sc_hd__and4_4 _2299_ (.A(net261),
    .B(net226),
    .C(net219),
    .D(net139),
    .X(_1395_));
 sky130_fd_sc_hd__o41a_4 _2300_ (.A1(net211),
    .A2(net177),
    .A3(net141),
    .A4(net134),
    .B1(net83),
    .X(_1396_));
 sky130_fd_sc_hd__and4_4 _2301_ (.A(net260),
    .B(net235),
    .C(net216),
    .D(net180),
    .X(_1397_));
 sky130_fd_sc_hd__or3_2 _2302_ (.A(_1365_),
    .B(_1369_),
    .C(_1397_),
    .X(_1398_));
 sky130_fd_sc_hd__o31a_1 _2303_ (.A1(_1393_),
    .A2(_1396_),
    .A3(_1398_),
    .B1(net44),
    .X(_1399_));
 sky130_fd_sc_hd__or4_4 _2304_ (.A(_1352_),
    .B(_1371_),
    .C(_1385_),
    .D(_1399_),
    .X(_1400_));
 sky130_fd_sc_hd__and2b_2 _2305_ (.A_N(_0539_),
    .B(_0561_),
    .X(_1401_));
 sky130_fd_sc_hd__nand2b_4 _2306_ (.A_N(_0539_),
    .B(_0561_),
    .Y(_1402_));
 sky130_fd_sc_hd__and3b_4 _2307_ (.A_N(_1313_),
    .B(_1401_),
    .C(_0605_),
    .X(_1403_));
 sky130_fd_sc_hd__or3_4 _2308_ (.A(net263),
    .B(net229),
    .C(_1287_),
    .X(_1404_));
 sky130_fd_sc_hd__nor2_4 _2309_ (.A(net150),
    .B(_1404_),
    .Y(_1405_));
 sky130_fd_sc_hd__and4_4 _2310_ (.A(net250),
    .B(net236),
    .C(net197),
    .D(net162),
    .X(_1406_));
 sky130_fd_sc_hd__o2111a_4 _2311_ (.A1(net198),
    .A2(net152),
    .B1(net163),
    .C1(net251),
    .D1(net238),
    .X(_1407_));
 sky130_fd_sc_hd__and4_4 _2312_ (.A(_0814_),
    .B(_0836_),
    .C(net262),
    .D(net239),
    .X(_1408_));
 sky130_fd_sc_hd__or4_4 _2313_ (.A(_0803_),
    .B(_0825_),
    .C(net253),
    .D(net229),
    .X(_1409_));
 sky130_fd_sc_hd__nor2_8 _2314_ (.A(net142),
    .B(net77),
    .Y(_1410_));
 sky130_fd_sc_hd__nor2_4 _2315_ (.A(net241),
    .B(net80),
    .Y(_1411_));
 sky130_fd_sc_hd__or3_2 _2316_ (.A(_1407_),
    .B(_1410_),
    .C(_1411_),
    .X(_1412_));
 sky130_fd_sc_hd__and4_4 _2317_ (.A(net247),
    .B(net222),
    .C(net172),
    .D(net157),
    .X(_1413_));
 sky130_fd_sc_hd__and4_4 _2318_ (.A(net248),
    .B(net225),
    .C(net209),
    .D(net159),
    .X(_1414_));
 sky130_fd_sc_hd__or2_1 _2319_ (.A(net76),
    .B(_1414_),
    .X(_1415_));
 sky130_fd_sc_hd__nor2_1 _2320_ (.A(net107),
    .B(_1389_),
    .Y(_1416_));
 sky130_fd_sc_hd__and4_4 _2321_ (.A(net255),
    .B(net222),
    .C(net180),
    .D(net156),
    .X(_1417_));
 sky130_fd_sc_hd__o2111a_4 _2322_ (.A1(net184),
    .A2(net181),
    .B1(net163),
    .C1(net227),
    .D1(net263),
    .X(_1418_));
 sky130_fd_sc_hd__or3_2 _2323_ (.A(net76),
    .B(_1414_),
    .C(_1418_),
    .X(_1419_));
 sky130_fd_sc_hd__nor2_8 _2324_ (.A(net96),
    .B(net167),
    .Y(_1420_));
 sky130_fd_sc_hd__nor2_8 _2325_ (.A(net95),
    .B(net132),
    .Y(_1421_));
 sky130_fd_sc_hd__a21oi_4 _2326_ (.A1(net167),
    .A2(net131),
    .B1(net96),
    .Y(_1422_));
 sky130_fd_sc_hd__and4_4 _2327_ (.A(net250),
    .B(net236),
    .C(net183),
    .D(net162),
    .X(_1423_));
 sky130_fd_sc_hd__and4_4 _2328_ (.A(net250),
    .B(net236),
    .C(net162),
    .D(net155),
    .X(_1424_));
 sky130_fd_sc_hd__or2_4 _2329_ (.A(_1423_),
    .B(_1424_),
    .X(_1425_));
 sky130_fd_sc_hd__or4_1 _2330_ (.A(_1412_),
    .B(_1419_),
    .C(_1422_),
    .D(_1425_),
    .X(_1426_));
 sky130_fd_sc_hd__and4_4 _2331_ (.A(net276),
    .B(_0594_),
    .C(_0616_),
    .D(_1401_),
    .X(_1427_));
 sky130_fd_sc_hd__nor2_2 _2332_ (.A(net186),
    .B(_1318_),
    .Y(_1428_));
 sky130_fd_sc_hd__o2111a_4 _2333_ (.A1(net187),
    .A2(net169),
    .B1(net260),
    .C1(net224),
    .D1(net216),
    .X(_1429_));
 sky130_fd_sc_hd__or2_4 _2334_ (.A(_1346_),
    .B(_1429_),
    .X(_1430_));
 sky130_fd_sc_hd__and4_4 _2335_ (.A(net247),
    .B(net231),
    .C(net212),
    .D(net138),
    .X(_1431_));
 sky130_fd_sc_hd__and4_4 _2336_ (.A(net247),
    .B(net230),
    .C(net212),
    .D(net133),
    .X(_1432_));
 sky130_fd_sc_hd__or2_4 _2337_ (.A(_1431_),
    .B(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__and4_4 _2338_ (.A(net249),
    .B(net235),
    .C(net216),
    .D(net169),
    .X(_1434_));
 sky130_fd_sc_hd__and4_4 _2339_ (.A(net245),
    .B(net232),
    .C(net213),
    .D(net179),
    .X(_1435_));
 sky130_fd_sc_hd__or2_1 _2340_ (.A(_1434_),
    .B(_1435_),
    .X(_1436_));
 sky130_fd_sc_hd__or3_4 _2341_ (.A(_1430_),
    .B(_1433_),
    .C(_1436_),
    .X(_1437_));
 sky130_fd_sc_hd__and4_4 _2342_ (.A(net258),
    .B(net223),
    .C(net196),
    .D(net158),
    .X(_1438_));
 sky130_fd_sc_hd__or2_2 _2343_ (.A(_1391_),
    .B(net75),
    .X(_1439_));
 sky130_fd_sc_hd__and4_4 _2344_ (.A(net254),
    .B(net236),
    .C(net162),
    .D(net145),
    .X(_1440_));
 sky130_fd_sc_hd__and4_4 _2345_ (.A(net242),
    .B(net248),
    .C(net233),
    .D(net158),
    .X(_1441_));
 sky130_fd_sc_hd__nor2_8 _2346_ (.A(net190),
    .B(net77),
    .Y(_1442_));
 sky130_fd_sc_hd__nor2_8 _2347_ (.A(net200),
    .B(net77),
    .Y(_1443_));
 sky130_fd_sc_hd__a21oi_2 _2348_ (.A1(net200),
    .A2(net190),
    .B1(net77),
    .Y(_1444_));
 sky130_fd_sc_hd__nor2_8 _2349_ (.A(net122),
    .B(net100),
    .Y(_1445_));
 sky130_fd_sc_hd__nor2_8 _2350_ (.A(net171),
    .B(net95),
    .Y(_1446_));
 sky130_fd_sc_hd__a22o_4 _2351_ (.A1(net125),
    .A2(net181),
    .B1(net173),
    .B2(net98),
    .X(_1447_));
 sky130_fd_sc_hd__or3_1 _2352_ (.A(_1440_),
    .B(net74),
    .C(_1447_),
    .X(_1448_));
 sky130_fd_sc_hd__or4_1 _2353_ (.A(_1437_),
    .B(_1439_),
    .C(_1444_),
    .D(_1448_),
    .X(_1449_));
 sky130_fd_sc_hd__a22o_1 _2354_ (.A1(_1403_),
    .A2(_1426_),
    .B1(_1427_),
    .B2(_1449_),
    .X(_1450_));
 sky130_fd_sc_hd__and3_4 _2355_ (.A(_0594_),
    .B(_1386_),
    .C(_1401_),
    .X(_1451_));
 sky130_fd_sc_hd__nor2_4 _2356_ (.A(net93),
    .B(net87),
    .Y(_1452_));
 sky130_fd_sc_hd__a21oi_4 _2357_ (.A1(net113),
    .A2(net91),
    .B1(net86),
    .Y(_1453_));
 sky130_fd_sc_hd__nor2_8 _2358_ (.A(net95),
    .B(net137),
    .Y(_1454_));
 sky130_fd_sc_hd__a21oi_4 _2359_ (.A1(net136),
    .A2(net130),
    .B1(net96),
    .Y(_1455_));
 sky130_fd_sc_hd__or4_1 _2360_ (.A(_1290_),
    .B(_1293_),
    .C(_1453_),
    .D(_1455_),
    .X(_1456_));
 sky130_fd_sc_hd__nor2_4 _2361_ (.A(net241),
    .B(net102),
    .Y(_1457_));
 sky130_fd_sc_hd__a21oi_4 _2362_ (.A1(_0770_),
    .A2(net185),
    .B1(net103),
    .Y(_1458_));
 sky130_fd_sc_hd__and4_4 _2363_ (.A(net246),
    .B(net223),
    .C(net169),
    .D(net157),
    .X(_1459_));
 sky130_fd_sc_hd__and4_4 _2364_ (.A(net250),
    .B(net226),
    .C(net203),
    .D(net162),
    .X(_1460_));
 sky130_fd_sc_hd__or2_4 _2365_ (.A(_1459_),
    .B(_1460_),
    .X(_1461_));
 sky130_fd_sc_hd__or3_1 _2366_ (.A(_1456_),
    .B(_1458_),
    .C(_1461_),
    .X(_1462_));
 sky130_fd_sc_hd__nor2_4 _2367_ (.A(_1278_),
    .B(_1404_),
    .Y(_1463_));
 sky130_fd_sc_hd__nor2_4 _2368_ (.A(net201),
    .B(_1404_),
    .Y(_1464_));
 sky130_fd_sc_hd__a21oi_4 _2369_ (.A1(net200),
    .A2(net167),
    .B1(_1404_),
    .Y(_1465_));
 sky130_fd_sc_hd__nor2_1 _2370_ (.A(net137),
    .B(net80),
    .Y(_1466_));
 sky130_fd_sc_hd__nor2_8 _2371_ (.A(net176),
    .B(net80),
    .Y(_1467_));
 sky130_fd_sc_hd__a21oi_4 _2372_ (.A1(net174),
    .A2(net136),
    .B1(net77),
    .Y(_1468_));
 sky130_fd_sc_hd__nor2_8 _2373_ (.A(net170),
    .B(net77),
    .Y(_1469_));
 sky130_fd_sc_hd__nor2_4 _2374_ (.A(net208),
    .B(net80),
    .Y(_1470_));
 sky130_fd_sc_hd__a21oi_4 _2375_ (.A1(net207),
    .A2(net170),
    .B1(net77),
    .Y(_1471_));
 sky130_fd_sc_hd__a21oi_2 _2376_ (.A1(net148),
    .A2(net142),
    .B1(_1404_),
    .Y(_1472_));
 sky130_fd_sc_hd__or4_1 _2377_ (.A(_1465_),
    .B(_1468_),
    .C(_1471_),
    .D(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__or2_1 _2378_ (.A(_1444_),
    .B(_1473_),
    .X(_1474_));
 sky130_fd_sc_hd__a22o_1 _2379_ (.A1(net40),
    .A2(_1462_),
    .B1(_1474_),
    .B2(net46),
    .X(_1475_));
 sky130_fd_sc_hd__or4_1 _2380_ (.A(_1335_),
    .B(_1400_),
    .C(_1450_),
    .D(_1475_),
    .X(_1476_));
 sky130_fd_sc_hd__or3_4 _2381_ (.A(net253),
    .B(net229),
    .C(_1287_),
    .X(_1477_));
 sky130_fd_sc_hd__and4_4 _2382_ (.A(net261),
    .B(net236),
    .C(net162),
    .D(net133),
    .X(_1478_));
 sky130_fd_sc_hd__nor2_8 _2383_ (.A(net96),
    .B(net92),
    .Y(_1479_));
 sky130_fd_sc_hd__and4_4 _2384_ (.A(net247),
    .B(net222),
    .C(net157),
    .D(net133),
    .X(_1480_));
 sky130_fd_sc_hd__a2111o_1 _2385_ (.A1(net98),
    .A2(net155),
    .B1(_1460_),
    .C1(_1478_),
    .D1(_1480_),
    .X(_1481_));
 sky130_fd_sc_hd__o41a_1 _2386_ (.A1(_1414_),
    .A2(_1439_),
    .A3(net74),
    .A4(_1481_),
    .B1(net55),
    .X(_1482_));
 sky130_fd_sc_hd__nor2_4 _2387_ (.A(_1336_),
    .B(_1402_),
    .Y(_1483_));
 sky130_fd_sc_hd__and4_4 _2388_ (.A(net249),
    .B(net224),
    .C(net217),
    .D(net169),
    .X(_1484_));
 sky130_fd_sc_hd__or2_4 _2389_ (.A(_1331_),
    .B(_1484_),
    .X(_1485_));
 sky130_fd_sc_hd__nor2_4 _2390_ (.A(net192),
    .B(net87),
    .Y(_1486_));
 sky130_fd_sc_hd__a21oi_4 _2391_ (.A1(net190),
    .A2(_1236_),
    .B1(net85),
    .Y(_1487_));
 sky130_fd_sc_hd__nor2_8 _2392_ (.A(net127),
    .B(net170),
    .Y(_1488_));
 sky130_fd_sc_hd__nor2_8 _2393_ (.A(net127),
    .B(net207),
    .Y(_1489_));
 sky130_fd_sc_hd__a21oi_4 _2394_ (.A1(net207),
    .A2(net170),
    .B1(net126),
    .Y(_1490_));
 sky130_fd_sc_hd__a21oi_4 _2395_ (.A1(net106),
    .A2(net91),
    .B1(net97),
    .Y(_1491_));
 sky130_fd_sc_hd__o41a_1 _2396_ (.A1(_1485_),
    .A2(_1487_),
    .A3(_1490_),
    .A4(_1491_),
    .B1(net36),
    .X(_1492_));
 sky130_fd_sc_hd__nor3_4 _2397_ (.A(_0605_),
    .B(_1313_),
    .C(_1402_),
    .Y(_1493_));
 sky130_fd_sc_hd__and4_4 _2398_ (.A(net245),
    .B(net221),
    .C(net213),
    .D(net193),
    .X(_1494_));
 sky130_fd_sc_hd__and4_4 _2399_ (.A(net245),
    .B(net221),
    .C(net214),
    .D(net187),
    .X(_1495_));
 sky130_fd_sc_hd__or2_1 _2400_ (.A(_1494_),
    .B(_1495_),
    .X(_1496_));
 sky130_fd_sc_hd__o21a_1 _2401_ (.A1(_1268_),
    .A2(_1496_),
    .B1(_1493_),
    .X(_1497_));
 sky130_fd_sc_hd__nor2_4 _2402_ (.A(net116),
    .B(net192),
    .Y(_1498_));
 sky130_fd_sc_hd__a21o_2 _2403_ (.A1(_1089_),
    .A2(net195),
    .B1(_1478_),
    .X(_1499_));
 sky130_fd_sc_hd__nor2_8 _2404_ (.A(net207),
    .B(net85),
    .Y(_1500_));
 sky130_fd_sc_hd__nor2_4 _2405_ (.A(net87),
    .B(net132),
    .Y(_1501_));
 sky130_fd_sc_hd__a21oi_4 _2406_ (.A1(net207),
    .A2(net130),
    .B1(net86),
    .Y(_1502_));
 sky130_fd_sc_hd__o31a_1 _2407_ (.A1(_1296_),
    .A2(_1499_),
    .A3(_1502_),
    .B1(net59),
    .X(_1503_));
 sky130_fd_sc_hd__or4_4 _2408_ (.A(_1482_),
    .B(_1492_),
    .C(_1497_),
    .D(_1503_),
    .X(_1504_));
 sky130_fd_sc_hd__nor3b_4 _2409_ (.A(_0605_),
    .B(_1313_),
    .C_N(_1337_),
    .Y(_1505_));
 sky130_fd_sc_hd__and4_4 _2410_ (.A(net260),
    .B(net223),
    .C(net209),
    .D(net161),
    .X(_1506_));
 sky130_fd_sc_hd__and4_4 _2411_ (.A(net255),
    .B(net222),
    .C(net172),
    .D(net156),
    .X(_1507_));
 sky130_fd_sc_hd__or2_4 _2412_ (.A(_1506_),
    .B(net73),
    .X(_1508_));
 sky130_fd_sc_hd__nor2_8 _2413_ (.A(net111),
    .B(_1307_),
    .Y(_1509_));
 sky130_fd_sc_hd__nor2_1 _2414_ (.A(net111),
    .B(net150),
    .Y(_1510_));
 sky130_fd_sc_hd__a21oi_4 _2415_ (.A1(net149),
    .A2(net143),
    .B1(net110),
    .Y(_1511_));
 sky130_fd_sc_hd__and4_4 _2416_ (.A(net258),
    .B(net233),
    .C(net196),
    .D(net158),
    .X(_1512_));
 sky130_fd_sc_hd__and4_4 _2417_ (.A(net255),
    .B(net230),
    .C(net156),
    .D(net154),
    .X(_1513_));
 sky130_fd_sc_hd__or2_2 _2418_ (.A(net72),
    .B(net71),
    .X(_1514_));
 sky130_fd_sc_hd__o41a_1 _2419_ (.A1(_1378_),
    .A2(_1508_),
    .A3(_1511_),
    .A4(_1514_),
    .B1(net34),
    .X(_1515_));
 sky130_fd_sc_hd__a21o_1 _2420_ (.A1(net169),
    .A2(net83),
    .B1(_1435_),
    .X(_1516_));
 sky130_fd_sc_hd__and4_4 _2421_ (.A(net245),
    .B(net232),
    .C(net213),
    .D(net144),
    .X(_1517_));
 sky130_fd_sc_hd__and4_4 _2422_ (.A(net248),
    .B(net233),
    .C(net218),
    .D(net193),
    .X(_1518_));
 sky130_fd_sc_hd__or2_4 _2423_ (.A(_1517_),
    .B(_1518_),
    .X(_1519_));
 sky130_fd_sc_hd__o31a_1 _2424_ (.A1(_1331_),
    .A2(_1516_),
    .A3(_1519_),
    .B1(net54),
    .X(_1520_));
 sky130_fd_sc_hd__nor2_8 _2425_ (.A(_1262_),
    .B(_1336_),
    .Y(_1521_));
 sky130_fd_sc_hd__o21a_1 _2426_ (.A1(_1362_),
    .A2(_1506_),
    .B1(net31),
    .X(_1522_));
 sky130_fd_sc_hd__a2111o_1 _2427_ (.A1(net49),
    .A2(_1442_),
    .B1(_1515_),
    .C1(_1520_),
    .D1(_1522_),
    .X(_1523_));
 sky130_fd_sc_hd__or3_4 _2428_ (.A(net272),
    .B(net267),
    .C(_1389_),
    .X(_1524_));
 sky130_fd_sc_hd__and4_4 _2429_ (.A(net248),
    .B(net234),
    .C(net161),
    .D(net133),
    .X(_1525_));
 sky130_fd_sc_hd__and4_4 _2430_ (.A(net248),
    .B(net234),
    .C(net160),
    .D(net139),
    .X(_1526_));
 sky130_fd_sc_hd__o2111a_2 _2431_ (.A1(net141),
    .A2(net134),
    .B1(net251),
    .C1(net238),
    .D1(net163),
    .X(_1527_));
 sky130_fd_sc_hd__and4_4 _2432_ (.A(net246),
    .B(net235),
    .C(net179),
    .D(net157),
    .X(_1528_));
 sky130_fd_sc_hd__and4_4 _2433_ (.A(net248),
    .B(net233),
    .C(net209),
    .D(net159),
    .X(_1529_));
 sky130_fd_sc_hd__or2_1 _2434_ (.A(_1528_),
    .B(_1529_),
    .X(_1530_));
 sky130_fd_sc_hd__or3_4 _2435_ (.A(_1527_),
    .B(_1528_),
    .C(_1529_),
    .X(_1531_));
 sky130_fd_sc_hd__nand2b_4 _2436_ (.A_N(_1531_),
    .B(_1524_),
    .Y(_1532_));
 sky130_fd_sc_hd__nor2_4 _2437_ (.A(net128),
    .B(net150),
    .Y(_1533_));
 sky130_fd_sc_hd__nor2_1 _2438_ (.A(net118),
    .B(net101),
    .Y(_1534_));
 sky130_fd_sc_hd__nor2_2 _2439_ (.A(net121),
    .B(net201),
    .Y(_1535_));
 sky130_fd_sc_hd__or4_1 _2440_ (.A(net72),
    .B(_1533_),
    .C(net27),
    .D(_1535_),
    .X(_1536_));
 sky130_fd_sc_hd__and4_4 _2441_ (.A(net258),
    .B(net233),
    .C(net159),
    .D(net151),
    .X(_1537_));
 sky130_fd_sc_hd__a21o_4 _2442_ (.A1(net119),
    .A2(net182),
    .B1(_1537_),
    .X(_1538_));
 sky130_fd_sc_hd__nor2_1 _2443_ (.A(net208),
    .B(net95),
    .Y(_1539_));
 sky130_fd_sc_hd__a21oi_2 _2444_ (.A1(net208),
    .A2(net171),
    .B1(net97),
    .Y(_1540_));
 sky130_fd_sc_hd__o2111a_2 _2445_ (.A1(net183),
    .A2(_1294_),
    .B1(net163),
    .C1(net263),
    .D1(net227),
    .X(_1541_));
 sky130_fd_sc_hd__or3_1 _2446_ (.A(_1538_),
    .B(_1540_),
    .C(_1541_),
    .X(_1542_));
 sky130_fd_sc_hd__o31a_1 _2447_ (.A1(_1532_),
    .A2(_1536_),
    .A3(_1542_),
    .B1(net49),
    .X(_1543_));
 sky130_fd_sc_hd__and4_4 _2448_ (.A(net249),
    .B(net224),
    .C(net216),
    .D(net154),
    .X(_1544_));
 sky130_fd_sc_hd__nor2_8 _2449_ (.A(net128),
    .B(net136),
    .Y(_1545_));
 sky130_fd_sc_hd__a221o_1 _2450_ (.A1(net129),
    .A2(net209),
    .B1(net119),
    .B2(net139),
    .C1(_1537_),
    .X(_1546_));
 sky130_fd_sc_hd__o31a_1 _2451_ (.A1(_1544_),
    .A2(_1545_),
    .A3(_1546_),
    .B1(net63),
    .X(_1547_));
 sky130_fd_sc_hd__and4_4 _2452_ (.A(net247),
    .B(net231),
    .C(net212),
    .D(net202),
    .X(_1548_));
 sky130_fd_sc_hd__o2111a_4 _2453_ (.A1(net204),
    .A2(net194),
    .B1(net251),
    .C1(net238),
    .D1(net220),
    .X(_1549_));
 sky130_fd_sc_hd__nor2_8 _2454_ (.A(net174),
    .B(net96),
    .Y(_1550_));
 sky130_fd_sc_hd__or4_1 _2455_ (.A(_1344_),
    .B(_1454_),
    .C(_1549_),
    .D(_1550_),
    .X(_1551_));
 sky130_fd_sc_hd__nor2_8 _2456_ (.A(net165),
    .B(net80),
    .Y(_1552_));
 sky130_fd_sc_hd__a221o_1 _2457_ (.A1(net43),
    .A2(_1551_),
    .B1(_1552_),
    .B2(net52),
    .C1(_1547_),
    .X(_1553_));
 sky130_fd_sc_hd__or4_1 _2458_ (.A(_1504_),
    .B(_1523_),
    .C(_1543_),
    .D(_1553_),
    .X(_1554_));
 sky130_fd_sc_hd__nor2_8 _2459_ (.A(net176),
    .B(_1289_),
    .Y(_1555_));
 sky130_fd_sc_hd__nor2_2 _2460_ (.A(net186),
    .B(net80),
    .Y(_1556_));
 sky130_fd_sc_hd__and4_4 _2461_ (.A(net250),
    .B(net236),
    .C(net180),
    .D(net162),
    .X(_1557_));
 sky130_fd_sc_hd__or4_1 _2462_ (.A(_1296_),
    .B(_1555_),
    .C(_1556_),
    .D(_1557_),
    .X(_1558_));
 sky130_fd_sc_hd__and4_4 _2463_ (.A(net255),
    .B(net230),
    .C(net215),
    .D(net193),
    .X(_1559_));
 sky130_fd_sc_hd__or2_4 _2464_ (.A(_1434_),
    .B(_1559_),
    .X(_1560_));
 sky130_fd_sc_hd__nor2_2 _2465_ (.A(net93),
    .B(net80),
    .Y(_1561_));
 sky130_fd_sc_hd__or4_1 _2466_ (.A(_1283_),
    .B(_1347_),
    .C(_1388_),
    .D(_1561_),
    .X(_1562_));
 sky130_fd_sc_hd__o31a_1 _2467_ (.A1(_1558_),
    .A2(_1560_),
    .A3(_1562_),
    .B1(_1403_),
    .X(_1563_));
 sky130_fd_sc_hd__nor2_8 _2468_ (.A(_1023_),
    .B(net114),
    .Y(_1564_));
 sky130_fd_sc_hd__and4_4 _2469_ (.A(net245),
    .B(net232),
    .C(net213),
    .D(net154),
    .X(_1565_));
 sky130_fd_sc_hd__a211o_1 _2470_ (.A1(net205),
    .A2(net89),
    .B1(_1342_),
    .C1(_1565_),
    .X(_1566_));
 sky130_fd_sc_hd__o211ai_2 _2471_ (.A1(_1564_),
    .A2(_1566_),
    .B1(_0594_),
    .C1(_1386_),
    .Y(_1567_));
 sky130_fd_sc_hd__and4_4 _2472_ (.A(net261),
    .B(net226),
    .C(net188),
    .D(net164),
    .X(_1568_));
 sky130_fd_sc_hd__and4_4 _2473_ (.A(net247),
    .B(net230),
    .C(net187),
    .D(net156),
    .X(_1569_));
 sky130_fd_sc_hd__nor2_8 _2474_ (.A(net191),
    .B(_1404_),
    .Y(_1570_));
 sky130_fd_sc_hd__nor3_1 _2475_ (.A(_1568_),
    .B(_1569_),
    .C(_1570_),
    .Y(_1571_));
 sky130_fd_sc_hd__o21ai_2 _2476_ (.A1(_1336_),
    .A2(_1571_),
    .B1(_1567_),
    .Y(_1572_));
 sky130_fd_sc_hd__and3_2 _2477_ (.A(_0572_),
    .B(_0594_),
    .C(_1386_),
    .X(_1573_));
 sky130_fd_sc_hd__and4_4 _2478_ (.A(net246),
    .B(net232),
    .C(net217),
    .D(net182),
    .X(_1574_));
 sky130_fd_sc_hd__and4_4 _2479_ (.A(net249),
    .B(net224),
    .C(net216),
    .D(net209),
    .X(_1575_));
 sky130_fd_sc_hd__o21a_1 _2480_ (.A1(net244),
    .A2(net146),
    .B1(_1340_),
    .X(_1576_));
 sky130_fd_sc_hd__and4_4 _2481_ (.A(net245),
    .B(net221),
    .C(net213),
    .D(net172),
    .X(_1577_));
 sky130_fd_sc_hd__and4_4 _2482_ (.A(net245),
    .B(net232),
    .C(net213),
    .D(net180),
    .X(_1578_));
 sky130_fd_sc_hd__or2_4 _2483_ (.A(_1574_),
    .B(_1578_),
    .X(_1579_));
 sky130_fd_sc_hd__or4_1 _2484_ (.A(_1575_),
    .B(_1576_),
    .C(_1577_),
    .D(_1579_),
    .X(_1580_));
 sky130_fd_sc_hd__nor2_1 _2485_ (.A(net201),
    .B(net95),
    .Y(_1581_));
 sky130_fd_sc_hd__a21oi_2 _2486_ (.A1(net199),
    .A2(net166),
    .B1(net97),
    .Y(_1582_));
 sky130_fd_sc_hd__nor2_8 _2487_ (.A(net190),
    .B(net96),
    .Y(_1583_));
 sky130_fd_sc_hd__a21oi_4 _2488_ (.A1(net192),
    .A2(net186),
    .B1(net97),
    .Y(_1584_));
 sky130_fd_sc_hd__or2_1 _2489_ (.A(_1582_),
    .B(_1584_),
    .X(_1585_));
 sky130_fd_sc_hd__a211o_1 _2490_ (.A1(net197),
    .A2(net84),
    .B1(_1321_),
    .C1(_1339_),
    .X(_1586_));
 sky130_fd_sc_hd__o31a_1 _2491_ (.A1(_1580_),
    .A2(_1585_),
    .A3(_1586_),
    .B1(net26),
    .X(_1587_));
 sky130_fd_sc_hd__nor3_4 _2492_ (.A(_0583_),
    .B(_0605_),
    .C(_1313_),
    .Y(_1588_));
 sky130_fd_sc_hd__nor2_8 _2493_ (.A(net127),
    .B(net200),
    .Y(_1589_));
 sky130_fd_sc_hd__nor2_8 _2494_ (.A(net127),
    .B(net191),
    .Y(_1590_));
 sky130_fd_sc_hd__nor2_8 _2495_ (.A(net126),
    .B(net142),
    .Y(_1591_));
 sky130_fd_sc_hd__o41a_4 _2496_ (.A1(net205),
    .A2(net194),
    .A3(net152),
    .A4(net146),
    .B1(net129),
    .X(_1592_));
 sky130_fd_sc_hd__nor2_4 _2497_ (.A(_0968_),
    .B(net142),
    .Y(_1593_));
 sky130_fd_sc_hd__or4b_1 _2498_ (.A(net262),
    .B(net142),
    .C(net237),
    .D_N(_0946_),
    .X(_1594_));
 sky130_fd_sc_hd__o2111a_4 _2499_ (.A1(net242),
    .A2(net144),
    .B1(net220),
    .C1(net227),
    .D1(net251),
    .X(_1595_));
 sky130_fd_sc_hd__nor2_8 _2500_ (.A(net126),
    .B(net165),
    .Y(_1596_));
 sky130_fd_sc_hd__nor2_4 _2501_ (.A(net126),
    .B(net132),
    .Y(_1597_));
 sky130_fd_sc_hd__a21oi_4 _2502_ (.A1(net165),
    .A2(net132),
    .B1(net126),
    .Y(_1598_));
 sky130_fd_sc_hd__and4_4 _2503_ (.A(net254),
    .B(net226),
    .C(net219),
    .D(net180),
    .X(_1599_));
 sky130_fd_sc_hd__nor2_2 _2504_ (.A(_0968_),
    .B(net107),
    .Y(_1600_));
 sky130_fd_sc_hd__a21oi_4 _2505_ (.A1(net107),
    .A2(net101),
    .B1(_0968_),
    .Y(_1601_));
 sky130_fd_sc_hd__or4_1 _2506_ (.A(_1268_),
    .B(_1595_),
    .C(_1598_),
    .D(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__o21a_2 _2507_ (.A1(_1592_),
    .A2(_1602_),
    .B1(net21),
    .X(_1603_));
 sky130_fd_sc_hd__a2111o_2 _2508_ (.A1(_0572_),
    .A2(_1572_),
    .B1(_1587_),
    .C1(_1603_),
    .D1(_1563_),
    .X(_1604_));
 sky130_fd_sc_hd__and3_4 _2509_ (.A(_0594_),
    .B(_1337_),
    .C(_1386_),
    .X(_1605_));
 sky130_fd_sc_hd__and4_4 _2510_ (.A(net261),
    .B(net239),
    .C(net219),
    .D(net188),
    .X(_1606_));
 sky130_fd_sc_hd__or2_4 _2511_ (.A(_1559_),
    .B(_1606_),
    .X(_1607_));
 sky130_fd_sc_hd__or4_2 _2512_ (.A(_1341_),
    .B(_1379_),
    .C(_1593_),
    .D(_1607_),
    .X(_1608_));
 sky130_fd_sc_hd__o21a_1 _2513_ (.A1(_1579_),
    .A2(_1608_),
    .B1(net34),
    .X(_1609_));
 sky130_fd_sc_hd__nor2_8 _2514_ (.A(net121),
    .B(net130),
    .Y(_1610_));
 sky130_fd_sc_hd__a2111o_1 _2515_ (.A1(net119),
    .A2(net144),
    .B1(_1363_),
    .C1(_1373_),
    .D1(_1545_),
    .X(_1611_));
 sky130_fd_sc_hd__o31a_1 _2516_ (.A1(net27),
    .A2(_1610_),
    .A3(_1611_),
    .B1(net29),
    .X(_1612_));
 sky130_fd_sc_hd__nor2_1 _2517_ (.A(net111),
    .B(net176),
    .Y(_1613_));
 sky130_fd_sc_hd__nor2_2 _2518_ (.A(net208),
    .B(net111),
    .Y(_1614_));
 sky130_fd_sc_hd__a21oi_4 _2519_ (.A1(net206),
    .A2(net175),
    .B1(net110),
    .Y(_1615_));
 sky130_fd_sc_hd__o31a_1 _2520_ (.A1(_1485_),
    .A2(_1598_),
    .A3(_1615_),
    .B1(net63),
    .X(_1616_));
 sky130_fd_sc_hd__a2111o_1 _2521_ (.A1(_1366_),
    .A2(net19),
    .B1(_1609_),
    .C1(_1612_),
    .D1(_1616_),
    .X(_1617_));
 sky130_fd_sc_hd__and4_4 _2522_ (.A(net256),
    .B(net231),
    .C(net213),
    .D(net172),
    .X(_1618_));
 sky130_fd_sc_hd__or2_1 _2523_ (.A(_1544_),
    .B(_1618_),
    .X(_1619_));
 sky130_fd_sc_hd__or3_1 _2524_ (.A(net76),
    .B(_1459_),
    .C(_1528_),
    .X(_1620_));
 sky130_fd_sc_hd__a22o_1 _2525_ (.A1(net21),
    .A2(_1619_),
    .B1(_1620_),
    .B2(net47),
    .X(_1621_));
 sky130_fd_sc_hd__nor2_2 _2526_ (.A(net102),
    .B(net132),
    .Y(_1622_));
 sky130_fd_sc_hd__a21oi_4 _2527_ (.A1(net167),
    .A2(net130),
    .B1(net103),
    .Y(_1623_));
 sky130_fd_sc_hd__nor2_8 _2528_ (.A(net240),
    .B(net109),
    .Y(_1624_));
 sky130_fd_sc_hd__a21oi_4 _2529_ (.A1(net240),
    .A2(net143),
    .B1(net110),
    .Y(_1625_));
 sky130_fd_sc_hd__nor2_4 _2530_ (.A(net111),
    .B(net107),
    .Y(_1626_));
 sky130_fd_sc_hd__nor2_8 _2531_ (.A(net111),
    .B(net101),
    .Y(_1627_));
 sky130_fd_sc_hd__a21oi_4 _2532_ (.A1(net106),
    .A2(net100),
    .B1(net109),
    .Y(_1628_));
 sky130_fd_sc_hd__nor2_8 _2533_ (.A(net110),
    .B(net92),
    .Y(_1629_));
 sky130_fd_sc_hd__a22o_1 _2534_ (.A1(net112),
    .A2(net155),
    .B1(net81),
    .B2(net173),
    .X(_1630_));
 sky130_fd_sc_hd__or3_4 _2535_ (.A(_1625_),
    .B(_1628_),
    .C(_1630_),
    .X(_1631_));
 sky130_fd_sc_hd__a221o_1 _2536_ (.A1(net36),
    .A2(_1623_),
    .B1(_1631_),
    .B2(net49),
    .C1(_1621_),
    .X(_1632_));
 sky130_fd_sc_hd__or4_2 _2537_ (.A(_1554_),
    .B(_1604_),
    .C(_1617_),
    .D(_1632_),
    .X(_1633_));
 sky130_fd_sc_hd__or2_4 _2538_ (.A(_1423_),
    .B(_1557_),
    .X(_1634_));
 sky130_fd_sc_hd__nor2_2 _2539_ (.A(net171),
    .B(net87),
    .Y(_1635_));
 sky130_fd_sc_hd__a21oi_2 _2540_ (.A1(net206),
    .A2(net170),
    .B1(net86),
    .Y(_1636_));
 sky130_fd_sc_hd__a21o_4 _2541_ (.A1(net173),
    .A2(net90),
    .B1(_1557_),
    .X(_1637_));
 sky130_fd_sc_hd__or2_1 _2542_ (.A(_1634_),
    .B(_1636_),
    .X(_1638_));
 sky130_fd_sc_hd__nor2_8 _2543_ (.A(net106),
    .B(net78),
    .Y(_1639_));
 sky130_fd_sc_hd__a21oi_2 _2544_ (.A1(net108),
    .A2(net92),
    .B1(net77),
    .Y(_1640_));
 sky130_fd_sc_hd__nor2_4 _2545_ (.A(net150),
    .B(net80),
    .Y(_1641_));
 sky130_fd_sc_hd__a21oi_4 _2546_ (.A1(net114),
    .A2(net148),
    .B1(net78),
    .Y(_1642_));
 sky130_fd_sc_hd__o41a_1 _2547_ (.A1(net198),
    .A2(net184),
    .A3(net155),
    .A4(net152),
    .B1(_1408_),
    .X(_1643_));
 sky130_fd_sc_hd__and4_4 _2548_ (.A(net243),
    .B(net251),
    .C(net227),
    .D(net163),
    .X(_1644_));
 sky130_fd_sc_hd__a21o_1 _2549_ (.A1(net240),
    .A2(net142),
    .B1(_1289_),
    .X(_1645_));
 sky130_fd_sc_hd__nor2_4 _2550_ (.A(net167),
    .B(net86),
    .Y(_1646_));
 sky130_fd_sc_hd__a21oi_2 _2551_ (.A1(net201),
    .A2(net165),
    .B1(net87),
    .Y(_1647_));
 sky130_fd_sc_hd__a211o_2 _2552_ (.A1(_1288_),
    .A2(net147),
    .B1(_1644_),
    .C1(_1647_),
    .X(_1648_));
 sky130_fd_sc_hd__nor2_8 _2553_ (.A(_1289_),
    .B(net137),
    .Y(_1649_));
 sky130_fd_sc_hd__a21oi_4 _2554_ (.A1(net174),
    .A2(net136),
    .B1(_1289_),
    .Y(_1650_));
 sky130_fd_sc_hd__a21oi_4 _2555_ (.A1(net199),
    .A2(net191),
    .B1(net96),
    .Y(_1651_));
 sky130_fd_sc_hd__nor2_2 _2556_ (.A(net186),
    .B(_1289_),
    .Y(_1652_));
 sky130_fd_sc_hd__o2111a_4 _2557_ (.A1(net194),
    .A2(net189),
    .B1(net163),
    .C1(net227),
    .D1(net252),
    .X(_1653_));
 sky130_fd_sc_hd__nor2_8 _2558_ (.A(net85),
    .B(net137),
    .Y(_1654_));
 sky130_fd_sc_hd__a21oi_1 _2559_ (.A1(net136),
    .A2(net130),
    .B1(net85),
    .Y(_1655_));
 sky130_fd_sc_hd__nor2_4 _2560_ (.A(net207),
    .B(net103),
    .Y(_1656_));
 sky130_fd_sc_hd__nor2_4 _2561_ (.A(net103),
    .B(net170),
    .Y(_1657_));
 sky130_fd_sc_hd__a21oi_2 _2562_ (.A1(net114),
    .A2(net148),
    .B1(net96),
    .Y(_1658_));
 sky130_fd_sc_hd__nand2_8 _2563_ (.A(net98),
    .B(net146),
    .Y(_1659_));
 sky130_fd_sc_hd__nor2_8 _2564_ (.A(net240),
    .B(net96),
    .Y(_1660_));
 sky130_fd_sc_hd__or3b_4 _2565_ (.A(_1660_),
    .B(_1658_),
    .C_N(_1659_),
    .X(_1661_));
 sky130_fd_sc_hd__or4_1 _2566_ (.A(_1642_),
    .B(_1656_),
    .C(net16),
    .D(_1661_),
    .X(_1662_));
 sky130_fd_sc_hd__or4_1 _2567_ (.A(_1422_),
    .B(_1488_),
    .C(_1578_),
    .D(_1640_),
    .X(_1663_));
 sky130_fd_sc_hd__o41a_4 _2568_ (.A1(net194),
    .A2(net189),
    .A3(net177),
    .A4(net140),
    .B1(_1288_),
    .X(_1664_));
 sky130_fd_sc_hd__or4_1 _2569_ (.A(_1447_),
    .B(_1651_),
    .C(_1655_),
    .D(_1664_),
    .X(_1665_));
 sky130_fd_sc_hd__or4_1 _2570_ (.A(_1638_),
    .B(_1648_),
    .C(_1663_),
    .D(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__o21a_1 _2571_ (.A1(_1662_),
    .A2(_1666_),
    .B1(net55),
    .X(_1667_));
 sky130_fd_sc_hd__a41o_1 _2572_ (.A1(net207),
    .A2(net176),
    .A3(net170),
    .A4(net136),
    .B1(net104),
    .X(_1668_));
 sky130_fd_sc_hd__nand2b_2 _2573_ (.A_N(_1642_),
    .B(_1668_),
    .Y(_1669_));
 sky130_fd_sc_hd__a21oi_2 _2574_ (.A1(net166),
    .A2(net130),
    .B1(net86),
    .Y(_1670_));
 sky130_fd_sc_hd__a21oi_4 _2575_ (.A1(net148),
    .A2(net142),
    .B1(net96),
    .Y(_1671_));
 sky130_fd_sc_hd__o2111a_4 _2576_ (.A1(net211),
    .A2(net177),
    .B1(net164),
    .C1(net227),
    .D1(net252),
    .X(_1672_));
 sky130_fd_sc_hd__o2111a_4 _2577_ (.A1(net140),
    .A2(net134),
    .B1(net251),
    .C1(net228),
    .D1(net163),
    .X(_1673_));
 sky130_fd_sc_hd__or2_4 _2578_ (.A(_1653_),
    .B(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__or4_1 _2579_ (.A(_1637_),
    .B(_1640_),
    .C(_1669_),
    .D(_1672_),
    .X(_1675_));
 sky130_fd_sc_hd__o41a_1 _2580_ (.A1(_1670_),
    .A2(_1671_),
    .A3(_1674_),
    .A4(_1675_),
    .B1(net26),
    .X(_1676_));
 sky130_fd_sc_hd__nor2_8 _2581_ (.A(net127),
    .B(net100),
    .Y(_1677_));
 sky130_fd_sc_hd__a21oi_4 _2582_ (.A1(net106),
    .A2(net100),
    .B1(net128),
    .Y(_1678_));
 sky130_fd_sc_hd__nor2_8 _2583_ (.A(net122),
    .B(net170),
    .Y(_1679_));
 sky130_fd_sc_hd__and4_4 _2584_ (.A(net260),
    .B(net235),
    .C(net217),
    .D(net139),
    .X(_1680_));
 sky130_fd_sc_hd__and4_4 _2585_ (.A(net255),
    .B(net230),
    .C(net215),
    .D(net133),
    .X(_1681_));
 sky130_fd_sc_hd__o2111a_4 _2586_ (.A1(net138),
    .A2(net133),
    .B1(net260),
    .C1(net235),
    .D1(net217),
    .X(_1682_));
 sky130_fd_sc_hd__and4_4 _2587_ (.A(net258),
    .B(net233),
    .C(net218),
    .D(net179),
    .X(_1683_));
 sky130_fd_sc_hd__o2111a_2 _2588_ (.A1(net177),
    .A2(net141),
    .B1(net263),
    .C1(net238),
    .D1(net220),
    .X(_1684_));
 sky130_fd_sc_hd__or3_1 _2589_ (.A(_1374_),
    .B(_1682_),
    .C(_1683_),
    .X(_1685_));
 sky130_fd_sc_hd__or4_1 _2590_ (.A(_1034_),
    .B(_1678_),
    .C(_1679_),
    .D(_1685_),
    .X(_1686_));
 sky130_fd_sc_hd__nor2_8 _2591_ (.A(net109),
    .B(net130),
    .Y(_1687_));
 sky130_fd_sc_hd__a21oi_4 _2592_ (.A1(net136),
    .A2(net131),
    .B1(net109),
    .Y(_1688_));
 sky130_fd_sc_hd__nor2_4 _2593_ (.A(net111),
    .B(net165),
    .Y(_1689_));
 sky130_fd_sc_hd__nor2_8 _2594_ (.A(net200),
    .B(net109),
    .Y(_1690_));
 sky130_fd_sc_hd__a21oi_4 _2595_ (.A1(net199),
    .A2(net166),
    .B1(net109),
    .Y(_1691_));
 sky130_fd_sc_hd__o41a_4 _2596_ (.A1(net204),
    .A2(net194),
    .A3(net189),
    .A4(net168),
    .B1(_1205_),
    .X(_1692_));
 sky130_fd_sc_hd__or2_2 _2597_ (.A(_1688_),
    .B(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__nor2_4 _2598_ (.A(net117),
    .B(net149),
    .Y(_1694_));
 sky130_fd_sc_hd__nor2_8 _2599_ (.A(net117),
    .B(net114),
    .Y(_1695_));
 sky130_fd_sc_hd__nor2_2 _2600_ (.A(net116),
    .B(net93),
    .Y(_1696_));
 sky130_fd_sc_hd__a21oi_4 _2601_ (.A1(net107),
    .A2(net93),
    .B1(net116),
    .Y(_1697_));
 sky130_fd_sc_hd__a41o_4 _2602_ (.A1(net113),
    .A2(net106),
    .A3(net91),
    .A4(net149),
    .B1(net117),
    .X(_1698_));
 sky130_fd_sc_hd__and4_4 _2603_ (.A(net258),
    .B(net233),
    .C(net158),
    .D(net144),
    .X(_1699_));
 sky130_fd_sc_hd__and4_4 _2604_ (.A(net242),
    .B(net259),
    .C(net234),
    .D(net160),
    .X(_1700_));
 sky130_fd_sc_hd__and4_4 _2605_ (.A(net261),
    .B(net236),
    .C(net187),
    .D(net162),
    .X(_1701_));
 sky130_fd_sc_hd__or2_1 _2606_ (.A(_1700_),
    .B(_1701_),
    .X(_1702_));
 sky130_fd_sc_hd__or4b_1 _2607_ (.A(_1537_),
    .B(_1699_),
    .C(_1702_),
    .D_N(_1698_),
    .X(_1703_));
 sky130_fd_sc_hd__or4_4 _2608_ (.A(_1511_),
    .B(_1686_),
    .C(_1693_),
    .D(_1703_),
    .X(_1704_));
 sky130_fd_sc_hd__or2_4 _2609_ (.A(_1599_),
    .B(_1618_),
    .X(_1705_));
 sky130_fd_sc_hd__or3_1 _2610_ (.A(_1677_),
    .B(_1679_),
    .C(_1705_),
    .X(_1706_));
 sky130_fd_sc_hd__and4_4 _2611_ (.A(net258),
    .B(net233),
    .C(net193),
    .D(net158),
    .X(_1707_));
 sky130_fd_sc_hd__a21o_4 _2612_ (.A1(net120),
    .A2(net145),
    .B1(_1707_),
    .X(_1708_));
 sky130_fd_sc_hd__and4_4 _2613_ (.A(net258),
    .B(net233),
    .C(net202),
    .D(net158),
    .X(_1709_));
 sky130_fd_sc_hd__a211o_1 _2614_ (.A1(net243),
    .A2(net120),
    .B1(_1708_),
    .C1(_1709_),
    .X(_1710_));
 sky130_fd_sc_hd__a21oi_4 _2615_ (.A1(net175),
    .A2(net166),
    .B1(net110),
    .Y(_1711_));
 sky130_fd_sc_hd__or2_1 _2616_ (.A(_1688_),
    .B(_1711_),
    .X(_1712_));
 sky130_fd_sc_hd__nor2_8 _2617_ (.A(net128),
    .B(net93),
    .Y(_1713_));
 sky130_fd_sc_hd__a21oi_4 _2618_ (.A1(net106),
    .A2(net91),
    .B1(net127),
    .Y(_1714_));
 sky130_fd_sc_hd__nor2_4 _2619_ (.A(net126),
    .B(net115),
    .Y(_1715_));
 sky130_fd_sc_hd__a21oi_2 _2620_ (.A1(net113),
    .A2(net149),
    .B1(net128),
    .Y(_1716_));
 sky130_fd_sc_hd__nor2_8 _2621_ (.A(net167),
    .B(_1477_),
    .Y(_1717_));
 sky130_fd_sc_hd__a31o_1 _2622_ (.A1(net166),
    .A2(net148),
    .A3(net131),
    .B1(_1477_),
    .X(_1718_));
 sky130_fd_sc_hd__or3b_1 _2623_ (.A(_1714_),
    .B(_1716_),
    .C_N(_1718_),
    .X(_1719_));
 sky130_fd_sc_hd__or4_1 _2624_ (.A(_1706_),
    .B(_1710_),
    .C(_1712_),
    .D(_1719_),
    .X(_1720_));
 sky130_fd_sc_hd__a22o_1 _2625_ (.A1(net31),
    .A2(_1704_),
    .B1(_1720_),
    .B2(net66),
    .X(_1721_));
 sky130_fd_sc_hd__and4_4 _2626_ (.A(net256),
    .B(net230),
    .C(net172),
    .D(net156),
    .X(_1722_));
 sky130_fd_sc_hd__or2_1 _2627_ (.A(_1290_),
    .B(_1722_),
    .X(_1723_));
 sky130_fd_sc_hd__a21oi_4 _2628_ (.A1(net108),
    .A2(net92),
    .B1(net85),
    .Y(_1724_));
 sky130_fd_sc_hd__or2_1 _2629_ (.A(_1723_),
    .B(_1724_),
    .X(_1725_));
 sky130_fd_sc_hd__a21oi_1 _2630_ (.A1(net114),
    .A2(net148),
    .B1(net85),
    .Y(_1726_));
 sky130_fd_sc_hd__a21o_4 _2631_ (.A1(net198),
    .A2(net88),
    .B1(_1457_),
    .X(_1727_));
 sky130_fd_sc_hd__or4_2 _2632_ (.A(_1458_),
    .B(_1723_),
    .C(_1724_),
    .D(_1726_),
    .X(_1728_));
 sky130_fd_sc_hd__a21oi_4 _2633_ (.A1(net199),
    .A2(net190),
    .B1(net118),
    .Y(_1729_));
 sky130_fd_sc_hd__nor2_8 _2634_ (.A(net116),
    .B(net186),
    .Y(_1730_));
 sky130_fd_sc_hd__a21oi_4 _2635_ (.A1(net240),
    .A2(net186),
    .B1(net117),
    .Y(_1731_));
 sky130_fd_sc_hd__or3_1 _2636_ (.A(_1258_),
    .B(_1729_),
    .C(_1731_),
    .X(_1732_));
 sky130_fd_sc_hd__nor2_2 _2637_ (.A(net110),
    .B(net171),
    .Y(_1733_));
 sky130_fd_sc_hd__a21oi_4 _2638_ (.A1(net207),
    .A2(net171),
    .B1(net109),
    .Y(_1734_));
 sky130_fd_sc_hd__or3_1 _2639_ (.A(_1478_),
    .B(_1717_),
    .C(_1734_),
    .X(_1735_));
 sky130_fd_sc_hd__nor2_4 _2640_ (.A(net116),
    .B(net132),
    .Y(_1736_));
 sky130_fd_sc_hd__a21o_1 _2641_ (.A1(net137),
    .A2(net131),
    .B1(net117),
    .X(_1737_));
 sky130_fd_sc_hd__a21o_1 _2642_ (.A1(net174),
    .A2(net137),
    .B1(net110),
    .X(_1738_));
 sky130_fd_sc_hd__a21oi_2 _2643_ (.A1(net174),
    .A2(net136),
    .B1(net110),
    .Y(_1739_));
 sky130_fd_sc_hd__nand2_1 _2644_ (.A(_1737_),
    .B(_1738_),
    .Y(_1740_));
 sky130_fd_sc_hd__o41a_1 _2645_ (.A1(_1728_),
    .A2(_1732_),
    .A3(_1735_),
    .A4(_1740_),
    .B1(net23),
    .X(_1741_));
 sky130_fd_sc_hd__or3_2 _2646_ (.A(_1494_),
    .B(_1495_),
    .C(_1595_),
    .X(_1742_));
 sky130_fd_sc_hd__o41a_4 _2647_ (.A1(net211),
    .A2(net177),
    .A3(net140),
    .A4(net134),
    .B1(net120),
    .X(_1743_));
 sky130_fd_sc_hd__nor2_4 _2648_ (.A(net132),
    .B(net80),
    .Y(_1744_));
 sky130_fd_sc_hd__a21oi_4 _2649_ (.A1(net167),
    .A2(net131),
    .B1(net77),
    .Y(_1745_));
 sky130_fd_sc_hd__nor2_4 _2650_ (.A(net102),
    .B(net150),
    .Y(_1746_));
 sky130_fd_sc_hd__nor2_4 _2651_ (.A(net103),
    .B(net142),
    .Y(_1747_));
 sky130_fd_sc_hd__a21oi_2 _2652_ (.A1(net150),
    .A2(net143),
    .B1(net102),
    .Y(_1748_));
 sky130_fd_sc_hd__or4_4 _2653_ (.A(_1742_),
    .B(_1743_),
    .C(_1745_),
    .D(_1748_),
    .X(_1749_));
 sky130_fd_sc_hd__a21oi_4 _2654_ (.A1(net149),
    .A2(net143),
    .B1(net121),
    .Y(_1750_));
 sky130_fd_sc_hd__or4_1 _2655_ (.A(_1589_),
    .B(_1596_),
    .C(_1601_),
    .D(_1750_),
    .X(_1751_));
 sky130_fd_sc_hd__o31a_1 _2656_ (.A1(_1728_),
    .A2(_1749_),
    .A3(_1751_),
    .B1(net19),
    .X(_1752_));
 sky130_fd_sc_hd__nor2_4 _2657_ (.A(net121),
    .B(net107),
    .Y(_1753_));
 sky130_fd_sc_hd__nor2_8 _2658_ (.A(net122),
    .B(net92),
    .Y(_1754_));
 sky130_fd_sc_hd__a21oi_4 _2659_ (.A1(net106),
    .A2(net91),
    .B1(net122),
    .Y(_1755_));
 sky130_fd_sc_hd__a21oi_1 _2660_ (.A1(net136),
    .A2(net130),
    .B1(net77),
    .Y(_1756_));
 sky130_fd_sc_hd__or2_2 _2661_ (.A(_1628_),
    .B(_1756_),
    .X(_1757_));
 sky130_fd_sc_hd__or3_1 _2662_ (.A(_1471_),
    .B(_1750_),
    .C(_1755_),
    .X(_1758_));
 sky130_fd_sc_hd__o31a_1 _2663_ (.A1(_1532_),
    .A2(_1757_),
    .A3(_1758_),
    .B1(net52),
    .X(_1759_));
 sky130_fd_sc_hd__a21oi_4 _2664_ (.A1(net113),
    .A2(net91),
    .B1(net97),
    .Y(_1760_));
 sky130_fd_sc_hd__or2_2 _2665_ (.A(_1651_),
    .B(_1760_),
    .X(_1761_));
 sky130_fd_sc_hd__and4_4 _2666_ (.A(net249),
    .B(net224),
    .C(net216),
    .D(net202),
    .X(_1762_));
 sky130_fd_sc_hd__and4_4 _2667_ (.A(net247),
    .B(net231),
    .C(net212),
    .D(net151),
    .X(_1763_));
 sky130_fd_sc_hd__a21oi_4 _2668_ (.A1(net136),
    .A2(net130),
    .B1(net103),
    .Y(_1764_));
 sky130_fd_sc_hd__a21oi_4 _2669_ (.A1(net206),
    .A2(net175),
    .B1(net104),
    .Y(_1765_));
 sky130_fd_sc_hd__o41a_4 _2670_ (.A1(net211),
    .A2(net178),
    .A3(net140),
    .A4(net134),
    .B1(net105),
    .X(_1766_));
 sky130_fd_sc_hd__and4_4 _2671_ (.A(net246),
    .B(net221),
    .C(net157),
    .D(net151),
    .X(_1767_));
 sky130_fd_sc_hd__o2111a_4 _2672_ (.A1(net152),
    .A2(net146),
    .B1(net251),
    .C1(net227),
    .D1(net163),
    .X(_1768_));
 sky130_fd_sc_hd__or3_4 _2673_ (.A(_1291_),
    .B(_1644_),
    .C(_1768_),
    .X(_1769_));
 sky130_fd_sc_hd__o41a_2 _2674_ (.A1(net204),
    .A2(net194),
    .A3(net189),
    .A4(net168),
    .B1(net89),
    .X(_1770_));
 sky130_fd_sc_hd__or2_1 _2675_ (.A(_1769_),
    .B(_1770_),
    .X(_1771_));
 sky130_fd_sc_hd__a21oi_2 _2676_ (.A1(net113),
    .A2(net91),
    .B1(net79),
    .Y(_1772_));
 sky130_fd_sc_hd__or3_2 _2677_ (.A(_1490_),
    .B(_1637_),
    .C(_1772_),
    .X(_1773_));
 sky130_fd_sc_hd__or4_2 _2678_ (.A(_1494_),
    .B(_1517_),
    .C(_1762_),
    .D(_1763_),
    .X(_1774_));
 sky130_fd_sc_hd__or2_1 _2679_ (.A(_1343_),
    .B(_1673_),
    .X(_1775_));
 sky130_fd_sc_hd__or4_1 _2680_ (.A(_1769_),
    .B(_1770_),
    .C(_1774_),
    .D(_1775_),
    .X(_1776_));
 sky130_fd_sc_hd__o41a_2 _2681_ (.A1(_1761_),
    .A2(_1766_),
    .A3(_1773_),
    .A4(_1776_),
    .B1(net59),
    .X(_1777_));
 sky130_fd_sc_hd__or4_1 _2682_ (.A(_1741_),
    .B(_1752_),
    .C(_1759_),
    .D(_1777_),
    .X(_1778_));
 sky130_fd_sc_hd__or4_4 _2683_ (.A(_1667_),
    .B(_1676_),
    .C(_1721_),
    .D(_1778_),
    .X(_1779_));
 sky130_fd_sc_hd__or3_4 _2684_ (.A(_1476_),
    .B(_1633_),
    .C(_1779_),
    .X(_1780_));
 sky130_fd_sc_hd__and4_4 _2685_ (.A(net259),
    .B(net234),
    .C(net160),
    .D(net138),
    .X(_1781_));
 sky130_fd_sc_hd__a21o_2 _2686_ (.A1(net123),
    .A2(net173),
    .B1(_1781_),
    .X(_1782_));
 sky130_fd_sc_hd__o31a_1 _2687_ (.A1(net27),
    .A2(_1768_),
    .A3(_1782_),
    .B1(net36),
    .X(_1783_));
 sky130_fd_sc_hd__a21o_1 _2688_ (.A1(net197),
    .A2(net88),
    .B1(_1257_),
    .X(_1784_));
 sky130_fd_sc_hd__and4_4 _2689_ (.A(net259),
    .B(net233),
    .C(net209),
    .D(net159),
    .X(_1785_));
 sky130_fd_sc_hd__o31a_1 _2690_ (.A1(_1495_),
    .A2(net71),
    .A3(net69),
    .B1(net21),
    .X(_1786_));
 sky130_fd_sc_hd__a21o_1 _2691_ (.A1(net88),
    .A2(net153),
    .B1(_1722_),
    .X(_1787_));
 sky130_fd_sc_hd__or3_4 _2692_ (.A(_1654_),
    .B(_1701_),
    .C(_1787_),
    .X(_1788_));
 sky130_fd_sc_hd__a21o_1 _2693_ (.A1(net209),
    .A2(net83),
    .B1(_1365_),
    .X(_1789_));
 sky130_fd_sc_hd__o41a_1 _2694_ (.A1(_1388_),
    .A2(_1518_),
    .A3(_1788_),
    .A4(_1789_),
    .B1(net39),
    .X(_1790_));
 sky130_fd_sc_hd__a2111o_1 _2695_ (.A1(net63),
    .A2(_1784_),
    .B1(_1786_),
    .C1(_1790_),
    .D1(_1783_),
    .X(_1791_));
 sky130_fd_sc_hd__and4_4 _2696_ (.A(net256),
    .B(net231),
    .C(net182),
    .D(net156),
    .X(_1792_));
 sky130_fd_sc_hd__or2_2 _2697_ (.A(_1525_),
    .B(_1792_),
    .X(_1793_));
 sky130_fd_sc_hd__nor2_8 _2698_ (.A(net206),
    .B(_1359_),
    .Y(_1794_));
 sky130_fd_sc_hd__and4_4 _2699_ (.A(net257),
    .B(net221),
    .C(net202),
    .D(net157),
    .X(_1795_));
 sky130_fd_sc_hd__or4_1 _2700_ (.A(_1707_),
    .B(_1793_),
    .C(_1794_),
    .D(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__a22o_1 _2701_ (.A1(net32),
    .A2(_1792_),
    .B1(_1796_),
    .B2(net29),
    .X(_1797_));
 sky130_fd_sc_hd__o21a_1 _2702_ (.A1(_1431_),
    .A2(_1574_),
    .B1(net54),
    .X(_1798_));
 sky130_fd_sc_hd__or2_1 _2703_ (.A(_1366_),
    .B(_1548_),
    .X(_1799_));
 sky130_fd_sc_hd__a211o_1 _2704_ (.A1(net44),
    .A2(_1799_),
    .B1(_1798_),
    .C1(_1797_),
    .X(_1800_));
 sky130_fd_sc_hd__a21o_1 _2705_ (.A1(net64),
    .A2(_1627_),
    .B1(net44),
    .X(_1801_));
 sky130_fd_sc_hd__and4_4 _2706_ (.A(net242),
    .B(net261),
    .C(net226),
    .D(net162),
    .X(_1802_));
 sky130_fd_sc_hd__or2_4 _2707_ (.A(_1568_),
    .B(_1802_),
    .X(_1803_));
 sky130_fd_sc_hd__a21oi_4 _2708_ (.A1(net114),
    .A2(net148),
    .B1(net122),
    .Y(_1804_));
 sky130_fd_sc_hd__and4_4 _2709_ (.A(net263),
    .B(net227),
    .C(net194),
    .D(net164),
    .X(_1805_));
 sky130_fd_sc_hd__a21o_4 _2710_ (.A1(net125),
    .A2(net146),
    .B1(_1805_),
    .X(_1806_));
 sky130_fd_sc_hd__or3_1 _2711_ (.A(_1362_),
    .B(_1795_),
    .C(_1806_),
    .X(_1807_));
 sky130_fd_sc_hd__or4_1 _2712_ (.A(_1433_),
    .B(_1540_),
    .C(_1803_),
    .D(_1804_),
    .X(_1808_));
 sky130_fd_sc_hd__or4_2 _2713_ (.A(_1527_),
    .B(_1755_),
    .C(_1807_),
    .D(_1808_),
    .X(_1809_));
 sky130_fd_sc_hd__o21a_1 _2714_ (.A1(_1627_),
    .A2(_1809_),
    .B1(_1801_),
    .X(_1810_));
 sky130_fd_sc_hd__and4_4 _2715_ (.A(net258),
    .B(net223),
    .C(net158),
    .D(net151),
    .X(_1811_));
 sky130_fd_sc_hd__or2_4 _2716_ (.A(_1390_),
    .B(_1811_),
    .X(_1812_));
 sky130_fd_sc_hd__or4_2 _2717_ (.A(_1323_),
    .B(_1561_),
    .C(_1649_),
    .D(_1812_),
    .X(_1813_));
 sky130_fd_sc_hd__a21o_1 _2718_ (.A1(net129),
    .A2(net139),
    .B1(_1578_),
    .X(_1814_));
 sky130_fd_sc_hd__a2111o_1 _2719_ (.A1(net196),
    .A2(_1340_),
    .B1(_1420_),
    .C1(_1577_),
    .D1(_1814_),
    .X(_1815_));
 sky130_fd_sc_hd__o21a_1 _2720_ (.A1(_1470_),
    .A2(_1762_),
    .B1(net29),
    .X(_1816_));
 sky130_fd_sc_hd__a221o_1 _2721_ (.A1(net51),
    .A2(_1813_),
    .B1(_1815_),
    .B2(net57),
    .C1(_1816_),
    .X(_1817_));
 sky130_fd_sc_hd__or4_4 _2722_ (.A(_1791_),
    .B(_1800_),
    .C(_1810_),
    .D(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__or2_2 _2723_ (.A(_1424_),
    .B(net74),
    .X(_1819_));
 sky130_fd_sc_hd__or4_1 _2724_ (.A(_1410_),
    .B(_1454_),
    .C(_1556_),
    .D(_1570_),
    .X(_1820_));
 sky130_fd_sc_hd__o31a_1 _2725_ (.A1(_1416_),
    .A2(_1819_),
    .A3(_1820_),
    .B1(net46),
    .X(_1821_));
 sky130_fd_sc_hd__or4_1 _2726_ (.A(net28),
    .B(_1590_),
    .C(_1610_),
    .D(_1624_),
    .X(_1822_));
 sky130_fd_sc_hd__o21a_1 _2727_ (.A1(_0935_),
    .A2(_1822_),
    .B1(net33),
    .X(_1823_));
 sky130_fd_sc_hd__nor2_4 _2728_ (.A(net100),
    .B(net78),
    .Y(_1824_));
 sky130_fd_sc_hd__or4_1 _2729_ (.A(_1544_),
    .B(_1624_),
    .C(_1681_),
    .D(net14),
    .X(_1825_));
 sky130_fd_sc_hd__a211o_1 _2730_ (.A1(net19),
    .A2(_1825_),
    .B1(_1823_),
    .C1(_1821_),
    .X(_1826_));
 sky130_fd_sc_hd__o22ai_4 _2731_ (.A1(net208),
    .A2(net95),
    .B1(_1389_),
    .B2(net107),
    .Y(_1827_));
 sky130_fd_sc_hd__or3_1 _2732_ (.A(_1322_),
    .B(_1556_),
    .C(_1827_),
    .X(_1828_));
 sky130_fd_sc_hd__a22o_4 _2733_ (.A1(net154),
    .A2(net88),
    .B1(net144),
    .B2(net105),
    .X(_1829_));
 sky130_fd_sc_hd__a22o_1 _2734_ (.A1(net42),
    .A2(_1828_),
    .B1(_1829_),
    .B2(net24),
    .X(_1830_));
 sky130_fd_sc_hd__a221o_1 _2735_ (.A1(net58),
    .A2(_1349_),
    .B1(_1509_),
    .B2(net22),
    .C1(_1830_),
    .X(_1831_));
 sky130_fd_sc_hd__o31a_1 _2736_ (.A1(_1360_),
    .A2(_1682_),
    .A3(_1794_),
    .B1(net64),
    .X(_1832_));
 sky130_fd_sc_hd__o31a_1 _2737_ (.A1(_1349_),
    .A2(_1421_),
    .A3(_1763_),
    .B1(net24),
    .X(_1833_));
 sky130_fd_sc_hd__o21a_1 _2738_ (.A1(_1342_),
    .A2(_1420_),
    .B1(net35),
    .X(_1834_));
 sky130_fd_sc_hd__or2_2 _2739_ (.A(_0935_),
    .B(_1591_),
    .X(_1835_));
 sky130_fd_sc_hd__o41a_1 _2740_ (.A1(_1034_),
    .A2(_1499_),
    .A3(_1589_),
    .A4(_1835_),
    .B1(net63),
    .X(_1836_));
 sky130_fd_sc_hd__or4_1 _2741_ (.A(_1832_),
    .B(_1833_),
    .C(_1834_),
    .D(_1836_),
    .X(_1837_));
 sky130_fd_sc_hd__a21o_1 _2742_ (.A1(net198),
    .A2(net98),
    .B1(_1644_),
    .X(_1838_));
 sky130_fd_sc_hd__or2_1 _2743_ (.A(_1722_),
    .B(_1802_),
    .X(_1839_));
 sky130_fd_sc_hd__or4_2 _2744_ (.A(_1423_),
    .B(_1500_),
    .C(_1838_),
    .D(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__or4_1 _2745_ (.A(_1111_),
    .B(_1680_),
    .C(_1687_),
    .D(_1696_),
    .X(_1841_));
 sky130_fd_sc_hd__o41a_1 _2746_ (.A1(net82),
    .A2(_1375_),
    .A3(net15),
    .A4(_1841_),
    .B1(net37),
    .X(_1842_));
 sky130_fd_sc_hd__o21a_1 _2747_ (.A1(_1339_),
    .A2(_1598_),
    .B1(net35),
    .X(_1843_));
 sky130_fd_sc_hd__nor2_8 _2748_ (.A(net103),
    .B(net92),
    .Y(_1844_));
 sky130_fd_sc_hd__o31a_1 _2749_ (.A1(_1656_),
    .A2(_1747_),
    .A3(_1844_),
    .B1(net23),
    .X(_1845_));
 sky130_fd_sc_hd__a2111o_1 _2750_ (.A1(net24),
    .A2(_1840_),
    .B1(_1842_),
    .C1(_1843_),
    .D1(_1845_),
    .X(_1846_));
 sky130_fd_sc_hd__or4_1 _2751_ (.A(_1826_),
    .B(_1831_),
    .C(_1837_),
    .D(_1846_),
    .X(_1847_));
 sky130_fd_sc_hd__or4_1 _2752_ (.A(_1354_),
    .B(_1432_),
    .C(_1559_),
    .D(_1610_),
    .X(_1848_));
 sky130_fd_sc_hd__a21o_2 _2753_ (.A1(net209),
    .A2(net123),
    .B1(_1681_),
    .X(_1849_));
 sky130_fd_sc_hd__a22o_1 _2754_ (.A1(_0957_),
    .A2(net182),
    .B1(net83),
    .B2(net193),
    .X(_1850_));
 sky130_fd_sc_hd__and4_4 _2755_ (.A(net255),
    .B(net230),
    .C(net212),
    .D(net144),
    .X(_1851_));
 sky130_fd_sc_hd__or4_1 _2756_ (.A(_1366_),
    .B(_1849_),
    .C(_1850_),
    .D(_1851_),
    .X(_1852_));
 sky130_fd_sc_hd__o21a_1 _2757_ (.A1(_1848_),
    .A2(_1852_),
    .B1(net48),
    .X(_1853_));
 sky130_fd_sc_hd__o21a_1 _2758_ (.A1(net51),
    .A2(net39),
    .B1(_1794_),
    .X(_1854_));
 sky130_fd_sc_hd__a2111o_2 _2759_ (.A1(net124),
    .A2(net188),
    .B1(_1486_),
    .C1(_1596_),
    .D1(_1614_),
    .X(_1855_));
 sky130_fd_sc_hd__or4_1 _2760_ (.A(_1528_),
    .B(_1622_),
    .C(_1694_),
    .D(_1730_),
    .X(_1856_));
 sky130_fd_sc_hd__or4_1 _2761_ (.A(_1697_),
    .B(_1699_),
    .C(_1855_),
    .D(_1856_),
    .X(_1857_));
 sky130_fd_sc_hd__a211o_1 _2762_ (.A1(net64),
    .A2(_1857_),
    .B1(_1854_),
    .C1(_1853_),
    .X(_1858_));
 sky130_fd_sc_hd__or4_1 _2763_ (.A(net94),
    .B(_1709_),
    .C(_1715_),
    .D(_1781_),
    .X(_1859_));
 sky130_fd_sc_hd__a21o_2 _2764_ (.A1(net124),
    .A2(_1329_),
    .B1(_1506_),
    .X(_1860_));
 sky130_fd_sc_hd__o21a_1 _2765_ (.A1(_1859_),
    .A2(_1860_),
    .B1(net22),
    .X(_1861_));
 sky130_fd_sc_hd__or2_1 _2766_ (.A(net16),
    .B(_1747_),
    .X(_1862_));
 sky130_fd_sc_hd__o21a_1 _2767_ (.A1(_1689_),
    .A2(_1862_),
    .B1(net40),
    .X(_1863_));
 sky130_fd_sc_hd__o21a_1 _2768_ (.A1(_1254_),
    .A2(_1614_),
    .B1(net53),
    .X(_1864_));
 sky130_fd_sc_hd__o31a_1 _2769_ (.A1(_1341_),
    .A2(_1445_),
    .A3(_1581_),
    .B1(net50),
    .X(_1865_));
 sky130_fd_sc_hd__or4_1 _2770_ (.A(_1861_),
    .B(_1863_),
    .C(_1864_),
    .D(_1865_),
    .X(_1866_));
 sky130_fd_sc_hd__and4_4 _2771_ (.A(net258),
    .B(net223),
    .C(net158),
    .D(net138),
    .X(_1867_));
 sky130_fd_sc_hd__and4_4 _2772_ (.A(net247),
    .B(net230),
    .C(net172),
    .D(net156),
    .X(_1868_));
 sky130_fd_sc_hd__or4_1 _2773_ (.A(net73),
    .B(net71),
    .C(_1867_),
    .D(net68),
    .X(_1869_));
 sky130_fd_sc_hd__or2_4 _2774_ (.A(_1243_),
    .B(_1470_),
    .X(_1870_));
 sky130_fd_sc_hd__o41a_1 _2775_ (.A1(_1440_),
    .A2(_1443_),
    .A3(_1869_),
    .A4(_1870_),
    .B1(net48),
    .X(_1871_));
 sky130_fd_sc_hd__nor2_8 _2776_ (.A(net174),
    .B(net85),
    .Y(_1872_));
 sky130_fd_sc_hd__o31a_1 _2777_ (.A1(_1405_),
    .A2(_1459_),
    .A3(_1872_),
    .B1(net41),
    .X(_1873_));
 sky130_fd_sc_hd__or4_1 _2778_ (.A(_1279_),
    .B(_1283_),
    .C(_1614_),
    .D(_1652_),
    .X(_1874_));
 sky130_fd_sc_hd__o31a_1 _2779_ (.A1(_1459_),
    .A2(_1555_),
    .A3(_1874_),
    .B1(net58),
    .X(_1875_));
 sky130_fd_sc_hd__a22o_1 _2780_ (.A1(net129),
    .A2(net184),
    .B1(net153),
    .B2(net120),
    .X(_1876_));
 sky130_fd_sc_hd__o41a_1 _2781_ (.A1(_1347_),
    .A2(_1480_),
    .A3(_1548_),
    .A4(_1876_),
    .B1(net38),
    .X(_1877_));
 sky130_fd_sc_hd__or4_1 _2782_ (.A(_1871_),
    .B(_1873_),
    .C(_1875_),
    .D(_1877_),
    .X(_1878_));
 sky130_fd_sc_hd__or3_1 _2783_ (.A(_1858_),
    .B(_1866_),
    .C(_1878_),
    .X(_1879_));
 sky130_fd_sc_hd__or3_4 _2784_ (.A(_1818_),
    .B(_1847_),
    .C(_1879_),
    .X(_1880_));
 sky130_fd_sc_hd__and4_4 _2785_ (.A(net249),
    .B(net224),
    .C(net217),
    .D(net151),
    .X(_1881_));
 sky130_fd_sc_hd__a22o_1 _2786_ (.A1(net66),
    .A2(_1600_),
    .B1(net20),
    .B2(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__o21a_1 _2787_ (.A1(_1283_),
    .A2(_1443_),
    .B1(net55),
    .X(_1883_));
 sky130_fd_sc_hd__o21a_1 _2788_ (.A1(_1320_),
    .A2(_1763_),
    .B1(net45),
    .X(_1884_));
 sky130_fd_sc_hd__o2111a_4 _2789_ (.A1(net211),
    .A2(net177),
    .B1(net251),
    .C1(net227),
    .D1(net220),
    .X(_1885_));
 sky130_fd_sc_hd__o31a_1 _2790_ (.A1(_1163_),
    .A2(_1323_),
    .A3(_1885_),
    .B1(net33),
    .X(_1886_));
 sky130_fd_sc_hd__a2111o_1 _2791_ (.A1(_1254_),
    .A2(net59),
    .B1(_1883_),
    .C1(_1884_),
    .D1(_1886_),
    .X(_1887_));
 sky130_fd_sc_hd__or2_1 _2792_ (.A(_1882_),
    .B(_1887_),
    .X(_1888_));
 sky130_fd_sc_hd__o31a_1 _2793_ (.A1(_1435_),
    .A2(_1463_),
    .A3(_1635_),
    .B1(net50),
    .X(_1889_));
 sky130_fd_sc_hd__nor2_8 _2794_ (.A(net165),
    .B(_1389_),
    .Y(_1890_));
 sky130_fd_sc_hd__or2_1 _2795_ (.A(_1701_),
    .B(_1890_),
    .X(_1891_));
 sky130_fd_sc_hd__or2_1 _2796_ (.A(_1411_),
    .B(_1457_),
    .X(_1892_));
 sky130_fd_sc_hd__a221o_1 _2797_ (.A1(net65),
    .A2(_1891_),
    .B1(_1892_),
    .B2(net61),
    .C1(_1889_),
    .X(_1893_));
 sky130_fd_sc_hd__or2_1 _2798_ (.A(net94),
    .B(net72),
    .X(_1894_));
 sky130_fd_sc_hd__or4_2 _2799_ (.A(_1561_),
    .B(_1627_),
    .C(net69),
    .D(_1894_),
    .X(_1895_));
 sky130_fd_sc_hd__or3_1 _2800_ (.A(_1590_),
    .B(_1591_),
    .C(_1597_),
    .X(_1896_));
 sky130_fd_sc_hd__or4_2 _2801_ (.A(_1034_),
    .B(_1533_),
    .C(net27),
    .D(_1805_),
    .X(_1897_));
 sky130_fd_sc_hd__or4_1 _2802_ (.A(_1365_),
    .B(_1568_),
    .C(_1895_),
    .D(_1897_),
    .X(_1898_));
 sky130_fd_sc_hd__o21a_1 _2803_ (.A1(_1896_),
    .A2(_1898_),
    .B1(net20),
    .X(_1899_));
 sky130_fd_sc_hd__or2_1 _2804_ (.A(_1559_),
    .B(_1881_),
    .X(_1900_));
 sky130_fd_sc_hd__a22o_1 _2805_ (.A1(net61),
    .A2(_1762_),
    .B1(_1900_),
    .B2(net23),
    .X(_1901_));
 sky130_fd_sc_hd__and3_4 _2806_ (.A(_0605_),
    .B(_1386_),
    .C(_1401_),
    .X(_1902_));
 sky130_fd_sc_hd__o21a_1 _2807_ (.A1(_1464_),
    .A2(_1654_),
    .B1(net25),
    .X(_1903_));
 sky130_fd_sc_hd__a2111o_1 _2808_ (.A1(_1254_),
    .A2(net59),
    .B1(_1883_),
    .C1(_1884_),
    .D1(_1886_),
    .X(_1904_));
 sky130_fd_sc_hd__a2111o_1 _2809_ (.A1(_1829_),
    .A2(_1902_),
    .B1(_1903_),
    .C1(_1893_),
    .D1(_1901_),
    .X(_1905_));
 sky130_fd_sc_hd__or4_2 _2810_ (.A(_1882_),
    .B(_1899_),
    .C(_1904_),
    .D(_1905_),
    .X(_1906_));
 sky130_fd_sc_hd__a22o_2 _2811_ (.A1(net173),
    .A2(net99),
    .B1(net84),
    .B2(net202),
    .X(_1907_));
 sky130_fd_sc_hd__or4_1 _2812_ (.A(_1361_),
    .B(_1423_),
    .C(_1528_),
    .D(_1907_),
    .X(_1908_));
 sky130_fd_sc_hd__or4_1 _2813_ (.A(_1414_),
    .B(_1440_),
    .C(_1570_),
    .D(_1872_),
    .X(_1909_));
 sky130_fd_sc_hd__or4_1 _2814_ (.A(_1368_),
    .B(_1391_),
    .C(_1395_),
    .D(_1431_),
    .X(_1910_));
 sky130_fd_sc_hd__or4_1 _2815_ (.A(_1390_),
    .B(_1754_),
    .C(_1890_),
    .D(_1910_),
    .X(_1911_));
 sky130_fd_sc_hd__o31a_1 _2816_ (.A1(_1908_),
    .A2(_1909_),
    .A3(_1911_),
    .B1(net39),
    .X(_1912_));
 sky130_fd_sc_hd__a21o_1 _2817_ (.A1(net188),
    .A2(net81),
    .B1(_1781_),
    .X(_1913_));
 sky130_fd_sc_hd__or4_1 _2818_ (.A(_1736_),
    .B(_1747_),
    .C(_1767_),
    .D(_1913_),
    .X(_1914_));
 sky130_fd_sc_hd__and4_4 _2819_ (.A(net258),
    .B(net223),
    .C(net158),
    .D(net133),
    .X(_1915_));
 sky130_fd_sc_hd__a21o_1 _2820_ (.A1(net124),
    .A2(net195),
    .B1(_1915_),
    .X(_1916_));
 sky130_fd_sc_hd__or3_1 _2821_ (.A(_1529_),
    .B(_1626_),
    .C(_1916_),
    .X(_1917_));
 sky130_fd_sc_hd__o31a_1 _2822_ (.A1(_1431_),
    .A2(_1851_),
    .A3(_1917_),
    .B1(net64),
    .X(_1918_));
 sky130_fd_sc_hd__o31a_1 _2823_ (.A1(_1347_),
    .A2(_1424_),
    .A3(_1660_),
    .B1(net24),
    .X(_1919_));
 sky130_fd_sc_hd__nor2_8 _2824_ (.A(net115),
    .B(_1253_),
    .Y(_1920_));
 sky130_fd_sc_hd__and3_4 _2825_ (.A(net267),
    .B(_1121_),
    .C(_1252_),
    .X(_1921_));
 sky130_fd_sc_hd__a22o_1 _2826_ (.A1(_1163_),
    .A2(net22),
    .B1(_1921_),
    .B2(net41),
    .X(_1922_));
 sky130_fd_sc_hd__nor2_8 _2827_ (.A(net100),
    .B(net86),
    .Y(_1923_));
 sky130_fd_sc_hd__or3_1 _2828_ (.A(_1296_),
    .B(_1308_),
    .C(_1923_),
    .X(_1924_));
 sky130_fd_sc_hd__o31a_1 _2829_ (.A1(_1376_),
    .A2(_1377_),
    .A3(_1924_),
    .B1(net22),
    .X(_1925_));
 sky130_fd_sc_hd__nor2_8 _2830_ (.A(net175),
    .B(_1477_),
    .Y(_1926_));
 sky130_fd_sc_hd__or4_1 _2831_ (.A(_1279_),
    .B(net94),
    .C(_1305_),
    .D(net13),
    .X(_1927_));
 sky130_fd_sc_hd__o31a_1 _2832_ (.A1(_1767_),
    .A2(_1923_),
    .A3(_1927_),
    .B1(net41),
    .X(_1928_));
 sky130_fd_sc_hd__o21a_1 _2833_ (.A1(net66),
    .A2(net49),
    .B1(_1345_),
    .X(_1929_));
 sky130_fd_sc_hd__a211o_1 _2834_ (.A1(net195),
    .A2(_1288_),
    .B1(_1339_),
    .C1(_1574_),
    .X(_1930_));
 sky130_fd_sc_hd__a21o_2 _2835_ (.A1(net123),
    .A2(net182),
    .B1(_1367_),
    .X(_1931_));
 sky130_fd_sc_hd__or4_1 _2836_ (.A(_1111_),
    .B(_1357_),
    .C(_1930_),
    .D(_1931_),
    .X(_1932_));
 sky130_fd_sc_hd__or3_2 _2837_ (.A(_1423_),
    .B(_1624_),
    .C(net14),
    .X(_1933_));
 sky130_fd_sc_hd__or3_2 _2838_ (.A(net15),
    .B(_1781_),
    .C(_1844_),
    .X(_1934_));
 sky130_fd_sc_hd__o31a_1 _2839_ (.A1(_1932_),
    .A2(_1933_),
    .A3(_1934_),
    .B1(net57),
    .X(_1935_));
 sky130_fd_sc_hd__o2111a_4 _2840_ (.A1(net179),
    .A2(net169),
    .B1(net157),
    .C1(net232),
    .D1(net246),
    .X(_1936_));
 sky130_fd_sc_hd__a21o_1 _2841_ (.A1(net209),
    .A2(net83),
    .B1(_1936_),
    .X(_1937_));
 sky130_fd_sc_hd__or4_1 _2842_ (.A(_1467_),
    .B(_1578_),
    .C(_1890_),
    .D(_1937_),
    .X(_1938_));
 sky130_fd_sc_hd__a22o_2 _2843_ (.A1(_0957_),
    .A2(net179),
    .B1(net99),
    .B2(net196),
    .X(_1939_));
 sky130_fd_sc_hd__a22o_2 _2844_ (.A1(net193),
    .A2(net105),
    .B1(net88),
    .B2(net144),
    .X(_1940_));
 sky130_fd_sc_hd__o41a_1 _2845_ (.A1(_1361_),
    .A2(_1938_),
    .A3(_1939_),
    .A4(_1940_),
    .B1(net17),
    .X(_1941_));
 sky130_fd_sc_hd__a21o_1 _2846_ (.A1(net112),
    .A2(net133),
    .B1(_1707_),
    .X(_1942_));
 sky130_fd_sc_hd__or3_1 _2847_ (.A(net70),
    .B(_1811_),
    .C(_1942_),
    .X(_1943_));
 sky130_fd_sc_hd__or4_1 _2848_ (.A(_1454_),
    .B(_1548_),
    .C(_1552_),
    .D(net14),
    .X(_1944_));
 sky130_fd_sc_hd__o31a_1 _2849_ (.A1(_1931_),
    .A2(_1943_),
    .A3(_1944_),
    .B1(net54),
    .X(_1945_));
 sky130_fd_sc_hd__a32o_1 _2850_ (.A1(net197),
    .A2(_1340_),
    .A3(net33),
    .B1(net75),
    .B2(net48),
    .X(_1946_));
 sky130_fd_sc_hd__a21o_4 _2851_ (.A1(net119),
    .A2(net154),
    .B1(_1699_),
    .X(_1947_));
 sky130_fd_sc_hd__or4_1 _2852_ (.A(_1319_),
    .B(_1345_),
    .C(_1890_),
    .D(_1947_),
    .X(_1948_));
 sky130_fd_sc_hd__o31a_1 _2853_ (.A1(_1222_),
    .A2(_1552_),
    .A3(_1948_),
    .B1(net45),
    .X(_1949_));
 sky130_fd_sc_hd__or2_2 _2854_ (.A(_1360_),
    .B(_1484_),
    .X(_1950_));
 sky130_fd_sc_hd__nor2_8 _2855_ (.A(net127),
    .B(net174),
    .Y(_1951_));
 sky130_fd_sc_hd__or3_2 _2856_ (.A(_1257_),
    .B(_1950_),
    .C(_1951_),
    .X(_1952_));
 sky130_fd_sc_hd__o31a_1 _2857_ (.A1(_1469_),
    .A2(net73),
    .A3(_1952_),
    .B1(net29),
    .X(_1953_));
 sky130_fd_sc_hd__a21o_1 _2858_ (.A1(net129),
    .A2(net180),
    .B1(_1683_),
    .X(_1954_));
 sky130_fd_sc_hd__a21o_4 _2859_ (.A1(net124),
    .A2(net203),
    .B1(_1867_),
    .X(_1955_));
 sky130_fd_sc_hd__or4_2 _2860_ (.A(net72),
    .B(_1690_),
    .C(_1700_),
    .D(net68),
    .X(_1956_));
 sky130_fd_sc_hd__and4_4 _2861_ (.A(net242),
    .B(net255),
    .C(net230),
    .D(net215),
    .X(_1957_));
 sky130_fd_sc_hd__or3_1 _2862_ (.A(_1254_),
    .B(_1629_),
    .C(_1695_),
    .X(_1958_));
 sky130_fd_sc_hd__or4_1 _2863_ (.A(_1624_),
    .B(_1954_),
    .C(_1955_),
    .D(net67),
    .X(_1959_));
 sky130_fd_sc_hd__o31a_1 _2864_ (.A1(_1956_),
    .A2(_1958_),
    .A3(_1959_),
    .B1(net36),
    .X(_1960_));
 sky130_fd_sc_hd__o21ai_1 _2865_ (.A1(_1324_),
    .A2(_1681_),
    .B1(net32),
    .Y(_1961_));
 sky130_fd_sc_hd__a211o_1 _2866_ (.A1(net99),
    .A2(net169),
    .B1(_1339_),
    .C1(_1342_),
    .X(_1962_));
 sky130_fd_sc_hd__o41ai_1 _2867_ (.A1(_1555_),
    .A2(_1557_),
    .A3(_1629_),
    .A4(_1962_),
    .B1(net50),
    .Y(_1963_));
 sky130_fd_sc_hd__nand2_1 _2868_ (.A(_1961_),
    .B(_1963_),
    .Y(_1964_));
 sky130_fd_sc_hd__or4_1 _2869_ (.A(_1922_),
    .B(_1941_),
    .C(_1960_),
    .D(_1964_),
    .X(_1965_));
 sky130_fd_sc_hd__a221o_1 _2870_ (.A1(net53),
    .A2(_1388_),
    .B1(_1914_),
    .B2(net63),
    .C1(_1929_),
    .X(_1966_));
 sky130_fd_sc_hd__or3_1 _2871_ (.A(_1949_),
    .B(_1953_),
    .C(_1966_),
    .X(_1967_));
 sky130_fd_sc_hd__or4_1 _2872_ (.A(_1912_),
    .B(_1918_),
    .C(_1919_),
    .D(_1945_),
    .X(_1968_));
 sky130_fd_sc_hd__or4_1 _2873_ (.A(_1925_),
    .B(_1928_),
    .C(_1935_),
    .D(_1946_),
    .X(_1969_));
 sky130_fd_sc_hd__or4_4 _2874_ (.A(_1965_),
    .B(_1967_),
    .C(_1968_),
    .D(_1969_),
    .X(_1970_));
 sky130_fd_sc_hd__or2_2 _2875_ (.A(_1635_),
    .B(_1639_),
    .X(_1971_));
 sky130_fd_sc_hd__a21oi_1 _2876_ (.A1(net192),
    .A2(net150),
    .B1(net80),
    .Y(_1972_));
 sky130_fd_sc_hd__or2_1 _2877_ (.A(_1627_),
    .B(_1744_),
    .X(_1973_));
 sky130_fd_sc_hd__o31a_1 _2878_ (.A1(net14),
    .A2(_1972_),
    .A3(_1973_),
    .B1(net38),
    .X(_1974_));
 sky130_fd_sc_hd__o21a_1 _2879_ (.A1(_0979_),
    .A2(_1479_),
    .B1(net61),
    .X(_1975_));
 sky130_fd_sc_hd__a22o_1 _2880_ (.A1(net129),
    .A2(net210),
    .B1(net183),
    .B2(net99),
    .X(_1976_));
 sky130_fd_sc_hd__or4_1 _2881_ (.A(_1316_),
    .B(_1574_),
    .C(_1575_),
    .D(_1976_),
    .X(_1977_));
 sky130_fd_sc_hd__o21a_1 _2882_ (.A1(_1331_),
    .A2(_1977_),
    .B1(net35),
    .X(_1978_));
 sky130_fd_sc_hd__a2111o_2 _2883_ (.A1(net43),
    .A2(_1971_),
    .B1(_1974_),
    .C1(_1975_),
    .D1(_1978_),
    .X(_1979_));
 sky130_fd_sc_hd__o21a_1 _2884_ (.A1(_1377_),
    .A2(_1539_),
    .B1(net43),
    .X(_1980_));
 sky130_fd_sc_hd__a2111o_1 _2885_ (.A1(_1727_),
    .A2(_1902_),
    .B1(_1970_),
    .C1(_1979_),
    .D1(_1980_),
    .X(_1981_));
 sky130_fd_sc_hd__or4_1 _2886_ (.A(_1780_),
    .B(_1880_),
    .C(_1906_),
    .D(_1981_),
    .X(_1982_));
 sky130_fd_sc_hd__nor2_8 _2887_ (.A(net126),
    .B(net185),
    .Y(_1983_));
 sky130_fd_sc_hd__or2_1 _2888_ (.A(_1365_),
    .B(_1983_),
    .X(_1984_));
 sky130_fd_sc_hd__nor2_8 _2889_ (.A(net118),
    .B(net165),
    .Y(_1985_));
 sky130_fd_sc_hd__or2_2 _2890_ (.A(net13),
    .B(_1985_),
    .X(_1986_));
 sky130_fd_sc_hd__a21oi_1 _2891_ (.A1(net186),
    .A2(net150),
    .B1(_1023_),
    .Y(_1987_));
 sky130_fd_sc_hd__or3_1 _2892_ (.A(_1568_),
    .B(_1890_),
    .C(_1987_),
    .X(_1988_));
 sky130_fd_sc_hd__or4_4 _2893_ (.A(_1360_),
    .B(_1881_),
    .C(_1937_),
    .D(_1984_),
    .X(_1989_));
 sky130_fd_sc_hd__or3_1 _2894_ (.A(_1986_),
    .B(_1988_),
    .C(_1989_),
    .X(_1990_));
 sky130_fd_sc_hd__a21oi_2 _2895_ (.A1(net241),
    .A2(net201),
    .B1(net95),
    .Y(_1991_));
 sky130_fd_sc_hd__a21o_4 _2896_ (.A1(net242),
    .A2(net81),
    .B1(_1406_),
    .X(_1992_));
 sky130_fd_sc_hd__or4_1 _2897_ (.A(_1283_),
    .B(_1561_),
    .C(_1955_),
    .D(_1991_),
    .X(_1993_));
 sky130_fd_sc_hd__or4_1 _2898_ (.A(_1325_),
    .B(_1635_),
    .C(_1992_),
    .D(_1993_),
    .X(_1994_));
 sky130_fd_sc_hd__o21a_1 _2899_ (.A1(_1464_),
    .A2(_1687_),
    .B1(net51),
    .X(_1995_));
 sky130_fd_sc_hd__or2_2 _2900_ (.A(_1163_),
    .B(_1851_),
    .X(_1996_));
 sky130_fd_sc_hd__or3_1 _2901_ (.A(_1500_),
    .B(_1529_),
    .C(_1996_),
    .X(_1997_));
 sky130_fd_sc_hd__a221o_1 _2902_ (.A1(net38),
    .A2(_1994_),
    .B1(_1997_),
    .B2(net20),
    .C1(_1995_),
    .X(_1998_));
 sky130_fd_sc_hd__o21a_1 _2903_ (.A1(_1443_),
    .A2(_1641_),
    .B1(net57),
    .X(_1999_));
 sky130_fd_sc_hd__o41a_1 _2904_ (.A1(_1442_),
    .A2(_1459_),
    .A3(net14),
    .A4(_1872_),
    .B1(_1403_),
    .X(_2000_));
 sky130_fd_sc_hd__o41a_1 _2905_ (.A1(_1111_),
    .A2(_1163_),
    .A3(_1254_),
    .A4(_1622_),
    .B1(net63),
    .X(_2001_));
 sky130_fd_sc_hd__o31a_1 _2906_ (.A1(_1411_),
    .A2(net14),
    .A3(_1872_),
    .B1(net45),
    .X(_2002_));
 sky130_fd_sc_hd__or4_1 _2907_ (.A(_1999_),
    .B(_2000_),
    .C(_2001_),
    .D(_2002_),
    .X(_2003_));
 sky130_fd_sc_hd__a21o_1 _2908_ (.A1(net119),
    .A2(net139),
    .B1(_1460_),
    .X(_2004_));
 sky130_fd_sc_hd__o31a_1 _2909_ (.A1(_1410_),
    .A2(_1467_),
    .A3(_2004_),
    .B1(net25),
    .X(_2005_));
 sky130_fd_sc_hd__o41a_1 _2910_ (.A1(_1460_),
    .A2(net73),
    .A3(_1654_),
    .A4(_1660_),
    .B1(net22),
    .X(_2006_));
 sky130_fd_sc_hd__a21o_2 _2911_ (.A1(net129),
    .A2(net145),
    .B1(_1544_),
    .X(_2007_));
 sky130_fd_sc_hd__o221a_2 _2912_ (.A1(net126),
    .A2(net192),
    .B1(net132),
    .B2(net116),
    .C1(_1594_),
    .X(_2008_));
 sky130_fd_sc_hd__inv_2 _2913_ (.A(_2008_),
    .Y(_2009_));
 sky130_fd_sc_hd__o41a_1 _2914_ (.A1(_1590_),
    .A2(_1593_),
    .A3(_1736_),
    .A4(_2007_),
    .B1(net35),
    .X(_2010_));
 sky130_fd_sc_hd__a2111o_1 _2915_ (.A1(net35),
    .A2(_1498_),
    .B1(_2005_),
    .C1(_2006_),
    .D1(_2010_),
    .X(_2011_));
 sky130_fd_sc_hd__o41a_1 _2916_ (.A1(_0979_),
    .A2(_1518_),
    .A3(_1589_),
    .A4(_1789_),
    .B1(net24),
    .X(_2012_));
 sky130_fd_sc_hd__a2111o_1 _2917_ (.A1(net198),
    .A2(net81),
    .B1(_1708_),
    .C1(_1713_),
    .D1(_1381_),
    .X(_2013_));
 sky130_fd_sc_hd__a21oi_4 _2918_ (.A1(net92),
    .A2(_1303_),
    .B1(net104),
    .Y(_2014_));
 sky130_fd_sc_hd__o31a_1 _2919_ (.A1(_1781_),
    .A2(net69),
    .A3(_2014_),
    .B1(net54),
    .X(_2015_));
 sky130_fd_sc_hd__and4_4 _2920_ (.A(net256),
    .B(net231),
    .C(net180),
    .D(net156),
    .X(_2016_));
 sky130_fd_sc_hd__nor2_1 _2921_ (.A(net115),
    .B(net111),
    .Y(_2017_));
 sky130_fd_sc_hd__a21o_2 _2922_ (.A1(net197),
    .A2(net112),
    .B1(_2016_),
    .X(_2018_));
 sky130_fd_sc_hd__o31a_1 _2923_ (.A1(_1283_),
    .A2(_1526_),
    .A3(_2018_),
    .B1(net29),
    .X(_2019_));
 sky130_fd_sc_hd__a2111o_2 _2924_ (.A1(net51),
    .A2(_2013_),
    .B1(_2015_),
    .C1(_2019_),
    .D1(_2012_),
    .X(_2020_));
 sky130_fd_sc_hd__o41a_1 _2925_ (.A1(_1163_),
    .A2(_1280_),
    .A3(net74),
    .A4(net71),
    .B1(net57),
    .X(_2021_));
 sky130_fd_sc_hd__o41a_1 _2926_ (.A1(_1254_),
    .A2(_1614_),
    .A3(_1639_),
    .A4(_1942_),
    .B1(net41),
    .X(_2022_));
 sky130_fd_sc_hd__o21a_1 _2927_ (.A1(_1308_),
    .A2(_1629_),
    .B1(net38),
    .X(_2023_));
 sky130_fd_sc_hd__o41a_1 _2928_ (.A1(_1405_),
    .A2(_1495_),
    .A3(_1498_),
    .A4(_1827_),
    .B1(net65),
    .X(_2024_));
 sky130_fd_sc_hd__or4_1 _2929_ (.A(_2021_),
    .B(_2022_),
    .C(_2023_),
    .D(_2024_),
    .X(_2025_));
 sky130_fd_sc_hd__or4_4 _2930_ (.A(_2003_),
    .B(_2011_),
    .C(_2020_),
    .D(_2025_),
    .X(_2027_));
 sky130_fd_sc_hd__a211oi_2 _2931_ (.A1(net37),
    .A2(_1990_),
    .B1(_1998_),
    .C1(_2027_),
    .Y(_2028_));
 sky130_fd_sc_hd__a22o_1 _2932_ (.A1(net181),
    .A2(net90),
    .B1(net139),
    .B2(net112),
    .X(_2029_));
 sky130_fd_sc_hd__or4_1 _2933_ (.A(_1467_),
    .B(_1627_),
    .C(_1920_),
    .D(_2029_),
    .X(_2030_));
 sky130_fd_sc_hd__a22o_1 _2934_ (.A1(_1354_),
    .A2(net40),
    .B1(net37),
    .B2(_2030_),
    .X(_2031_));
 sky130_fd_sc_hd__or4_1 _2935_ (.A(_1480_),
    .B(_1583_),
    .C(_1626_),
    .D(_1916_),
    .X(_2032_));
 sky130_fd_sc_hd__a211o_1 _2936_ (.A1(net197),
    .A2(_1340_),
    .B1(_1494_),
    .C1(_1324_),
    .X(_2033_));
 sky130_fd_sc_hd__or4_1 _2937_ (.A(_0935_),
    .B(_1283_),
    .C(_1920_),
    .D(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__a22o_1 _2938_ (.A1(net17),
    .A2(_2032_),
    .B1(_2034_),
    .B2(net21),
    .X(_2035_));
 sky130_fd_sc_hd__a211o_1 _2939_ (.A1(net210),
    .A2(net124),
    .B1(_1339_),
    .C1(_1342_),
    .X(_2036_));
 sky130_fd_sc_hd__o31a_1 _2940_ (.A1(_1243_),
    .A2(_1538_),
    .A3(_2036_),
    .B1(net32),
    .X(_0051_));
 sky130_fd_sc_hd__o31a_1 _2941_ (.A1(_1431_),
    .A2(net74),
    .A3(net67),
    .B1(net48),
    .X(_0052_));
 sky130_fd_sc_hd__o31a_1 _2942_ (.A1(_1363_),
    .A2(net75),
    .A3(_1849_),
    .B1(net44),
    .X(_0053_));
 sky130_fd_sc_hd__a2111o_1 _2943_ (.A1(net51),
    .A2(_1395_),
    .B1(_0051_),
    .C1(_0052_),
    .D1(_0053_),
    .X(_0054_));
 sky130_fd_sc_hd__or4_1 _2944_ (.A(_1296_),
    .B(_1417_),
    .C(_1649_),
    .D(net68),
    .X(_0055_));
 sky130_fd_sc_hd__o41a_1 _2945_ (.A1(net71),
    .A2(_1559_),
    .A3(_1709_),
    .A4(_1713_),
    .B1(net29),
    .X(_0056_));
 sky130_fd_sc_hd__a221oi_1 _2946_ (.A1(net64),
    .A2(_1690_),
    .B1(_0055_),
    .B2(net39),
    .C1(_0056_),
    .Y(_0057_));
 sky130_fd_sc_hd__o2111a_1 _2947_ (.A1(net244),
    .A2(net197),
    .B1(net219),
    .C1(net239),
    .D1(net250),
    .X(_0058_));
 sky130_fd_sc_hd__or3_1 _2948_ (.A(_1366_),
    .B(net67),
    .C(_0058_),
    .X(_0059_));
 sky130_fd_sc_hd__a22o_1 _2949_ (.A1(net41),
    .A2(_1478_),
    .B1(_0059_),
    .B2(net39),
    .X(_0060_));
 sky130_fd_sc_hd__a21o_1 _2950_ (.A1(net183),
    .A2(net90),
    .B1(_1424_),
    .X(_0062_));
 sky130_fd_sc_hd__o41a_1 _2951_ (.A1(_1410_),
    .A2(net76),
    .A3(net15),
    .A4(_0062_),
    .B1(net53),
    .X(_0063_));
 sky130_fd_sc_hd__or4_1 _2952_ (.A(_0935_),
    .B(_1376_),
    .C(net75),
    .D(net73),
    .X(_0064_));
 sky130_fd_sc_hd__a211oi_1 _2953_ (.A1(net58),
    .A2(_0064_),
    .B1(_0063_),
    .C1(_0060_),
    .Y(_0065_));
 sky130_fd_sc_hd__or4bb_4 _2954_ (.A(_2035_),
    .B(_0054_),
    .C_N(_0057_),
    .D_N(_0065_),
    .X(_0066_));
 sky130_fd_sc_hd__or2_1 _2955_ (.A(_2031_),
    .B(_0066_),
    .X(_0067_));
 sky130_fd_sc_hd__and2_1 _2956_ (.A(net55),
    .B(_1459_),
    .X(_0068_));
 sky130_fd_sc_hd__o21a_1 _2957_ (.A1(_1452_),
    .A2(_1746_),
    .B1(net61),
    .X(_0069_));
 sky130_fd_sc_hd__o21a_1 _2958_ (.A1(_1544_),
    .A2(net15),
    .B1(net65),
    .X(_0070_));
 sky130_fd_sc_hd__a211o_1 _2959_ (.A1(net45),
    .A2(_1550_),
    .B1(_0069_),
    .C1(_0070_),
    .X(_0071_));
 sky130_fd_sc_hd__a221o_2 _2960_ (.A1(_1521_),
    .A2(_1606_),
    .B1(net16),
    .B2(net60),
    .C1(_0071_),
    .X(_0073_));
 sky130_fd_sc_hd__a22o_1 _2961_ (.A1(net45),
    .A2(_1479_),
    .B1(net31),
    .B2(_1445_),
    .X(_0074_));
 sky130_fd_sc_hd__a22o_1 _2962_ (.A1(net52),
    .A2(_1564_),
    .B1(_1695_),
    .B2(net66),
    .X(_0075_));
 sky130_fd_sc_hd__a221oi_4 _2963_ (.A1(_1274_),
    .A2(net59),
    .B1(_1322_),
    .B2(net56),
    .C1(_0075_),
    .Y(_0076_));
 sky130_fd_sc_hd__a21oi_4 _2964_ (.A1(net108),
    .A2(net100),
    .B1(net85),
    .Y(_0077_));
 sky130_fd_sc_hd__a21oi_4 _2965_ (.A1(net114),
    .A2(_1303_),
    .B1(net103),
    .Y(_0078_));
 sky130_fd_sc_hd__or2_4 _2966_ (.A(_0077_),
    .B(_0078_),
    .X(_0079_));
 sky130_fd_sc_hd__a22o_1 _2967_ (.A1(_1441_),
    .A2(net31),
    .B1(_0079_),
    .B2(_1403_),
    .X(_0080_));
 sky130_fd_sc_hd__nand2_1 _2968_ (.A(net82),
    .B(net46),
    .Y(_0081_));
 sky130_fd_sc_hd__or4_2 _2969_ (.A(_1606_),
    .B(net68),
    .C(_1957_),
    .D(_2016_),
    .X(_0082_));
 sky130_fd_sc_hd__and4_4 _2970_ (.A(net255),
    .B(net222),
    .C(net179),
    .D(net156),
    .X(_0084_));
 sky130_fd_sc_hd__nor2_8 _2971_ (.A(net121),
    .B(net166),
    .Y(_0085_));
 sky130_fd_sc_hd__a21o_4 _2972_ (.A1(net123),
    .A2(net169),
    .B1(_0084_),
    .X(_0086_));
 sky130_fd_sc_hd__nor2_1 _2973_ (.A(_1867_),
    .B(_0084_),
    .Y(_0087_));
 sky130_fd_sc_hd__a21oi_4 _2974_ (.A1(net199),
    .A2(net166),
    .B1(net122),
    .Y(_0088_));
 sky130_fd_sc_hd__o31a_1 _2975_ (.A1(_1955_),
    .A2(_0082_),
    .A3(_0086_),
    .B1(net62),
    .X(_0089_));
 sky130_fd_sc_hd__or4bb_1 _2976_ (.A(_0089_),
    .B(_0080_),
    .C_N(_0076_),
    .D_N(_0081_),
    .X(_0090_));
 sky130_fd_sc_hd__or4_1 _2977_ (.A(_0068_),
    .B(_0073_),
    .C(_0074_),
    .D(_0090_),
    .X(_0091_));
 sky130_fd_sc_hd__nor2_1 _2978_ (.A(_0067_),
    .B(_0091_),
    .Y(_0092_));
 sky130_fd_sc_hd__nand2_1 _2979_ (.A(_2028_),
    .B(_0092_),
    .Y(_0093_));
 sky130_fd_sc_hd__o21a_1 _2980_ (.A1(_1583_),
    .A2(_1713_),
    .B1(net39),
    .X(_0095_));
 sky130_fd_sc_hd__a21o_1 _2981_ (.A1(net123),
    .A2(net187),
    .B1(_1618_),
    .X(_0096_));
 sky130_fd_sc_hd__o21a_1 _2982_ (.A1(_1414_),
    .A2(_1538_),
    .B1(net57),
    .X(_0097_));
 sky130_fd_sc_hd__o41a_1 _2983_ (.A1(_1494_),
    .A2(_1517_),
    .A3(_1597_),
    .A4(_1618_),
    .B1(net39),
    .X(_0098_));
 sky130_fd_sc_hd__o41a_1 _2984_ (.A1(_1322_),
    .A2(_1390_),
    .A3(_1679_),
    .A4(_1696_),
    .B1(net19),
    .X(_0099_));
 sky130_fd_sc_hd__o31a_1 _2985_ (.A1(_1701_),
    .A2(_1876_),
    .A3(net67),
    .B1(net50),
    .X(_0100_));
 sky130_fd_sc_hd__o21a_1 _2986_ (.A1(_1280_),
    .A2(_1915_),
    .B1(net54),
    .X(_0101_));
 sky130_fd_sc_hd__or3_4 _2987_ (.A(_1380_),
    .B(_1381_),
    .C(_1690_),
    .X(_0102_));
 sky130_fd_sc_hd__o31a_1 _2988_ (.A1(net75),
    .A2(_1445_),
    .A3(_1985_),
    .B1(net64),
    .X(_0103_));
 sky130_fd_sc_hd__o31a_1 _2989_ (.A1(_0979_),
    .A2(_1345_),
    .A3(_1367_),
    .B1(net32),
    .X(_0104_));
 sky130_fd_sc_hd__a211o_1 _2990_ (.A1(net244),
    .A2(net120),
    .B1(net70),
    .C1(_1624_),
    .X(_0106_));
 sky130_fd_sc_hd__a22o_4 _2991_ (.A1(net120),
    .A2(net173),
    .B1(net98),
    .B2(net146),
    .X(_0107_));
 sky130_fd_sc_hd__or2_4 _2992_ (.A(_1296_),
    .B(_1699_),
    .X(_0108_));
 sky130_fd_sc_hd__o21a_1 _2993_ (.A1(_1452_),
    .A2(_1781_),
    .B1(net32),
    .X(_0109_));
 sky130_fd_sc_hd__o31a_1 _2994_ (.A1(_1291_),
    .A2(net94),
    .A3(_1700_),
    .B1(net54),
    .X(_0110_));
 sky130_fd_sc_hd__or3_1 _2995_ (.A(_1222_),
    .B(_1459_),
    .C(_1872_),
    .X(_0111_));
 sky130_fd_sc_hd__a22o_1 _2996_ (.A1(net76),
    .A2(net24),
    .B1(net17),
    .B2(_0111_),
    .X(_0112_));
 sky130_fd_sc_hd__o31a_1 _2997_ (.A1(_1271_),
    .A2(_1320_),
    .A3(_1339_),
    .B1(net19),
    .X(_0113_));
 sky130_fd_sc_hd__a22o_1 _2998_ (.A1(net44),
    .A2(_1494_),
    .B1(_1577_),
    .B2(net21),
    .X(_0114_));
 sky130_fd_sc_hd__or4_1 _2999_ (.A(_0109_),
    .B(_0110_),
    .C(_0113_),
    .D(_0114_),
    .X(_0115_));
 sky130_fd_sc_hd__a22o_1 _3000_ (.A1(net22),
    .A2(_1624_),
    .B1(_1689_),
    .B2(net50),
    .X(_0117_));
 sky130_fd_sc_hd__o21a_1 _3001_ (.A1(_1552_),
    .A2(_0084_),
    .B1(net42),
    .X(_0118_));
 sky130_fd_sc_hd__a211oi_1 _3002_ (.A1(net32),
    .A2(_1722_),
    .B1(_0117_),
    .C1(_0118_),
    .Y(_0119_));
 sky130_fd_sc_hd__a22o_1 _3003_ (.A1(net44),
    .A2(_1445_),
    .B1(net29),
    .B2(_1753_),
    .X(_0120_));
 sky130_fd_sc_hd__a22o_1 _3004_ (.A1(net119),
    .A2(net182),
    .B1(net105),
    .B2(net138),
    .X(_0121_));
 sky130_fd_sc_hd__o31a_1 _3005_ (.A1(_1849_),
    .A2(_1939_),
    .A3(_0121_),
    .B1(net36),
    .X(_0122_));
 sky130_fd_sc_hd__a211oi_1 _3006_ (.A1(_1034_),
    .A2(net57),
    .B1(_0120_),
    .C1(_0122_),
    .Y(_0123_));
 sky130_fd_sc_hd__or4bb_1 _3007_ (.A(_0112_),
    .B(_0115_),
    .C_N(_0119_),
    .D_N(_0123_),
    .X(_0124_));
 sky130_fd_sc_hd__o31a_1 _3008_ (.A1(net70),
    .A2(_1811_),
    .A3(_2018_),
    .B1(net42),
    .X(_0125_));
 sky130_fd_sc_hd__a211o_1 _3009_ (.A1(_1388_),
    .A2(net36),
    .B1(_0103_),
    .C1(_0125_),
    .X(_0126_));
 sky130_fd_sc_hd__a221o_1 _3010_ (.A1(net43),
    .A2(_1440_),
    .B1(_0102_),
    .B2(net54),
    .C1(_0104_),
    .X(_0128_));
 sky130_fd_sc_hd__or4_1 _3011_ (.A(_0097_),
    .B(_0098_),
    .C(_0126_),
    .D(_0128_),
    .X(_0129_));
 sky130_fd_sc_hd__or3_2 _3012_ (.A(_1397_),
    .B(_1457_),
    .C(_1466_),
    .X(_0130_));
 sky130_fd_sc_hd__a221o_1 _3013_ (.A1(net30),
    .A2(_0106_),
    .B1(_0130_),
    .B2(net25),
    .C1(_0100_),
    .X(_0131_));
 sky130_fd_sc_hd__a221o_2 _3014_ (.A1(_1349_),
    .A2(net44),
    .B1(_1699_),
    .B2(net48),
    .C1(_0099_),
    .X(_0132_));
 sky130_fd_sc_hd__a22o_1 _3015_ (.A1(net57),
    .A2(_1421_),
    .B1(_1488_),
    .B2(net63),
    .X(_0133_));
 sky130_fd_sc_hd__a211o_1 _3016_ (.A1(_1394_),
    .A2(net24),
    .B1(_0095_),
    .C1(_0133_),
    .X(_0134_));
 sky130_fd_sc_hd__a22o_1 _3017_ (.A1(net21),
    .A2(_0107_),
    .B1(_0108_),
    .B2(net17),
    .X(_0135_));
 sky130_fd_sc_hd__a211o_1 _3018_ (.A1(net29),
    .A2(_0096_),
    .B1(_0101_),
    .C1(_0135_),
    .X(_0136_));
 sky130_fd_sc_hd__or4_1 _3019_ (.A(_0131_),
    .B(_0132_),
    .C(_0134_),
    .D(_0136_),
    .X(_0137_));
 sky130_fd_sc_hd__or3_4 _3020_ (.A(_0124_),
    .B(_0129_),
    .C(_0137_),
    .X(_0139_));
 sky130_fd_sc_hd__o21a_1 _3021_ (.A1(_1548_),
    .A2(_1578_),
    .B1(net36),
    .X(_0140_));
 sky130_fd_sc_hd__a22o_4 _3022_ (.A1(net129),
    .A2(net204),
    .B1(net120),
    .B2(net140),
    .X(_0141_));
 sky130_fd_sc_hd__a211o_1 _3023_ (.A1(net202),
    .A2(net119),
    .B1(_1357_),
    .C1(_1431_),
    .X(_0142_));
 sky130_fd_sc_hd__o31a_1 _3024_ (.A1(net15),
    .A2(_0141_),
    .A3(_0142_),
    .B1(net32),
    .X(_0143_));
 sky130_fd_sc_hd__a211o_1 _3025_ (.A1(net54),
    .A2(_1357_),
    .B1(_0140_),
    .C1(_0143_),
    .X(_0144_));
 sky130_fd_sc_hd__a221o_1 _3026_ (.A1(net123),
    .A2(net187),
    .B1(net99),
    .B2(net196),
    .C1(_1517_),
    .X(_0145_));
 sky130_fd_sc_hd__o31a_1 _3027_ (.A1(_1583_),
    .A2(_1626_),
    .A3(_0145_),
    .B1(net44),
    .X(_0146_));
 sky130_fd_sc_hd__a32o_1 _3028_ (.A1(net196),
    .A2(net81),
    .A3(net17),
    .B1(_1983_),
    .B2(net64),
    .X(_0147_));
 sky130_fd_sc_hd__a211o_1 _3029_ (.A1(net193),
    .A2(_1288_),
    .B1(_1501_),
    .C1(_1565_),
    .X(_0148_));
 sky130_fd_sc_hd__o21a_1 _3030_ (.A1(_1552_),
    .A2(_2017_),
    .B1(net48),
    .X(_0150_));
 sky130_fd_sc_hd__a211o_1 _3031_ (.A1(net21),
    .A2(_0148_),
    .B1(_0150_),
    .C1(_0147_),
    .X(_0151_));
 sky130_fd_sc_hd__a2111o_4 _3032_ (.A1(net51),
    .A2(net68),
    .B1(_0144_),
    .C1(_0146_),
    .D1(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__nand2_1 _3033_ (.A(_1282_),
    .B(net56),
    .Y(_0153_));
 sky130_fd_sc_hd__a22o_1 _3034_ (.A1(_1375_),
    .A2(net18),
    .B1(net13),
    .B2(net22),
    .X(_0154_));
 sky130_fd_sc_hd__a22o_1 _3035_ (.A1(net198),
    .A2(_1340_),
    .B1(net81),
    .B2(net181),
    .X(_0155_));
 sky130_fd_sc_hd__a22o_1 _3036_ (.A1(net61),
    .A2(_1951_),
    .B1(_0155_),
    .B2(net25),
    .X(_0156_));
 sky130_fd_sc_hd__a22o_1 _3037_ (.A1(net45),
    .A2(net70),
    .B1(_1649_),
    .B2(net43),
    .X(_0157_));
 sky130_fd_sc_hd__or4b_2 _3038_ (.A(_0154_),
    .B(_0156_),
    .C(_0157_),
    .D_N(_0153_),
    .X(_0158_));
 sky130_fd_sc_hd__o41a_1 _3039_ (.A1(net74),
    .A2(_1920_),
    .A3(_1923_),
    .A4(net13),
    .B1(net65),
    .X(_0159_));
 sky130_fd_sc_hd__or4_4 _3040_ (.A(_1309_),
    .B(_1470_),
    .C(_1525_),
    .D(_1626_),
    .X(_0161_));
 sky130_fd_sc_hd__o31ai_1 _3041_ (.A1(_1304_),
    .A2(_1529_),
    .A3(_0161_),
    .B1(net53),
    .Y(_0162_));
 sky130_fd_sc_hd__o21a_1 _3042_ (.A1(_1222_),
    .A2(_2016_),
    .B1(net48),
    .X(_0163_));
 sky130_fd_sc_hd__o41a_1 _3043_ (.A1(_1420_),
    .A2(_1557_),
    .A3(_1570_),
    .A4(_1754_),
    .B1(net18),
    .X(_0164_));
 sky130_fd_sc_hd__and2_1 _3044_ (.A(net61),
    .B(_1486_),
    .X(_0165_));
 sky130_fd_sc_hd__a2111o_1 _3045_ (.A1(_1264_),
    .A2(net38),
    .B1(_0163_),
    .C1(_0164_),
    .D1(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__or4b_4 _3046_ (.A(_0158_),
    .B(_0159_),
    .C(_0166_),
    .D_N(_0162_),
    .X(_0167_));
 sky130_fd_sc_hd__or2_1 _3047_ (.A(_1406_),
    .B(_1417_),
    .X(_0168_));
 sky130_fd_sc_hd__or2_1 _3048_ (.A(_1802_),
    .B(_1851_),
    .X(_0169_));
 sky130_fd_sc_hd__a22o_1 _3049_ (.A1(net45),
    .A2(_0168_),
    .B1(_0169_),
    .B2(net50),
    .X(_0170_));
 sky130_fd_sc_hd__a221o_4 _3050_ (.A1(net53),
    .A2(_1872_),
    .B1(_0086_),
    .B2(net30),
    .C1(_0170_),
    .X(_0171_));
 sky130_fd_sc_hd__a22o_1 _3051_ (.A1(_1309_),
    .A2(net59),
    .B1(_1844_),
    .B2(net66),
    .X(_0172_));
 sky130_fd_sc_hd__or2_1 _3052_ (.A(_1565_),
    .B(_1805_),
    .X(_0173_));
 sky130_fd_sc_hd__a21o_2 _3053_ (.A1(net99),
    .A2(_1326_),
    .B1(_1413_),
    .X(_0174_));
 sky130_fd_sc_hd__a22o_2 _3054_ (.A1(net205),
    .A2(net89),
    .B1(net147),
    .B2(_1408_),
    .X(_0175_));
 sky130_fd_sc_hd__or4_1 _3055_ (.A(_1424_),
    .B(_1644_),
    .C(_0174_),
    .D(_0175_),
    .X(_0176_));
 sky130_fd_sc_hd__a22o_1 _3056_ (.A1(net55),
    .A2(_0173_),
    .B1(_0176_),
    .B2(net37),
    .X(_0177_));
 sky130_fd_sc_hd__or3_1 _3057_ (.A(_0935_),
    .B(_1342_),
    .C(_1763_),
    .X(_0178_));
 sky130_fd_sc_hd__or2_2 _3058_ (.A(_1395_),
    .B(_1680_),
    .X(_0179_));
 sky130_fd_sc_hd__o41a_1 _3059_ (.A1(_1368_),
    .A2(_1555_),
    .A3(_0178_),
    .A4(_0179_),
    .B1(net19),
    .X(_0180_));
 sky130_fd_sc_hd__o21a_1 _3060_ (.A1(_1591_),
    .A2(_1700_),
    .B1(_0627_),
    .X(_0182_));
 sky130_fd_sc_hd__or4_1 _3061_ (.A(_0172_),
    .B(_0177_),
    .C(_0180_),
    .D(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__or4_1 _3062_ (.A(_0152_),
    .B(_0167_),
    .C(_0171_),
    .D(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__or4_1 _3063_ (.A(_1982_),
    .B(_0093_),
    .C(_0139_),
    .D(_0184_),
    .X(_0047_));
 sky130_fd_sc_hd__a31o_2 _3064_ (.A1(net174),
    .A2(net170),
    .A3(net167),
    .B1(_1477_),
    .X(_0185_));
 sky130_fd_sc_hd__or3b_1 _3065_ (.A(_1373_),
    .B(_1593_),
    .C_N(_0185_),
    .X(_0186_));
 sky130_fd_sc_hd__or4_2 _3066_ (.A(_1388_),
    .B(net72),
    .C(_1548_),
    .D(_0062_),
    .X(_0187_));
 sky130_fd_sc_hd__o31a_1 _3067_ (.A1(_0174_),
    .A2(_0186_),
    .A3(_0187_),
    .B1(net62),
    .X(_0188_));
 sky130_fd_sc_hd__or2_1 _3068_ (.A(_1860_),
    .B(_1955_),
    .X(_0189_));
 sky130_fd_sc_hd__or3_1 _3069_ (.A(_1510_),
    .B(_1793_),
    .C(net68),
    .X(_0190_));
 sky130_fd_sc_hd__or4_1 _3070_ (.A(_1470_),
    .B(_1629_),
    .C(_1983_),
    .D(_1985_),
    .X(_0192_));
 sky130_fd_sc_hd__o31a_1 _3071_ (.A1(_0189_),
    .A2(_0190_),
    .A3(_0192_),
    .B1(net17),
    .X(_0193_));
 sky130_fd_sc_hd__or4_1 _3072_ (.A(_1440_),
    .B(_1489_),
    .C(_1709_),
    .D(net13),
    .X(_0194_));
 sky130_fd_sc_hd__or4_2 _3073_ (.A(_1320_),
    .B(_1722_),
    .C(_1829_),
    .D(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__o31a_1 _3074_ (.A1(_1920_),
    .A2(_2029_),
    .A3(_0195_),
    .B1(net53),
    .X(_0196_));
 sky130_fd_sc_hd__or2_1 _3075_ (.A(_1394_),
    .B(_1397_),
    .X(_0197_));
 sky130_fd_sc_hd__or2_1 _3076_ (.A(net75),
    .B(net74),
    .X(_0198_));
 sky130_fd_sc_hd__or4_1 _3077_ (.A(_1443_),
    .B(_1467_),
    .C(_0197_),
    .D(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__a22o_1 _3078_ (.A1(net41),
    .A2(_1550_),
    .B1(_0199_),
    .B2(net50),
    .X(_0200_));
 sky130_fd_sc_hd__a221o_1 _3079_ (.A1(net188),
    .A2(net105),
    .B1(net99),
    .B2(net203),
    .C1(net94),
    .X(_0201_));
 sky130_fd_sc_hd__or4_1 _3080_ (.A(net16),
    .B(_2018_),
    .C(_0086_),
    .D(_0201_),
    .X(_0203_));
 sky130_fd_sc_hd__o21a_1 _3081_ (.A1(_1405_),
    .A2(_1506_),
    .B1(net48),
    .X(_0204_));
 sky130_fd_sc_hd__or4_1 _3082_ (.A(_1264_),
    .B(_1431_),
    .C(_1484_),
    .D(_1660_),
    .X(_0205_));
 sky130_fd_sc_hd__a21oi_4 _3083_ (.A1(net176),
    .A2(net132),
    .B1(net126),
    .Y(_0206_));
 sky130_fd_sc_hd__o41a_1 _3084_ (.A1(_1907_),
    .A2(_2007_),
    .A3(_0205_),
    .A4(_0206_),
    .B1(net58),
    .X(_0207_));
 sky130_fd_sc_hd__o41a_1 _3085_ (.A1(_1267_),
    .A2(_1593_),
    .A3(_1683_),
    .A4(_1781_),
    .B1(net64),
    .X(_0208_));
 sky130_fd_sc_hd__or4_1 _3086_ (.A(net27),
    .B(_1654_),
    .C(net16),
    .D(_1744_),
    .X(_0209_));
 sky130_fd_sc_hd__a21o_1 _3087_ (.A1(net242),
    .A2(net112),
    .B1(net72),
    .X(_0210_));
 sky130_fd_sc_hd__o31a_1 _3088_ (.A1(_1429_),
    .A2(_0209_),
    .A3(_0210_),
    .B1(net44),
    .X(_0211_));
 sky130_fd_sc_hd__or4_1 _3089_ (.A(_1708_),
    .B(_1713_),
    .C(_1746_),
    .D(_1983_),
    .X(_0212_));
 sky130_fd_sc_hd__o31ai_1 _3090_ (.A1(_1510_),
    .A2(_1792_),
    .A3(_0212_),
    .B1(net22),
    .Y(_0214_));
 sky130_fd_sc_hd__o31a_1 _3091_ (.A1(_1243_),
    .A2(_1537_),
    .A3(_1951_),
    .B1(net36),
    .X(_0215_));
 sky130_fd_sc_hd__o41a_1 _3092_ (.A1(net82),
    .A2(_1354_),
    .A3(_1559_),
    .A4(net67),
    .B1(net18),
    .X(_0216_));
 sky130_fd_sc_hd__o41a_1 _3093_ (.A1(_1356_),
    .A2(_1500_),
    .A3(_1639_),
    .A4(_1683_),
    .B1(net39),
    .X(_0217_));
 sky130_fd_sc_hd__nand2b_2 _3094_ (.A_N(_1459_),
    .B(_2008_),
    .Y(_0218_));
 sky130_fd_sc_hd__a22o_1 _3095_ (.A1(net43),
    .A2(_0203_),
    .B1(_0218_),
    .B2(net25),
    .X(_0219_));
 sky130_fd_sc_hd__o31a_1 _3096_ (.A1(_1518_),
    .A2(_1763_),
    .A3(_0086_),
    .B1(net33),
    .X(_0220_));
 sky130_fd_sc_hd__o41a_1 _3097_ (.A1(_1320_),
    .A2(_1347_),
    .A3(_1428_),
    .A4(_1434_),
    .B1(net34),
    .X(_0221_));
 sky130_fd_sc_hd__or4_1 _3098_ (.A(_0204_),
    .B(_0216_),
    .C(_0220_),
    .D(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__or4_1 _3099_ (.A(_0188_),
    .B(_0200_),
    .C(_0219_),
    .D(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__a2111o_1 _3100_ (.A1(net29),
    .A2(_1806_),
    .B1(_0208_),
    .C1(_0215_),
    .D1(_0217_),
    .X(_0225_));
 sky130_fd_sc_hd__or4b_2 _3101_ (.A(_0193_),
    .B(_0211_),
    .C(_0225_),
    .D_N(_0214_),
    .X(_0226_));
 sky130_fd_sc_hd__nor4_2 _3102_ (.A(_0196_),
    .B(_0207_),
    .C(_0223_),
    .D(_0226_),
    .Y(_0227_));
 sky130_fd_sc_hd__nand2_1 _3103_ (.A(_2028_),
    .B(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__a221o_1 _3104_ (.A1(net46),
    .A2(_1488_),
    .B1(net31),
    .B2(_1443_),
    .C1(_0172_),
    .X(_0229_));
 sky130_fd_sc_hd__or2_1 _3105_ (.A(_0171_),
    .B(_0229_),
    .X(_0230_));
 sky130_fd_sc_hd__a211o_1 _3106_ (.A1(_1438_),
    .A2(net31),
    .B1(_0182_),
    .C1(_0230_),
    .X(_0231_));
 sky130_fd_sc_hd__a21o_1 _3107_ (.A1(_1288_),
    .A2(net145),
    .B1(net69),
    .X(_0232_));
 sky130_fd_sc_hd__a22o_2 _3108_ (.A1(net35),
    .A2(_0197_),
    .B1(_0232_),
    .B2(net61),
    .X(_0233_));
 sky130_fd_sc_hd__o21a_1 _3109_ (.A1(_1983_),
    .A2(_1985_),
    .B1(net62),
    .X(_0234_));
 sky130_fd_sc_hd__a21o_1 _3110_ (.A1(_1290_),
    .A2(net46),
    .B1(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__o21a_1 _3111_ (.A1(_1410_),
    .A2(_1414_),
    .B1(net30),
    .X(_0236_));
 sky130_fd_sc_hd__a221o_1 _3112_ (.A1(net46),
    .A2(_1597_),
    .B1(_1881_),
    .B2(net61),
    .C1(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__or4_1 _3113_ (.A(_0231_),
    .B(_0233_),
    .C(_0235_),
    .D(_0237_),
    .X(_0238_));
 sky130_fd_sc_hd__or4_1 _3114_ (.A(_1982_),
    .B(_0067_),
    .C(_0228_),
    .D(_0238_),
    .X(_0048_));
 sky130_fd_sc_hd__o21a_1 _3115_ (.A1(_1690_),
    .A2(_1954_),
    .B1(net50),
    .X(_0239_));
 sky130_fd_sc_hd__o31a_1 _3116_ (.A1(_1282_),
    .A2(_1304_),
    .A3(_1639_),
    .B1(net58),
    .X(_0240_));
 sky130_fd_sc_hd__o31a_2 _3117_ (.A1(_1279_),
    .A2(_1301_),
    .A3(_1374_),
    .B1(net65),
    .X(_0241_));
 sky130_fd_sc_hd__a2111o_1 _3118_ (.A1(net119),
    .A2(net183),
    .B1(net73),
    .C1(_1649_),
    .D1(net13),
    .X(_0242_));
 sky130_fd_sc_hd__or2_4 _3119_ (.A(_1460_),
    .B(_1811_),
    .X(_0243_));
 sky130_fd_sc_hd__o31a_1 _3120_ (.A1(_1991_),
    .A2(_0242_),
    .A3(_0243_),
    .B1(net18),
    .X(_0245_));
 sky130_fd_sc_hd__or4_1 _3121_ (.A(_0239_),
    .B(_0240_),
    .C(_0241_),
    .D(_0245_),
    .X(_0246_));
 sky130_fd_sc_hd__o21a_1 _3122_ (.A1(_1715_),
    .A2(_1792_),
    .B1(net49),
    .X(_0247_));
 sky130_fd_sc_hd__or2_1 _3123_ (.A(_1478_),
    .B(net69),
    .X(_0248_));
 sky130_fd_sc_hd__o31a_1 _3124_ (.A1(_1395_),
    .A2(_1570_),
    .A3(net69),
    .B1(net25),
    .X(_0249_));
 sky130_fd_sc_hd__o41a_4 _3125_ (.A1(_1316_),
    .A2(_1574_),
    .A3(_1575_),
    .A4(_1985_),
    .B1(net21),
    .X(_0250_));
 sky130_fd_sc_hd__a2111o_1 _3126_ (.A1(net33),
    .A2(_0248_),
    .B1(_0249_),
    .C1(_0250_),
    .D1(_0247_),
    .X(_0251_));
 sky130_fd_sc_hd__o211a_1 _3127_ (.A1(net210),
    .A2(net188),
    .B1(net84),
    .C1(net49),
    .X(_0252_));
 sky130_fd_sc_hd__o21a_1 _3128_ (.A1(_1315_),
    .A2(_1590_),
    .B1(net61),
    .X(_0253_));
 sky130_fd_sc_hd__o21a_1 _3129_ (.A1(_1480_),
    .A2(_1583_),
    .B1(net43),
    .X(_0254_));
 sky130_fd_sc_hd__a2111o_1 _3130_ (.A1(net210),
    .A2(net112),
    .B1(_1291_),
    .C1(_1478_),
    .D1(_1518_),
    .X(_0256_));
 sky130_fd_sc_hd__o31a_2 _3131_ (.A1(_1347_),
    .A2(_1423_),
    .A3(_0256_),
    .B1(net37),
    .X(_0257_));
 sky130_fd_sc_hd__or2_1 _3132_ (.A(_1394_),
    .B(_1495_),
    .X(_0258_));
 sky130_fd_sc_hd__o31a_1 _3133_ (.A1(_1267_),
    .A2(_1322_),
    .A3(_0258_),
    .B1(net38),
    .X(_0259_));
 sky130_fd_sc_hd__a211o_4 _3134_ (.A1(net124),
    .A2(net203),
    .B1(_1366_),
    .C1(net67),
    .X(_0260_));
 sky130_fd_sc_hd__o31a_2 _3135_ (.A1(net72),
    .A2(_1867_),
    .A3(_0260_),
    .B1(net30),
    .X(_0261_));
 sky130_fd_sc_hd__a21oi_4 _3136_ (.A1(net192),
    .A2(_1278_),
    .B1(_1318_),
    .Y(_0262_));
 sky130_fd_sc_hd__a21oi_4 _3137_ (.A1(net191),
    .A2(net130),
    .B1(net118),
    .Y(_0263_));
 sky130_fd_sc_hd__o21a_1 _3138_ (.A1(_0262_),
    .A2(_0263_),
    .B1(net34),
    .X(_0264_));
 sky130_fd_sc_hd__or4_1 _3139_ (.A(_0257_),
    .B(_0259_),
    .C(_0261_),
    .D(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__or4_1 _3140_ (.A(_0252_),
    .B(_0253_),
    .C(_0254_),
    .D(_0265_),
    .X(_0267_));
 sky130_fd_sc_hd__or3_1 _3141_ (.A(_0246_),
    .B(_0251_),
    .C(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__or4_1 _3142_ (.A(net71),
    .B(_1537_),
    .C(_1635_),
    .D(net16),
    .X(_0269_));
 sky130_fd_sc_hd__a2111o_1 _3143_ (.A1(net112),
    .A2(net144),
    .B1(_1357_),
    .C1(_1377_),
    .D1(net70),
    .X(_0270_));
 sky130_fd_sc_hd__or4_1 _3144_ (.A(_1243_),
    .B(_1325_),
    .C(_1654_),
    .D(_0270_),
    .X(_0271_));
 sky130_fd_sc_hd__o21a_1 _3145_ (.A1(_0269_),
    .A2(_0271_),
    .B1(net18),
    .X(_0272_));
 sky130_fd_sc_hd__o31a_2 _3146_ (.A1(_1367_),
    .A2(_1488_),
    .A3(_0058_),
    .B1(net17),
    .X(_0273_));
 sky130_fd_sc_hd__o21a_1 _3147_ (.A1(_1641_),
    .A2(_1689_),
    .B1(_1483_),
    .X(_0274_));
 sky130_fd_sc_hd__a22o_1 _3148_ (.A1(net182),
    .A2(net88),
    .B1(net151),
    .B2(net105),
    .X(_0275_));
 sky130_fd_sc_hd__or4_1 _3149_ (.A(_1390_),
    .B(_1744_),
    .C(_1754_),
    .D(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__or4_1 _3150_ (.A(_1324_),
    .B(net82),
    .C(_1368_),
    .D(_1488_),
    .X(_0278_));
 sky130_fd_sc_hd__o31a_4 _3151_ (.A1(_1872_),
    .A2(_0276_),
    .A3(_0278_),
    .B1(net24),
    .X(_0279_));
 sky130_fd_sc_hd__a21oi_4 _3152_ (.A1(net114),
    .A2(_1307_),
    .B1(net85),
    .Y(_0280_));
 sky130_fd_sc_hd__or4_1 _3153_ (.A(_1467_),
    .B(_1627_),
    .C(_0108_),
    .D(_0280_),
    .X(_0281_));
 sky130_fd_sc_hd__or4_1 _3154_ (.A(_1222_),
    .B(_1457_),
    .C(_1486_),
    .D(_1763_),
    .X(_0282_));
 sky130_fd_sc_hd__or3_1 _3155_ (.A(_1290_),
    .B(_1432_),
    .C(_1936_),
    .X(_0283_));
 sky130_fd_sc_hd__or3_1 _3156_ (.A(_0281_),
    .B(_0282_),
    .C(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__a21o_1 _3157_ (.A1(net53),
    .A2(_0284_),
    .B1(_0279_),
    .X(_0285_));
 sky130_fd_sc_hd__or4_1 _3158_ (.A(_0272_),
    .B(_0273_),
    .C(_0274_),
    .D(_0285_),
    .X(_0286_));
 sky130_fd_sc_hd__a21o_4 _3159_ (.A1(net119),
    .A2(net196),
    .B1(_1700_),
    .X(_0287_));
 sky130_fd_sc_hd__o21a_1 _3160_ (.A1(_1730_),
    .A2(_1923_),
    .B1(net61),
    .X(_0289_));
 sky130_fd_sc_hd__o31a_2 _3161_ (.A1(_1373_),
    .A2(net28),
    .A3(_1894_),
    .B1(net57),
    .X(_0290_));
 sky130_fd_sc_hd__o41a_1 _3162_ (.A1(_1391_),
    .A2(_1440_),
    .A3(_1446_),
    .A4(_1589_),
    .B1(net65),
    .X(_0291_));
 sky130_fd_sc_hd__a2111o_1 _3163_ (.A1(net50),
    .A2(_0287_),
    .B1(_0289_),
    .C1(_0290_),
    .D1(_0291_),
    .X(_0292_));
 sky130_fd_sc_hd__a21o_1 _3164_ (.A1(net183),
    .A2(net90),
    .B1(_2016_),
    .X(_0293_));
 sky130_fd_sc_hd__or2_4 _3165_ (.A(_1432_),
    .B(_1435_),
    .X(_0294_));
 sky130_fd_sc_hd__or4_4 _3166_ (.A(_1614_),
    .B(_2007_),
    .C(_0293_),
    .D(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__a211o_1 _3167_ (.A1(net112),
    .A2(net155),
    .B1(_1417_),
    .C1(_1867_),
    .X(_0296_));
 sky130_fd_sc_hd__or3_2 _3168_ (.A(_1654_),
    .B(_1660_),
    .C(_0296_),
    .X(_0297_));
 sky130_fd_sc_hd__a22o_1 _3169_ (.A1(net33),
    .A2(_0295_),
    .B1(_0297_),
    .B2(net41),
    .X(_0298_));
 sky130_fd_sc_hd__o21a_2 _3170_ (.A1(_1376_),
    .A2(_1753_),
    .B1(net17),
    .X(_0300_));
 sky130_fd_sc_hd__o21a_1 _3171_ (.A1(_1599_),
    .A2(_1606_),
    .B1(net49),
    .X(_0301_));
 sky130_fd_sc_hd__or4_1 _3172_ (.A(_0292_),
    .B(_0298_),
    .C(_0300_),
    .D(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__a21o_2 _3173_ (.A1(_1272_),
    .A2(net135),
    .B1(_1414_),
    .X(_0303_));
 sky130_fd_sc_hd__o31a_2 _3174_ (.A1(_1274_),
    .A2(_1498_),
    .A3(_0303_),
    .B1(net37),
    .X(_0304_));
 sky130_fd_sc_hd__or2_1 _3175_ (.A(_1460_),
    .B(net68),
    .X(_0305_));
 sky130_fd_sc_hd__o31a_1 _3176_ (.A1(_1323_),
    .A2(_1341_),
    .A3(_1581_),
    .B1(net35),
    .X(_0306_));
 sky130_fd_sc_hd__a21o_1 _3177_ (.A1(net41),
    .A2(_0305_),
    .B1(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__o41a_2 _3178_ (.A1(_1397_),
    .A2(_1596_),
    .A3(_1677_),
    .A4(_1763_),
    .B1(net40),
    .X(_0308_));
 sky130_fd_sc_hd__o21a_4 _3179_ (.A1(net197),
    .A2(net169),
    .B1(_1340_),
    .X(_0309_));
 sky130_fd_sc_hd__or3_2 _3180_ (.A(_1435_),
    .B(_1660_),
    .C(_0243_),
    .X(_0311_));
 sky130_fd_sc_hd__o21a_1 _3181_ (.A1(_0309_),
    .A2(_0311_),
    .B1(net45),
    .X(_0312_));
 sky130_fd_sc_hd__o41a_4 _3182_ (.A1(_1350_),
    .A2(_1646_),
    .A3(_1652_),
    .A4(_1687_),
    .B1(net22),
    .X(_0313_));
 sky130_fd_sc_hd__a2111o_1 _3183_ (.A1(net38),
    .A2(_1695_),
    .B1(_0308_),
    .C1(_0312_),
    .D1(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__a2111o_1 _3184_ (.A1(net57),
    .A2(_1565_),
    .B1(_0304_),
    .C1(_0307_),
    .D1(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__or4_2 _3185_ (.A(_0268_),
    .B(_0286_),
    .C(_0302_),
    .D(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__a22o_1 _3186_ (.A1(_1377_),
    .A2(net30),
    .B1(_1988_),
    .B2(net53),
    .X(_0317_));
 sky130_fd_sc_hd__a21oi_1 _3187_ (.A1(net62),
    .A2(_1920_),
    .B1(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__o21a_1 _3188_ (.A1(_1432_),
    .A2(_1763_),
    .B1(net53),
    .X(_0319_));
 sky130_fd_sc_hd__or4_1 _3189_ (.A(_0239_),
    .B(_0240_),
    .C(_0241_),
    .D(_0273_),
    .X(_0320_));
 sky130_fd_sc_hd__or4_1 _3190_ (.A(_0247_),
    .B(_0249_),
    .C(_0250_),
    .D(_0319_),
    .X(_0322_));
 sky130_fd_sc_hd__a221o_1 _3191_ (.A1(net33),
    .A2(_0295_),
    .B1(_0297_),
    .B2(net41),
    .C1(_0257_),
    .X(_0323_));
 sky130_fd_sc_hd__or4_1 _3192_ (.A(_0245_),
    .B(_0320_),
    .C(_0322_),
    .D(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__or4_1 _3193_ (.A(_1222_),
    .B(_1290_),
    .C(_1457_),
    .D(_1486_),
    .X(_0325_));
 sky130_fd_sc_hd__or4_1 _3194_ (.A(_1467_),
    .B(_1627_),
    .C(_1936_),
    .D(_0280_),
    .X(_0326_));
 sky130_fd_sc_hd__o31a_1 _3195_ (.A1(_0108_),
    .A2(_0325_),
    .A3(_0326_),
    .B1(net53),
    .X(_0327_));
 sky130_fd_sc_hd__a221o_1 _3196_ (.A1(net33),
    .A2(_0248_),
    .B1(_0287_),
    .B2(net50),
    .C1(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__or2_1 _3197_ (.A(_1391_),
    .B(_1440_),
    .X(_0329_));
 sky130_fd_sc_hd__o21a_1 _3198_ (.A1(_1446_),
    .A2(_1589_),
    .B1(net66),
    .X(_0330_));
 sky130_fd_sc_hd__a2111o_1 _3199_ (.A1(net65),
    .A2(_0329_),
    .B1(_0330_),
    .C1(_0274_),
    .D1(_0300_),
    .X(_0331_));
 sky130_fd_sc_hd__or4_1 _3200_ (.A(_0290_),
    .B(_0301_),
    .C(_0308_),
    .D(_0331_),
    .X(_0333_));
 sky130_fd_sc_hd__nor4_2 _3201_ (.A(_0289_),
    .B(_0324_),
    .C(_0328_),
    .D(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__a2111o_1 _3202_ (.A1(net38),
    .A2(_1695_),
    .B1(_0252_),
    .C1(_0304_),
    .D1(_0306_),
    .X(_0335_));
 sky130_fd_sc_hd__or4_1 _3203_ (.A(_0253_),
    .B(_0272_),
    .C(_0279_),
    .D(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__o21a_1 _3204_ (.A1(_1267_),
    .A2(_1322_),
    .B1(net38),
    .X(_0337_));
 sky130_fd_sc_hd__a211o_1 _3205_ (.A1(net45),
    .A2(_0309_),
    .B1(_0313_),
    .C1(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__a221o_1 _3206_ (.A1(net38),
    .A2(_0258_),
    .B1(_0311_),
    .B2(net45),
    .C1(_0261_),
    .X(_0339_));
 sky130_fd_sc_hd__a21o_1 _3207_ (.A1(net41),
    .A2(_0305_),
    .B1(_0264_),
    .X(_0340_));
 sky130_fd_sc_hd__a2111o_1 _3208_ (.A1(net58),
    .A2(_1565_),
    .B1(_0254_),
    .C1(_0339_),
    .D1(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__nor3_1 _3209_ (.A(_0336_),
    .B(_0338_),
    .C(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__and4_1 _3210_ (.A(_0227_),
    .B(_0318_),
    .C(_0334_),
    .D(_0342_),
    .X(_0344_));
 sky130_fd_sc_hd__or4b_1 _3211_ (.A(_1780_),
    .B(_1880_),
    .C(_1906_),
    .D_N(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__or3_2 _3212_ (.A(_1425_),
    .B(_1440_),
    .C(_1446_),
    .X(_0346_));
 sky130_fd_sc_hd__or3_1 _3213_ (.A(_1268_),
    .B(_1315_),
    .C(_1331_),
    .X(_0347_));
 sky130_fd_sc_hd__a221o_4 _3214_ (.A1(net30),
    .A2(_0346_),
    .B1(_0347_),
    .B2(net46),
    .C1(_0233_),
    .X(_0348_));
 sky130_fd_sc_hd__or4_1 _3215_ (.A(_0093_),
    .B(_0234_),
    .C(_0345_),
    .D(_0348_),
    .X(_0049_));
 sky130_fd_sc_hd__o2111a_2 _3216_ (.A1(net189),
    .A2(_1277_),
    .B1(net163),
    .C1(net238),
    .D1(net263),
    .X(_0349_));
 sky130_fd_sc_hd__o41a_4 _3217_ (.A1(_1257_),
    .A2(_1442_),
    .A3(_1711_),
    .A4(_0349_),
    .B1(net55),
    .X(_0350_));
 sky130_fd_sc_hd__o41a_1 _3218_ (.A1(_1362_),
    .A2(_1373_),
    .A3(net27),
    .A4(_1795_),
    .B1(net64),
    .X(_0351_));
 sky130_fd_sc_hd__a21o_1 _3219_ (.A1(net195),
    .A2(net84),
    .B1(_1432_),
    .X(_0352_));
 sky130_fd_sc_hd__or3_1 _3220_ (.A(_1469_),
    .B(_1526_),
    .C(_0210_),
    .X(_0354_));
 sky130_fd_sc_hd__or4_1 _3221_ (.A(_1354_),
    .B(_1391_),
    .C(net76),
    .D(net68),
    .X(_0355_));
 sky130_fd_sc_hd__o41a_1 _3222_ (.A1(_1376_),
    .A2(_1467_),
    .A3(_1629_),
    .A4(_0355_),
    .B1(net29),
    .X(_0356_));
 sky130_fd_sc_hd__a211o_1 _3223_ (.A1(_1288_),
    .A2(net145),
    .B1(_1479_),
    .C1(_1486_),
    .X(_0357_));
 sky130_fd_sc_hd__or2_1 _3224_ (.A(_1526_),
    .B(_1795_),
    .X(_0358_));
 sky130_fd_sc_hd__and3_2 _3225_ (.A(net267),
    .B(_1121_),
    .C(_1408_),
    .X(_0359_));
 sky130_fd_sc_hd__a21o_1 _3226_ (.A1(net123),
    .A2(net151),
    .B1(_1365_),
    .X(_0360_));
 sky130_fd_sc_hd__o21a_2 _3227_ (.A1(_1315_),
    .A2(_1539_),
    .B1(net56),
    .X(_0361_));
 sky130_fd_sc_hd__or4_4 _3228_ (.A(_1309_),
    .B(net71),
    .C(_1529_),
    .D(_1626_),
    .X(_0362_));
 sky130_fd_sc_hd__a22o_2 _3229_ (.A1(net202),
    .A2(net105),
    .B1(net88),
    .B2(net242),
    .X(_0363_));
 sky130_fd_sc_hd__or4_1 _3230_ (.A(_1727_),
    .B(_1934_),
    .C(_1992_),
    .D(_0363_),
    .X(_0365_));
 sky130_fd_sc_hd__a22o_4 _3231_ (.A1(net181),
    .A2(net98),
    .B1(net140),
    .B2(_1089_),
    .X(_0366_));
 sky130_fd_sc_hd__or4_1 _3232_ (.A(_0979_),
    .B(_1589_),
    .C(_1939_),
    .D(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__or4_1 _3233_ (.A(_1484_),
    .B(_1578_),
    .C(_1951_),
    .D(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__or4_1 _3234_ (.A(_1243_),
    .B(net94),
    .C(_1489_),
    .D(_1518_),
    .X(_0369_));
 sky130_fd_sc_hd__or2_2 _3235_ (.A(_1324_),
    .B(_1347_),
    .X(_0370_));
 sky130_fd_sc_hd__or4_1 _3236_ (.A(_1421_),
    .B(_1538_),
    .C(_1596_),
    .D(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__o21a_1 _3237_ (.A1(_0369_),
    .A2(_0371_),
    .B1(net44),
    .X(_0372_));
 sky130_fd_sc_hd__a21oi_4 _3238_ (.A1(net199),
    .A2(net137),
    .B1(net79),
    .Y(_0373_));
 sky130_fd_sc_hd__a21o_1 _3239_ (.A1(net172),
    .A2(net81),
    .B1(_1363_),
    .X(_0374_));
 sky130_fd_sc_hd__a21oi_1 _3240_ (.A1(net241),
    .A2(net115),
    .B1(net121),
    .Y(_0376_));
 sky130_fd_sc_hd__a22o_1 _3241_ (.A1(net124),
    .A2(net180),
    .B1(net179),
    .B2(net88),
    .X(_0377_));
 sky130_fd_sc_hd__o41a_1 _3242_ (.A1(_1509_),
    .A2(_1516_),
    .A3(_1575_),
    .A4(_0377_),
    .B1(net57),
    .X(_0378_));
 sky130_fd_sc_hd__o31a_2 _3243_ (.A1(_1357_),
    .A2(_1552_),
    .A3(_0359_),
    .B1(net40),
    .X(_0379_));
 sky130_fd_sc_hd__o21a_1 _3244_ (.A1(_1510_),
    .A2(_1556_),
    .B1(net48),
    .X(_0380_));
 sky130_fd_sc_hd__a22o_1 _3245_ (.A1(net22),
    .A2(_1606_),
    .B1(_1972_),
    .B2(net30),
    .X(_0381_));
 sky130_fd_sc_hd__a211o_1 _3246_ (.A1(net173),
    .A2(net81),
    .B1(_1394_),
    .C1(_1363_),
    .X(_0382_));
 sky130_fd_sc_hd__o41a_1 _3247_ (.A1(_1639_),
    .A2(_1920_),
    .A3(_0373_),
    .A4(_0382_),
    .B1(net17),
    .X(_0383_));
 sky130_fd_sc_hd__or4_1 _3248_ (.A(_0350_),
    .B(_0356_),
    .C(_0378_),
    .D(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__o31a_1 _3249_ (.A1(_1397_),
    .A2(_1795_),
    .A3(_0376_),
    .B1(net19),
    .X(_0385_));
 sky130_fd_sc_hd__or4_1 _3250_ (.A(_1700_),
    .B(_1811_),
    .C(_0352_),
    .D(_0358_),
    .X(_0387_));
 sky130_fd_sc_hd__or3_1 _3251_ (.A(_1362_),
    .B(_1363_),
    .C(_1931_),
    .X(_0388_));
 sky130_fd_sc_hd__or3_1 _3252_ (.A(_1555_),
    .B(_1827_),
    .C(_1962_),
    .X(_0389_));
 sky130_fd_sc_hd__o31a_1 _3253_ (.A1(_0387_),
    .A2(_0388_),
    .A3(_0389_),
    .B1(net39),
    .X(_0390_));
 sky130_fd_sc_hd__or2_2 _3254_ (.A(_1434_),
    .B(_0360_),
    .X(_0391_));
 sky130_fd_sc_hd__or4_1 _3255_ (.A(_1464_),
    .B(_1526_),
    .C(_1802_),
    .D(_1923_),
    .X(_0392_));
 sky130_fd_sc_hd__a221o_1 _3256_ (.A1(net42),
    .A2(_0365_),
    .B1(_0368_),
    .B2(net35),
    .C1(_0372_),
    .X(_0393_));
 sky130_fd_sc_hd__a221o_1 _3257_ (.A1(net64),
    .A2(_0352_),
    .B1(_0392_),
    .B2(net17),
    .C1(_0361_),
    .X(_0394_));
 sky130_fd_sc_hd__a2111o_1 _3258_ (.A1(net123),
    .A2(net195),
    .B1(net73),
    .C1(_1699_),
    .D1(_1915_),
    .X(_0395_));
 sky130_fd_sc_hd__a22o_1 _3259_ (.A1(_1292_),
    .A2(net42),
    .B1(net36),
    .B2(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__a221o_1 _3260_ (.A1(net65),
    .A2(_0354_),
    .B1(_0391_),
    .B2(net48),
    .C1(_0396_),
    .X(_0398_));
 sky130_fd_sc_hd__a211o_1 _3261_ (.A1(net24),
    .A2(_0357_),
    .B1(_0380_),
    .C1(_0381_),
    .X(_0399_));
 sky130_fd_sc_hd__or4_1 _3262_ (.A(_1257_),
    .B(_1376_),
    .C(_1377_),
    .D(_1851_),
    .X(_0400_));
 sky130_fd_sc_hd__o41a_1 _3263_ (.A1(_1222_),
    .A2(_1509_),
    .A3(_0362_),
    .A4(_0400_),
    .B1(net36),
    .X(_0401_));
 sky130_fd_sc_hd__or4_1 _3264_ (.A(_0394_),
    .B(_0398_),
    .C(_0399_),
    .D(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__or4_1 _3265_ (.A(_1517_),
    .B(_1881_),
    .C(_1983_),
    .D(_2017_),
    .X(_0403_));
 sky130_fd_sc_hd__o31a_1 _3266_ (.A1(_1488_),
    .A2(_1565_),
    .A3(_0403_),
    .B1(net32),
    .X(_0404_));
 sky130_fd_sc_hd__or3_1 _3267_ (.A(_1319_),
    .B(net82),
    .C(_1577_),
    .X(_0405_));
 sky130_fd_sc_hd__a22o_1 _3268_ (.A1(net63),
    .A2(_1533_),
    .B1(_0405_),
    .B2(net32),
    .X(_0406_));
 sky130_fd_sc_hd__a2111o_1 _3269_ (.A1(net21),
    .A2(_0085_),
    .B1(_0379_),
    .C1(_0385_),
    .D1(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__or4_1 _3270_ (.A(_0351_),
    .B(_0384_),
    .C(_0404_),
    .D(_0407_),
    .X(_0409_));
 sky130_fd_sc_hd__or4_4 _3271_ (.A(_0390_),
    .B(_0393_),
    .C(_0402_),
    .D(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__or2_1 _3272_ (.A(_1500_),
    .B(_1654_),
    .X(_0411_));
 sky130_fd_sc_hd__o41a_1 _3273_ (.A1(_1405_),
    .A2(_1469_),
    .A3(_1557_),
    .A4(net70),
    .B1(net40),
    .X(_0412_));
 sky130_fd_sc_hd__a21oi_1 _3274_ (.A1(net43),
    .A2(_0411_),
    .B1(_0412_),
    .Y(_0413_));
 sky130_fd_sc_hd__nand2_1 _3275_ (.A(_0076_),
    .B(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__or4_1 _3276_ (.A(_0068_),
    .B(_0073_),
    .C(_0158_),
    .D(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__or4_1 _3277_ (.A(_0231_),
    .B(_0345_),
    .C(_0410_),
    .D(_0415_),
    .X(_0050_));
 sky130_fd_sc_hd__or4_4 _3278_ (.A(_1700_),
    .B(_1701_),
    .C(_1707_),
    .D(_1709_),
    .X(_0416_));
 sky130_fd_sc_hd__or2_1 _3279_ (.A(_1540_),
    .B(_1753_),
    .X(_0417_));
 sky130_fd_sc_hd__a22o_1 _3280_ (.A1(_1012_),
    .A2(net184),
    .B1(net98),
    .B2(net211),
    .X(_0419_));
 sky130_fd_sc_hd__or3_1 _3281_ (.A(_1447_),
    .B(_0416_),
    .C(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__o41a_4 _3282_ (.A1(net178),
    .A2(net168),
    .A3(net140),
    .A4(net134),
    .B1(net89),
    .X(_0421_));
 sky130_fd_sc_hd__a21oi_2 _3283_ (.A1(net199),
    .A2(net190),
    .B1(net86),
    .Y(_0422_));
 sky130_fd_sc_hd__or4_1 _3284_ (.A(_1453_),
    .B(_1734_),
    .C(_0077_),
    .D(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__or3_2 _3285_ (.A(_1310_),
    .B(_0421_),
    .C(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__a21oi_4 _3286_ (.A1(net113),
    .A2(net148),
    .B1(net109),
    .Y(_0425_));
 sky130_fd_sc_hd__or3_1 _3287_ (.A(_1509_),
    .B(_1629_),
    .C(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__or2_1 _3288_ (.A(_1638_),
    .B(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__or2_2 _3289_ (.A(_1527_),
    .B(_1936_),
    .X(_0428_));
 sky130_fd_sc_hd__or3_2 _3290_ (.A(_1460_),
    .B(_1644_),
    .C(_1653_),
    .X(_0430_));
 sky130_fd_sc_hd__or4_4 _3291_ (.A(net72),
    .B(net71),
    .C(_1537_),
    .D(_1699_),
    .X(_0431_));
 sky130_fd_sc_hd__or2_2 _3292_ (.A(_1406_),
    .B(_1424_),
    .X(_0432_));
 sky130_fd_sc_hd__a41oi_4 _3293_ (.A1(net114),
    .A2(net93),
    .A3(net148),
    .A4(net142),
    .B1(_1404_),
    .Y(_0433_));
 sky130_fd_sc_hd__or2_1 _3294_ (.A(net74),
    .B(_1569_),
    .X(_0434_));
 sky130_fd_sc_hd__o2111a_4 _3295_ (.A1(net204),
    .A2(net194),
    .B1(net164),
    .C1(net238),
    .D1(net252),
    .X(_0435_));
 sky130_fd_sc_hd__or3_1 _3296_ (.A(net74),
    .B(net70),
    .C(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__or2_1 _3297_ (.A(_0433_),
    .B(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__o41a_1 _3298_ (.A1(net243),
    .A2(net204),
    .A3(net194),
    .A4(net189),
    .B1(_1205_),
    .X(_0438_));
 sky130_fd_sc_hd__or3_1 _3299_ (.A(_1688_),
    .B(_1711_),
    .C(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__or4_4 _3300_ (.A(_1508_),
    .B(net27),
    .C(_1695_),
    .D(_1697_),
    .X(_0441_));
 sky130_fd_sc_hd__o41a_2 _3301_ (.A1(net243),
    .A2(net204),
    .A3(net195),
    .A4(_1230_),
    .B1(net125),
    .X(_0442_));
 sky130_fd_sc_hd__or4_1 _3302_ (.A(_1564_),
    .B(_1750_),
    .C(_1754_),
    .D(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__or2_4 _3303_ (.A(_1529_),
    .B(_1868_),
    .X(_0444_));
 sky130_fd_sc_hd__a21oi_4 _3304_ (.A1(net149),
    .A2(net143),
    .B1(net117),
    .Y(_0445_));
 sky130_fd_sc_hd__or2_2 _3305_ (.A(_1459_),
    .B(_1480_),
    .X(_0446_));
 sky130_fd_sc_hd__or2_4 _3306_ (.A(_1722_),
    .B(net69),
    .X(_0447_));
 sky130_fd_sc_hd__or4_2 _3307_ (.A(_1292_),
    .B(_1297_),
    .C(_1768_),
    .D(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__or2_4 _3308_ (.A(_1478_),
    .B(_1781_),
    .X(_0449_));
 sky130_fd_sc_hd__a21oi_4 _3309_ (.A1(net199),
    .A2(net166),
    .B1(net117),
    .Y(_0450_));
 sky130_fd_sc_hd__or4_1 _3310_ (.A(_1717_),
    .B(_1926_),
    .C(_0449_),
    .D(_0450_),
    .X(_0452_));
 sky130_fd_sc_hd__or2_4 _3311_ (.A(_1792_),
    .B(_2016_),
    .X(_0453_));
 sky130_fd_sc_hd__a21oi_4 _3312_ (.A1(net240),
    .A2(net185),
    .B1(net97),
    .Y(_0454_));
 sky130_fd_sc_hd__or4_1 _3313_ (.A(_0430_),
    .B(_0431_),
    .C(_0439_),
    .D(_0452_),
    .X(_0455_));
 sky130_fd_sc_hd__or4_1 _3314_ (.A(_1419_),
    .B(_1471_),
    .C(_1628_),
    .D(_1731_),
    .X(_0456_));
 sky130_fd_sc_hd__or3_1 _3315_ (.A(_0444_),
    .B(_0446_),
    .C(_0453_),
    .X(_0457_));
 sky130_fd_sc_hd__or4b_1 _3316_ (.A(_1421_),
    .B(_1583_),
    .C(_1439_),
    .D_N(_1524_),
    .X(_0458_));
 sky130_fd_sc_hd__or3_2 _3317_ (.A(_0456_),
    .B(_0457_),
    .C(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__or4_1 _3318_ (.A(_0420_),
    .B(_0424_),
    .C(_0455_),
    .D(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__or3_1 _3319_ (.A(_0441_),
    .B(_0445_),
    .C(_0448_),
    .X(_0461_));
 sky130_fd_sc_hd__or2_1 _3320_ (.A(_0107_),
    .B(_0454_),
    .X(_0463_));
 sky130_fd_sc_hd__or3_2 _3321_ (.A(_1454_),
    .B(_1550_),
    .C(_0428_),
    .X(_0464_));
 sky130_fd_sc_hd__or4b_1 _3322_ (.A(_1650_),
    .B(_1803_),
    .C(_1812_),
    .D_N(_0087_),
    .X(_0465_));
 sky130_fd_sc_hd__or4_1 _3323_ (.A(_0437_),
    .B(_0463_),
    .C(_0464_),
    .D(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__or4_1 _3324_ (.A(_0427_),
    .B(_0443_),
    .C(_0461_),
    .D(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__or3_1 _3325_ (.A(_1695_),
    .B(_1696_),
    .C(_0445_),
    .X(_0468_));
 sky130_fd_sc_hd__o21a_1 _3326_ (.A1(_0460_),
    .A2(_0467_),
    .B1(net35),
    .X(_0469_));
 sky130_fd_sc_hd__a21oi_4 _3327_ (.A1(net106),
    .A2(net100),
    .B1(net97),
    .Y(_0470_));
 sky130_fd_sc_hd__or4_2 _3328_ (.A(_1671_),
    .B(_1760_),
    .C(_0454_),
    .D(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__or3_2 _3329_ (.A(_1568_),
    .B(_1890_),
    .C(_1936_),
    .X(_0472_));
 sky130_fd_sc_hd__a21oi_4 _3330_ (.A1(net206),
    .A2(net175),
    .B1(_1359_),
    .Y(_0474_));
 sky130_fd_sc_hd__or2_2 _3331_ (.A(_1682_),
    .B(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__or4_2 _3332_ (.A(net71),
    .B(_1529_),
    .C(_1792_),
    .D(net68),
    .X(_0476_));
 sky130_fd_sc_hd__or4_2 _3333_ (.A(_0436_),
    .B(_0472_),
    .C(_0475_),
    .D(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__or3_4 _3334_ (.A(net82),
    .B(_1331_),
    .C(_1885_),
    .X(_0478_));
 sky130_fd_sc_hd__or4_4 _3335_ (.A(_1163_),
    .B(_1595_),
    .C(_1881_),
    .D(_0478_),
    .X(_0479_));
 sky130_fd_sc_hd__o2111a_2 _3336_ (.A1(net204),
    .A2(net168),
    .B1(net252),
    .C1(net228),
    .D1(net220),
    .X(_0480_));
 sky130_fd_sc_hd__or3_2 _3337_ (.A(_1494_),
    .B(_1495_),
    .C(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__or4_2 _3338_ (.A(_1601_),
    .B(_1619_),
    .C(_0479_),
    .D(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__or3_2 _3339_ (.A(_1707_),
    .B(_1709_),
    .C(_0349_),
    .X(_0483_));
 sky130_fd_sc_hd__or3_1 _3340_ (.A(_1291_),
    .B(_1391_),
    .C(_1767_),
    .X(_0485_));
 sky130_fd_sc_hd__or4_1 _3341_ (.A(net72),
    .B(_1537_),
    .C(_1699_),
    .D(_1700_),
    .X(_0486_));
 sky130_fd_sc_hd__or4_2 _3342_ (.A(net75),
    .B(_1811_),
    .C(_0449_),
    .D(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__or3_1 _3343_ (.A(_0483_),
    .B(_0485_),
    .C(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__or4_1 _3344_ (.A(_0471_),
    .B(_0477_),
    .C(_0482_),
    .D(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__or4_1 _3345_ (.A(_1305_),
    .B(_1642_),
    .C(_1723_),
    .D(_1734_),
    .X(_0490_));
 sky130_fd_sc_hd__a21o_1 _3346_ (.A1(net125),
    .A2(net198),
    .B1(_1431_),
    .X(_0491_));
 sky130_fd_sc_hd__or4_4 _3347_ (.A(_1369_),
    .B(_1447_),
    .C(_1453_),
    .D(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__a21oi_4 _3348_ (.A1(net240),
    .A2(net143),
    .B1(net104),
    .Y(_0493_));
 sky130_fd_sc_hd__or2_4 _3349_ (.A(_1390_),
    .B(_1802_),
    .X(_0494_));
 sky130_fd_sc_hd__and3_2 _3350_ (.A(_0682_),
    .B(net270),
    .C(_1252_),
    .X(_0496_));
 sky130_fd_sc_hd__and3_2 _3351_ (.A(_0682_),
    .B(net267),
    .C(net125),
    .X(_0497_));
 sky130_fd_sc_hd__or4_1 _3352_ (.A(_0493_),
    .B(_0494_),
    .C(_0496_),
    .D(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__or2_4 _3353_ (.A(_1851_),
    .B(net67),
    .X(_0499_));
 sky130_fd_sc_hd__or4_1 _3354_ (.A(_1670_),
    .B(_0294_),
    .C(_0373_),
    .D(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__or4_2 _3355_ (.A(_0490_),
    .B(_0492_),
    .C(_0498_),
    .D(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__a211o_2 _3356_ (.A1(_1288_),
    .A2(net146),
    .B1(_1644_),
    .C1(_1653_),
    .X(_0502_));
 sky130_fd_sc_hd__or3_1 _3357_ (.A(_1258_),
    .B(_1511_),
    .C(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__o31a_2 _3358_ (.A1(net178),
    .A2(net140),
    .A3(net134),
    .B1(net125),
    .X(_0504_));
 sky130_fd_sc_hd__nor2_4 _3359_ (.A(_1867_),
    .B(_1915_),
    .Y(_0505_));
 sky130_fd_sc_hd__or3b_1 _3360_ (.A(_1785_),
    .B(net13),
    .C_N(_0505_),
    .X(_0507_));
 sky130_fd_sc_hd__or4b_1 _3361_ (.A(_1785_),
    .B(net13),
    .C(_0504_),
    .D_N(_0505_),
    .X(_0508_));
 sky130_fd_sc_hd__and3_4 _3362_ (.A(net272),
    .B(net264),
    .C(net120),
    .X(_0509_));
 sky130_fd_sc_hd__or4_1 _3363_ (.A(_1366_),
    .B(_1374_),
    .C(_1460_),
    .D(_1606_),
    .X(_0510_));
 sky130_fd_sc_hd__or4_4 _3364_ (.A(_1535_),
    .B(_1753_),
    .C(_0509_),
    .D(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__or3_1 _3365_ (.A(_1382_),
    .B(_1383_),
    .C(_1766_),
    .X(_0512_));
 sky130_fd_sc_hd__or4_1 _3366_ (.A(_0503_),
    .B(_0508_),
    .C(_0511_),
    .D(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__o41a_2 _3367_ (.A1(net178),
    .A2(net168),
    .A3(net140),
    .A4(net135),
    .B1(_0913_),
    .X(_0514_));
 sky130_fd_sc_hd__a21oi_4 _3368_ (.A1(net240),
    .A2(net185),
    .B1(net128),
    .Y(_0515_));
 sky130_fd_sc_hd__or4_1 _3369_ (.A(_1589_),
    .B(_1590_),
    .C(_0514_),
    .D(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__a21oi_4 _3370_ (.A1(net240),
    .A2(net143),
    .B1(net117),
    .Y(_0518_));
 sky130_fd_sc_hd__or2_1 _3371_ (.A(_1731_),
    .B(_0445_),
    .X(_0519_));
 sky130_fd_sc_hd__or4_2 _3372_ (.A(_1731_),
    .B(_0263_),
    .C(_0445_),
    .D(_0450_),
    .X(_0520_));
 sky130_fd_sc_hd__a21oi_4 _3373_ (.A1(net113),
    .A2(net91),
    .B1(net128),
    .Y(_0521_));
 sky130_fd_sc_hd__o41a_1 _3374_ (.A1(_1146_),
    .A2(net155),
    .A3(net152),
    .A4(net146),
    .B1(_0913_),
    .X(_0522_));
 sky130_fd_sc_hd__or4_2 _3375_ (.A(_1034_),
    .B(_1678_),
    .C(_1679_),
    .D(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__or4_4 _3376_ (.A(_0441_),
    .B(_0516_),
    .C(_0520_),
    .D(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__a21oi_4 _3377_ (.A1(net206),
    .A2(net175),
    .B1(net79),
    .Y(_0525_));
 sky130_fd_sc_hd__or4_2 _3378_ (.A(_1628_),
    .B(_1630_),
    .C(_0422_),
    .D(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__o21a_4 _3379_ (.A1(net198),
    .A2(net152),
    .B1(_1340_),
    .X(_0527_));
 sky130_fd_sc_hd__a2111o_2 _3380_ (.A1(net198),
    .A2(_1340_),
    .B1(_1517_),
    .C1(_1565_),
    .D1(_1763_),
    .X(_0529_));
 sky130_fd_sc_hd__or3_4 _3381_ (.A(_1490_),
    .B(_1579_),
    .C(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__or3_1 _3382_ (.A(_0439_),
    .B(_0526_),
    .C(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__or4_1 _3383_ (.A(_0501_),
    .B(_0513_),
    .C(_0524_),
    .D(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__o21a_1 _3384_ (.A1(_0489_),
    .A2(_0532_),
    .B1(net43),
    .X(_0533_));
 sky130_fd_sc_hd__or3_2 _3385_ (.A(_1590_),
    .B(_1591_),
    .C(_0515_),
    .X(_0534_));
 sky130_fd_sc_hd__or3b_1 _3386_ (.A(_1420_),
    .B(_1651_),
    .C_N(_1659_),
    .X(_0535_));
 sky130_fd_sc_hd__or3_1 _3387_ (.A(_0475_),
    .B(_0534_),
    .C(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__or2_4 _3388_ (.A(_1368_),
    .B(_1397_),
    .X(_0537_));
 sky130_fd_sc_hd__or3_1 _3389_ (.A(_1677_),
    .B(_1679_),
    .C(_0537_),
    .X(_0538_));
 sky130_fd_sc_hd__or2_2 _3390_ (.A(_1382_),
    .B(_0494_),
    .X(_0540_));
 sky130_fd_sc_hd__or2_1 _3391_ (.A(_1491_),
    .B(_1658_),
    .X(_0541_));
 sky130_fd_sc_hd__or4_2 _3392_ (.A(_1757_),
    .B(_0538_),
    .C(_0540_),
    .D(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__or3_1 _3393_ (.A(_1343_),
    .B(_1367_),
    .C(_1548_),
    .X(_0543_));
 sky130_fd_sc_hd__o2111a_4 _3394_ (.A1(net184),
    .A2(net155),
    .B1(net252),
    .C1(net238),
    .D1(net220),
    .X(_0544_));
 sky130_fd_sc_hd__or3_1 _3395_ (.A(_1607_),
    .B(_0543_),
    .C(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__or4_1 _3396_ (.A(_1519_),
    .B(_0502_),
    .C(_0527_),
    .D(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__or4_1 _3397_ (.A(_0482_),
    .B(_0536_),
    .C(_0542_),
    .D(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__a22o_1 _3398_ (.A1(net211),
    .A2(net125),
    .B1(_1252_),
    .B2(net181),
    .X(_0548_));
 sky130_fd_sc_hd__a21o_1 _3399_ (.A1(net112),
    .A2(net152),
    .B1(_1365_),
    .X(_0549_));
 sky130_fd_sc_hd__a21o_1 _3400_ (.A1(net194),
    .A2(net89),
    .B1(_1480_),
    .X(_0551_));
 sky130_fd_sc_hd__or4_1 _3401_ (.A(_0085_),
    .B(_0548_),
    .C(_0549_),
    .D(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__or4_1 _3402_ (.A(_1268_),
    .B(_1275_),
    .C(_1378_),
    .D(_1379_),
    .X(_0553_));
 sky130_fd_sc_hd__or4_1 _3403_ (.A(_1647_),
    .B(_1702_),
    .C(_1829_),
    .D(_1940_),
    .X(_0554_));
 sky130_fd_sc_hd__or4_1 _3404_ (.A(_1415_),
    .B(_1530_),
    .C(_1625_),
    .D(_1764_),
    .X(_0555_));
 sky130_fd_sc_hd__or4_1 _3405_ (.A(_0552_),
    .B(_0553_),
    .C(_0554_),
    .D(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__or4_2 _3406_ (.A(_1488_),
    .B(_1578_),
    .C(_1650_),
    .D(_0260_),
    .X(_0557_));
 sky130_fd_sc_hd__or3_4 _3407_ (.A(net16),
    .B(_1765_),
    .C(net14),
    .X(_0558_));
 sky130_fd_sc_hd__a41o_1 _3408_ (.A1(net113),
    .A2(net91),
    .A3(net149),
    .A4(net143),
    .B1(net79),
    .X(_0559_));
 sky130_fd_sc_hd__or4b_1 _3409_ (.A(net16),
    .B(_1765_),
    .C(net14),
    .D_N(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__nand3_1 _3410_ (.A(_1698_),
    .B(_1737_),
    .C(_1738_),
    .Y(_0562_));
 sky130_fd_sc_hd__or3_1 _3411_ (.A(_1692_),
    .B(_1714_),
    .C(_1716_),
    .X(_0563_));
 sky130_fd_sc_hd__or4_4 _3412_ (.A(_0557_),
    .B(_0560_),
    .C(_0562_),
    .D(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__or2_1 _3413_ (.A(_1296_),
    .B(_1526_),
    .X(_0565_));
 sky130_fd_sc_hd__or4_2 _3414_ (.A(_1502_),
    .B(_1637_),
    .C(_0447_),
    .D(_0565_),
    .X(_0566_));
 sky130_fd_sc_hd__or3_1 _3415_ (.A(_1508_),
    .B(net28),
    .C(_1915_),
    .X(_0567_));
 sky130_fd_sc_hd__a21oi_4 _3416_ (.A1(net190),
    .A2(net185),
    .B1(net117),
    .Y(_0568_));
 sky130_fd_sc_hd__or3_1 _3417_ (.A(_0431_),
    .B(_0518_),
    .C(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__or3_1 _3418_ (.A(_0566_),
    .B(_0567_),
    .C(_0569_),
    .X(_0570_));
 sky130_fd_sc_hd__a21oi_4 _3419_ (.A1(net201),
    .A2(net165),
    .B1(_1389_),
    .Y(_0571_));
 sky130_fd_sc_hd__o211a_1 _3420_ (.A1(net204),
    .A2(net168),
    .B1(net163),
    .C1(net263),
    .X(_0573_));
 sky130_fd_sc_hd__or3_1 _3421_ (.A(_1610_),
    .B(_1792_),
    .C(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__or4_4 _3422_ (.A(_0275_),
    .B(_0374_),
    .C(_0376_),
    .D(_0450_),
    .X(_0575_));
 sky130_fd_sc_hd__or3_1 _3423_ (.A(_1545_),
    .B(_1589_),
    .C(_1598_),
    .X(_0576_));
 sky130_fd_sc_hd__a21oi_1 _3424_ (.A1(net206),
    .A2(net175),
    .B1(net128),
    .Y(_0577_));
 sky130_fd_sc_hd__or4_1 _3425_ (.A(_1545_),
    .B(_1589_),
    .C(_1598_),
    .D(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__or2_1 _3426_ (.A(_1425_),
    .B(_1455_),
    .X(_0579_));
 sky130_fd_sc_hd__or4_2 _3427_ (.A(_1425_),
    .B(_1455_),
    .C(_1755_),
    .D(_0435_),
    .X(_0580_));
 sky130_fd_sc_hd__or4_1 _3428_ (.A(_0574_),
    .B(_0575_),
    .C(_0578_),
    .D(_0580_),
    .X(_0581_));
 sky130_fd_sc_hd__or4_1 _3429_ (.A(_0556_),
    .B(_0564_),
    .C(_0570_),
    .D(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__or4_1 _3430_ (.A(_1343_),
    .B(_1519_),
    .C(_0527_),
    .D(_0544_),
    .X(_0584_));
 sky130_fd_sc_hd__o41a_1 _3431_ (.A1(net205),
    .A2(_1277_),
    .A3(_1326_),
    .A4(net135),
    .B1(_1089_),
    .X(_0585_));
 sky130_fd_sc_hd__or3_1 _3432_ (.A(_1367_),
    .B(_1548_),
    .C(_1607_),
    .X(_0586_));
 sky130_fd_sc_hd__o21a_1 _3433_ (.A1(_0547_),
    .A2(_0582_),
    .B1(_1427_),
    .X(_0587_));
 sky130_fd_sc_hd__or4_2 _3434_ (.A(_1717_),
    .B(_1926_),
    .C(_0449_),
    .D(_0585_),
    .X(_0588_));
 sky130_fd_sc_hd__or3_2 _3435_ (.A(_1034_),
    .B(_1679_),
    .C(_1716_),
    .X(_0589_));
 sky130_fd_sc_hd__or3_4 _3436_ (.A(_1291_),
    .B(_1767_),
    .C(_0480_),
    .X(_0590_));
 sky130_fd_sc_hd__or4_2 _3437_ (.A(_1529_),
    .B(_1544_),
    .C(_1600_),
    .D(_1915_),
    .X(_0591_));
 sky130_fd_sc_hd__or4_1 _3438_ (.A(_0534_),
    .B(_0589_),
    .C(_0590_),
    .D(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__or2_4 _3439_ (.A(_1506_),
    .B(_0084_),
    .X(_0593_));
 sky130_fd_sc_hd__or2_1 _3440_ (.A(_0453_),
    .B(_0593_),
    .X(_0595_));
 sky130_fd_sc_hd__or2_4 _3441_ (.A(_1625_),
    .B(_0425_),
    .X(_0596_));
 sky130_fd_sc_hd__or4_1 _3442_ (.A(_0102_),
    .B(_0161_),
    .C(_0595_),
    .D(_0596_),
    .X(_0597_));
 sky130_fd_sc_hd__or3_1 _3443_ (.A(_0588_),
    .B(_0592_),
    .C(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__or2_1 _3444_ (.A(_0085_),
    .B(_0504_),
    .X(_0599_));
 sky130_fd_sc_hd__or3_1 _3445_ (.A(_1379_),
    .B(_1559_),
    .C(_1681_),
    .X(_0600_));
 sky130_fd_sc_hd__or4_4 _3446_ (.A(net73),
    .B(net27),
    .C(_1697_),
    .D(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__or4_2 _3447_ (.A(_0479_),
    .B(_0569_),
    .C(_0599_),
    .D(_0601_),
    .X(_0602_));
 sky130_fd_sc_hd__or4_2 _3448_ (.A(_1320_),
    .B(_1434_),
    .C(_1599_),
    .D(_1606_),
    .X(_0603_));
 sky130_fd_sc_hd__or3_1 _3449_ (.A(_1438_),
    .B(_1443_),
    .C(_0175_),
    .X(_0604_));
 sky130_fd_sc_hd__or4_1 _3450_ (.A(_1653_),
    .B(_1658_),
    .C(_1670_),
    .D(_1819_),
    .X(_0606_));
 sky130_fd_sc_hd__or3_1 _3451_ (.A(_0603_),
    .B(_0604_),
    .C(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__a211o_1 _3452_ (.A1(_0913_),
    .A2(net173),
    .B1(_1578_),
    .C1(_0544_),
    .X(_0608_));
 sky130_fd_sc_hd__or3_1 _3453_ (.A(_1275_),
    .B(_1491_),
    .C(_0608_),
    .X(_0609_));
 sky130_fd_sc_hd__or3_1 _3454_ (.A(_1707_),
    .B(_1709_),
    .C(_0577_),
    .X(_0610_));
 sky130_fd_sc_hd__or4_2 _3455_ (.A(_1805_),
    .B(_1851_),
    .C(_0609_),
    .D(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__a31o_1 _3456_ (.A1(net272),
    .A2(_1045_),
    .A3(net99),
    .B1(_1785_),
    .X(_0612_));
 sky130_fd_sc_hd__or3_1 _3457_ (.A(_1465_),
    .B(_1468_),
    .C(_0612_),
    .X(_0613_));
 sky130_fd_sc_hd__or4_1 _3458_ (.A(_1803_),
    .B(_1804_),
    .C(_0079_),
    .D(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__or4_1 _3459_ (.A(_1249_),
    .B(_1734_),
    .C(_1739_),
    .D(_1765_),
    .X(_0615_));
 sky130_fd_sc_hd__or4_2 _3460_ (.A(_1435_),
    .B(_1545_),
    .C(_1680_),
    .D(_1687_),
    .X(_0617_));
 sky130_fd_sc_hd__or3_1 _3461_ (.A(_1281_),
    .B(_1577_),
    .C(_1589_),
    .X(_0618_));
 sky130_fd_sc_hd__or3_1 _3462_ (.A(_0615_),
    .B(_0617_),
    .C(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__or4_1 _3463_ (.A(_0607_),
    .B(_0611_),
    .C(_0614_),
    .D(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__or3_1 _3464_ (.A(_0598_),
    .B(_0602_),
    .C(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__a2111o_1 _3465_ (.A1(net40),
    .A2(_0621_),
    .B1(_0587_),
    .C1(_0533_),
    .D1(_0469_),
    .X(_0622_));
 sky130_fd_sc_hd__a21oi_4 _3466_ (.A1(net206),
    .A2(net170),
    .B1(net117),
    .Y(_0623_));
 sky130_fd_sc_hd__or4_4 _3467_ (.A(_1671_),
    .B(_1760_),
    .C(_0470_),
    .D(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__or4_2 _3468_ (.A(_1417_),
    .B(_1461_),
    .C(_1555_),
    .D(_1674_),
    .X(_0625_));
 sky130_fd_sc_hd__or3_2 _3469_ (.A(_1343_),
    .B(_1398_),
    .C(_1437_),
    .X(_0626_));
 sky130_fd_sc_hd__o41a_1 _3470_ (.A1(net243),
    .A2(_1146_),
    .A3(net152),
    .A4(net146),
    .B1(net83),
    .X(_0628_));
 sky130_fd_sc_hd__or2_4 _3471_ (.A(_1324_),
    .B(_1577_),
    .X(_0629_));
 sky130_fd_sc_hd__or3_4 _3472_ (.A(_1321_),
    .B(_1324_),
    .C(_1577_),
    .X(_0630_));
 sky130_fd_sc_hd__or2_4 _3473_ (.A(_0628_),
    .B(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__o41a_2 _3474_ (.A1(net178),
    .A2(net168),
    .A3(net140),
    .A4(net134),
    .B1(net98),
    .X(_0632_));
 sky130_fd_sc_hd__or3_2 _3475_ (.A(_1651_),
    .B(_0454_),
    .C(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__or3_1 _3476_ (.A(_1769_),
    .B(_0435_),
    .C(_0494_),
    .X(_0634_));
 sky130_fd_sc_hd__or4_2 _3477_ (.A(_0530_),
    .B(_0631_),
    .C(_0633_),
    .D(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__or4_1 _3478_ (.A(_1297_),
    .B(_1496_),
    .C(_1637_),
    .D(_1729_),
    .X(_0636_));
 sky130_fd_sc_hd__or4_1 _3479_ (.A(_0979_),
    .B(_1267_),
    .C(_1381_),
    .D(_1599_),
    .X(_0637_));
 sky130_fd_sc_hd__or4_1 _3480_ (.A(_1407_),
    .B(_1598_),
    .C(_0636_),
    .D(_0637_),
    .X(_0639_));
 sky130_fd_sc_hd__or4_1 _3481_ (.A(_1549_),
    .B(_1804_),
    .C(_1827_),
    .D(_1835_),
    .X(_0640_));
 sky130_fd_sc_hd__or4_2 _3482_ (.A(_1986_),
    .B(_1996_),
    .C(_0449_),
    .D(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__or4_1 _3483_ (.A(_1290_),
    .B(_1533_),
    .C(_1754_),
    .D(_1983_),
    .X(_0642_));
 sky130_fd_sc_hd__or4_1 _3484_ (.A(_1715_),
    .B(_1717_),
    .C(_1730_),
    .D(_1811_),
    .X(_0643_));
 sky130_fd_sc_hd__or3_1 _3485_ (.A(_1502_),
    .B(_1654_),
    .C(_1872_),
    .X(_0644_));
 sky130_fd_sc_hd__or4_1 _3486_ (.A(_1396_),
    .B(_0478_),
    .C(_0643_),
    .D(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__or4_1 _3487_ (.A(_0472_),
    .B(_0591_),
    .C(_0642_),
    .D(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__or4_1 _3488_ (.A(_0635_),
    .B(_0639_),
    .C(_0641_),
    .D(_0646_),
    .X(_0647_));
 sky130_fd_sc_hd__o41a_1 _3489_ (.A1(_0624_),
    .A2(_0625_),
    .A3(_0626_),
    .A4(_0647_),
    .B1(net31),
    .X(_0648_));
 sky130_fd_sc_hd__or4_4 _3490_ (.A(_1909_),
    .B(_1933_),
    .C(_1943_),
    .D(_1956_),
    .X(_0650_));
 sky130_fd_sc_hd__or3_1 _3491_ (.A(_1499_),
    .B(_1502_),
    .C(_1674_),
    .X(_0651_));
 sky130_fd_sc_hd__or3_1 _3492_ (.A(_1648_),
    .B(_1788_),
    .C(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__or2_2 _3493_ (.A(_1444_),
    .B(_1468_),
    .X(_0653_));
 sky130_fd_sc_hd__or2_4 _3494_ (.A(_1487_),
    .B(_1642_),
    .X(_0654_));
 sky130_fd_sc_hd__or4_2 _3495_ (.A(_1258_),
    .B(_1511_),
    .C(_0653_),
    .D(_0654_),
    .X(_0655_));
 sky130_fd_sc_hd__or4_1 _3496_ (.A(net76),
    .B(_1417_),
    .C(_1709_),
    .D(_1717_),
    .X(_0656_));
 sky130_fd_sc_hd__or3_4 _3497_ (.A(_1867_),
    .B(_1915_),
    .C(_0470_),
    .X(_0657_));
 sky130_fd_sc_hd__or4_1 _3498_ (.A(_0362_),
    .B(_0519_),
    .C(_0656_),
    .D(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__or4_1 _3499_ (.A(_0650_),
    .B(_0652_),
    .C(_0655_),
    .D(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__or3_4 _3500_ (.A(_1281_),
    .B(_1615_),
    .C(_1766_),
    .X(_0661_));
 sky130_fd_sc_hd__or2_2 _3501_ (.A(_1464_),
    .B(_1525_),
    .X(_0662_));
 sky130_fd_sc_hd__or2_2 _3502_ (.A(_1568_),
    .B(_1805_),
    .X(_0663_));
 sky130_fd_sc_hd__or4_1 _3503_ (.A(_1802_),
    .B(_0509_),
    .C(_0662_),
    .D(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__or3_1 _3504_ (.A(_1526_),
    .B(_1923_),
    .C(_0450_),
    .X(_0665_));
 sky130_fd_sc_hd__or4_1 _3505_ (.A(_1507_),
    .B(net28),
    .C(_0593_),
    .D(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__or3_1 _3506_ (.A(_0661_),
    .B(_0664_),
    .C(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__or4_1 _3507_ (.A(_1222_),
    .B(_1552_),
    .C(_1557_),
    .D(_1629_),
    .X(_0668_));
 sky130_fd_sc_hd__or4_1 _3508_ (.A(_1296_),
    .B(_1308_),
    .C(_1947_),
    .D(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__or4_1 _3509_ (.A(_1727_),
    .B(_1862_),
    .C(_1971_),
    .D(_1973_),
    .X(_0670_));
 sky130_fd_sc_hd__or2_1 _3510_ (.A(_2014_),
    .B(_0062_),
    .X(_0672_));
 sky130_fd_sc_hd__or4_1 _3511_ (.A(_1452_),
    .B(_1781_),
    .C(_2018_),
    .D(_0672_),
    .X(_0673_));
 sky130_fd_sc_hd__or3_1 _3512_ (.A(net94),
    .B(_1921_),
    .C(net13),
    .X(_0674_));
 sky130_fd_sc_hd__or4_1 _3513_ (.A(_1736_),
    .B(_1767_),
    .C(_1936_),
    .D(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__or4_4 _3514_ (.A(_0669_),
    .B(_0670_),
    .C(_0673_),
    .D(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__a2111o_1 _3515_ (.A1(net112),
    .A2(net139),
    .B1(_1689_),
    .C1(_1695_),
    .D1(net15),
    .X(_0677_));
 sky130_fd_sc_hd__or4_1 _3516_ (.A(_1390_),
    .B(net75),
    .C(_1441_),
    .D(_1469_),
    .X(_0678_));
 sky130_fd_sc_hd__or4_1 _3517_ (.A(net69),
    .B(_1792_),
    .C(_1795_),
    .D(_1890_),
    .X(_0679_));
 sky130_fd_sc_hd__or4_1 _3518_ (.A(_1412_),
    .B(_0677_),
    .C(_0678_),
    .D(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__or4_1 _3519_ (.A(_1538_),
    .B(_1541_),
    .C(_1760_),
    .D(_1870_),
    .X(_0681_));
 sky130_fd_sc_hd__or4_1 _3520_ (.A(_1283_),
    .B(_1555_),
    .C(_1556_),
    .D(_1561_),
    .X(_0683_));
 sky130_fd_sc_hd__or4_1 _3521_ (.A(_1292_),
    .B(_1461_),
    .C(_0681_),
    .D(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__or4_1 _3522_ (.A(_0667_),
    .B(_0676_),
    .C(_0680_),
    .D(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__o21a_1 _3523_ (.A1(_0659_),
    .A2(_0685_),
    .B1(_1902_),
    .X(_0686_));
 sky130_fd_sc_hd__or3_1 _3524_ (.A(_1513_),
    .B(_1792_),
    .C(_0571_),
    .X(_0687_));
 sky130_fd_sc_hd__or3_2 _3525_ (.A(_1694_),
    .B(_1695_),
    .C(_0474_),
    .X(_0688_));
 sky130_fd_sc_hd__o2111a_2 _3526_ (.A1(net211),
    .A2(net177),
    .B1(net251),
    .C1(net238),
    .D1(net220),
    .X(_0689_));
 sky130_fd_sc_hd__or2_1 _3527_ (.A(_1433_),
    .B(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__or4_2 _3528_ (.A(_0529_),
    .B(_0687_),
    .C(_0688_),
    .D(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__or3_4 _3529_ (.A(_1407_),
    .B(_1440_),
    .C(net74),
    .X(_0692_));
 sky130_fd_sc_hd__or4_1 _3530_ (.A(_1564_),
    .B(_1750_),
    .C(_1754_),
    .D(_0692_),
    .X(_0694_));
 sky130_fd_sc_hd__or4_1 _3531_ (.A(_1531_),
    .B(_1692_),
    .C(_0691_),
    .D(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__o41a_1 _3532_ (.A1(_0990_),
    .A2(net177),
    .A3(net141),
    .A4(net134),
    .B1(_1408_),
    .X(_0696_));
 sky130_fd_sc_hd__or4_2 _3533_ (.A(_1365_),
    .B(_1366_),
    .C(_0537_),
    .D(_0696_),
    .X(_0697_));
 sky130_fd_sc_hd__or3_2 _3534_ (.A(net75),
    .B(_1541_),
    .C(_1811_),
    .X(_0698_));
 sky130_fd_sc_hd__or3_1 _3535_ (.A(_0494_),
    .B(_0663_),
    .C(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__or4_2 _3536_ (.A(_1631_),
    .B(_0567_),
    .C(_0697_),
    .D(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__and3_2 _3537_ (.A(net264),
    .B(net125),
    .C(_1172_),
    .X(_0701_));
 sky130_fd_sc_hd__a21oi_4 _3538_ (.A1(net199),
    .A2(net166),
    .B1(net78),
    .Y(_0702_));
 sky130_fd_sc_hd__or4_1 _3539_ (.A(_1634_),
    .B(_0425_),
    .C(_0518_),
    .D(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__or4_1 _3540_ (.A(_1379_),
    .B(_1646_),
    .C(net15),
    .D(_0701_),
    .X(_0705_));
 sky130_fd_sc_hd__or4_1 _3541_ (.A(_1655_),
    .B(_1671_),
    .C(_1838_),
    .D(_0303_),
    .X(_0706_));
 sky130_fd_sc_hd__or4_1 _3542_ (.A(net70),
    .B(_1570_),
    .C(_1688_),
    .D(_1714_),
    .X(_0707_));
 sky130_fd_sc_hd__or4_2 _3543_ (.A(_1560_),
    .B(_0705_),
    .C(_0706_),
    .D(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__or4_1 _3544_ (.A(_1442_),
    .B(_1495_),
    .C(_1518_),
    .D(_1574_),
    .X(_0709_));
 sky130_fd_sc_hd__or4_1 _3545_ (.A(_1600_),
    .B(_1610_),
    .C(_1677_),
    .D(_1715_),
    .X(_0710_));
 sky130_fd_sc_hd__or4_4 _3546_ (.A(_1364_),
    .B(_1664_),
    .C(_0709_),
    .D(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__or4_1 _3547_ (.A(_1343_),
    .B(_1465_),
    .C(_1582_),
    .D(_1705_),
    .X(_0712_));
 sky130_fd_sc_hd__or4_1 _3548_ (.A(_1417_),
    .B(_1550_),
    .C(_1851_),
    .D(_1872_),
    .X(_0713_));
 sky130_fd_sc_hd__or3_2 _3549_ (.A(_1460_),
    .B(_1660_),
    .C(_0175_),
    .X(_0714_));
 sky130_fd_sc_hd__or3_1 _3550_ (.A(_0712_),
    .B(_0713_),
    .C(_0714_),
    .X(_0716_));
 sky130_fd_sc_hd__or4_1 _3551_ (.A(_0703_),
    .B(_0708_),
    .C(_0711_),
    .D(_0716_),
    .X(_0717_));
 sky130_fd_sc_hd__or4_1 _3552_ (.A(_0420_),
    .B(_0695_),
    .C(_0700_),
    .D(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__or3_1 _3553_ (.A(_1366_),
    .B(_1383_),
    .C(_1851_),
    .X(_0719_));
 sky130_fd_sc_hd__or2_1 _3554_ (.A(_0599_),
    .B(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__or3_1 _3555_ (.A(_1290_),
    .B(_1297_),
    .C(_1926_),
    .X(_0721_));
 sky130_fd_sc_hd__a41o_1 _3556_ (.A1(net240),
    .A2(net113),
    .A3(net149),
    .A4(net143),
    .B1(net86),
    .X(_0722_));
 sky130_fd_sc_hd__or4b_2 _3557_ (.A(_1694_),
    .B(_1695_),
    .C(_0518_),
    .D_N(_0722_),
    .X(_0723_));
 sky130_fd_sc_hd__or3_2 _3558_ (.A(_1618_),
    .B(_1794_),
    .C(_0568_),
    .X(_0724_));
 sky130_fd_sc_hd__or3_1 _3559_ (.A(_1867_),
    .B(_1915_),
    .C(_0593_),
    .X(_0725_));
 sky130_fd_sc_hd__or3_1 _3560_ (.A(_1445_),
    .B(_1550_),
    .C(_0450_),
    .X(_0727_));
 sky130_fd_sc_hd__or4_4 _3561_ (.A(_1301_),
    .B(_1469_),
    .C(net15),
    .D(_1923_),
    .X(_0728_));
 sky130_fd_sc_hd__or4_1 _3562_ (.A(_1442_),
    .B(_1454_),
    .C(_1976_),
    .D(_0082_),
    .X(_0729_));
 sky130_fd_sc_hd__or3_1 _3563_ (.A(_1431_),
    .B(_1463_),
    .C(_1615_),
    .X(_0730_));
 sky130_fd_sc_hd__or4_1 _3564_ (.A(_1418_),
    .B(_1684_),
    .C(_0729_),
    .D(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__or4_1 _3565_ (.A(_1276_),
    .B(_1531_),
    .C(_0417_),
    .D(_0687_),
    .X(_0732_));
 sky130_fd_sc_hd__or3_2 _3566_ (.A(_1470_),
    .B(_1629_),
    .C(_1806_),
    .X(_0733_));
 sky130_fd_sc_hd__or4_1 _3567_ (.A(_0434_),
    .B(_0515_),
    .C(_0689_),
    .D(_0702_),
    .X(_0734_));
 sky130_fd_sc_hd__or3_1 _3568_ (.A(_0728_),
    .B(_0733_),
    .C(_0734_),
    .X(_0735_));
 sky130_fd_sc_hd__or2_1 _3569_ (.A(_1693_),
    .B(_0601_),
    .X(_0736_));
 sky130_fd_sc_hd__or4_1 _3570_ (.A(_0731_),
    .B(_0732_),
    .C(_0735_),
    .D(_0736_),
    .X(_0738_));
 sky130_fd_sc_hd__or3_1 _3571_ (.A(_0488_),
    .B(_0523_),
    .C(_0723_),
    .X(_0739_));
 sky130_fd_sc_hd__or4_1 _3572_ (.A(_0442_),
    .B(_0596_),
    .C(_0725_),
    .D(_0727_),
    .X(_0740_));
 sky130_fd_sc_hd__or4_1 _3573_ (.A(_0514_),
    .B(_0721_),
    .C(_0724_),
    .D(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__or4_1 _3574_ (.A(_0720_),
    .B(_0738_),
    .C(_0739_),
    .D(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__a22o_1 _3575_ (.A1(net63),
    .A2(_0718_),
    .B1(_0742_),
    .B2(net26),
    .X(_0743_));
 sky130_fd_sc_hd__or4_4 _3576_ (.A(_0622_),
    .B(_0648_),
    .C(_0686_),
    .D(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__or4_2 _3577_ (.A(_1267_),
    .B(_1985_),
    .C(_0571_),
    .D(_0663_),
    .X(_0745_));
 sky130_fd_sc_hd__or3_1 _3578_ (.A(_1461_),
    .B(_1672_),
    .C(_1674_),
    .X(_0746_));
 sky130_fd_sc_hd__or4_1 _3579_ (.A(_1634_),
    .B(_1700_),
    .C(_1730_),
    .D(_0434_),
    .X(_0747_));
 sky130_fd_sc_hd__or4_1 _3580_ (.A(_1867_),
    .B(_1915_),
    .C(_0444_),
    .D(_0518_),
    .X(_0749_));
 sky130_fd_sc_hd__or4_1 _3581_ (.A(_0634_),
    .B(_0746_),
    .C(_0747_),
    .D(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__or4_1 _3582_ (.A(_0433_),
    .B(_0656_),
    .C(_0698_),
    .D(_0721_),
    .X(_0751_));
 sky130_fd_sc_hd__or4_1 _3583_ (.A(_1947_),
    .B(_0428_),
    .C(_0745_),
    .D(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__or3_1 _3584_ (.A(_0624_),
    .B(_0750_),
    .C(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__or3_2 _3585_ (.A(_1362_),
    .B(_1380_),
    .C(_1804_),
    .X(_0754_));
 sky130_fd_sc_hd__a21oi_4 _3586_ (.A1(net206),
    .A2(net175),
    .B1(net97),
    .Y(_0755_));
 sky130_fd_sc_hd__or3_2 _3587_ (.A(net76),
    .B(_1417_),
    .C(_1672_),
    .X(_0756_));
 sky130_fd_sc_hd__o41a_4 _3588_ (.A1(net211),
    .A2(net177),
    .A3(net172),
    .A4(net141),
    .B1(net84),
    .X(_0757_));
 sky130_fd_sc_hd__or2_2 _3589_ (.A(_1354_),
    .B(_1396_),
    .X(_0758_));
 sky130_fd_sc_hd__or4_1 _3590_ (.A(_1545_),
    .B(_1951_),
    .C(_0444_),
    .D(_0571_),
    .X(_0760_));
 sky130_fd_sc_hd__or4_1 _3591_ (.A(_0437_),
    .B(_0475_),
    .C(_0699_),
    .D(_0758_),
    .X(_0761_));
 sky130_fd_sc_hd__or4_1 _3592_ (.A(_1490_),
    .B(net72),
    .C(_1535_),
    .D(_1549_),
    .X(_0762_));
 sky130_fd_sc_hd__or4_1 _3593_ (.A(_1321_),
    .B(net82),
    .C(_1349_),
    .D(_1673_),
    .X(_0763_));
 sky130_fd_sc_hd__or4_1 _3594_ (.A(_1382_),
    .B(_1755_),
    .C(_0762_),
    .D(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__or4_1 _3595_ (.A(_1703_),
    .B(_0760_),
    .C(_0761_),
    .D(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__or4_1 _3596_ (.A(_1034_),
    .B(_1678_),
    .C(_1679_),
    .D(_0428_),
    .X(_0766_));
 sky130_fd_sc_hd__or4_1 _3597_ (.A(_1459_),
    .B(net67),
    .C(_2016_),
    .D(_0084_),
    .X(_0767_));
 sky130_fd_sc_hd__or4_1 _3598_ (.A(_1375_),
    .B(_1454_),
    .C(_1644_),
    .D(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__or4_1 _3599_ (.A(_1322_),
    .B(_1517_),
    .C(net27),
    .D(_1578_),
    .X(_0769_));
 sky130_fd_sc_hd__or3_1 _3600_ (.A(_1761_),
    .B(_0768_),
    .C(_0769_),
    .X(_0771_));
 sky130_fd_sc_hd__or4_1 _3601_ (.A(_0628_),
    .B(_0756_),
    .C(_0766_),
    .D(_0771_),
    .X(_0772_));
 sky130_fd_sc_hd__or4_1 _3602_ (.A(_1447_),
    .B(_0719_),
    .C(_0754_),
    .D(_0755_),
    .X(_0773_));
 sky130_fd_sc_hd__or3_1 _3603_ (.A(_0626_),
    .B(_0657_),
    .C(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__or3_1 _3604_ (.A(_0765_),
    .B(_0772_),
    .C(_0774_),
    .X(_0775_));
 sky130_fd_sc_hd__o41a_4 _3605_ (.A1(net205),
    .A2(net195),
    .A3(_1277_),
    .A4(net135),
    .B1(net105),
    .X(_0776_));
 sky130_fd_sc_hd__or2_1 _3606_ (.A(_1639_),
    .B(net14),
    .X(_0777_));
 sky130_fd_sc_hd__nand2_1 _3607_ (.A(_1668_),
    .B(_0559_),
    .Y(_0778_));
 sky130_fd_sc_hd__or4_4 _3608_ (.A(_1458_),
    .B(_0776_),
    .C(_0777_),
    .D(_0778_),
    .X(_0779_));
 sky130_fd_sc_hd__or3_1 _3609_ (.A(_1607_),
    .B(_1618_),
    .C(_1794_),
    .X(_0780_));
 sky130_fd_sc_hd__a21oi_4 _3610_ (.A1(net241),
    .A2(_1236_),
    .B1(net78),
    .Y(_0782_));
 sky130_fd_sc_hd__a21o_2 _3611_ (.A1(net187),
    .A2(net83),
    .B1(_1388_),
    .X(_0783_));
 sky130_fd_sc_hd__or4_1 _3612_ (.A(_0653_),
    .B(_0780_),
    .C(_0782_),
    .D(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__or2_4 _3613_ (.A(_1434_),
    .B(_1548_),
    .X(_0785_));
 sky130_fd_sc_hd__or4_2 _3614_ (.A(_1433_),
    .B(_1519_),
    .C(_0527_),
    .D(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__or4_1 _3615_ (.A(_1577_),
    .B(_1762_),
    .C(_0521_),
    .D(_0689_),
    .X(_0787_));
 sky130_fd_sc_hd__or3_1 _3616_ (.A(_1686_),
    .B(_0786_),
    .C(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__or4_1 _3617_ (.A(_1368_),
    .B(_1395_),
    .C(_1488_),
    .D(_1545_),
    .X(_0789_));
 sky130_fd_sc_hd__or4_2 _3618_ (.A(_0935_),
    .B(_1844_),
    .C(_1920_),
    .D(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__or3_1 _3619_ (.A(_1358_),
    .B(_1745_),
    .C(_1748_),
    .X(_0791_));
 sky130_fd_sc_hd__or4_1 _3620_ (.A(_1163_),
    .B(_1377_),
    .C(_1881_),
    .D(net67),
    .X(_0793_));
 sky130_fd_sc_hd__or2_1 _3621_ (.A(_1321_),
    .B(_1346_),
    .X(_0794_));
 sky130_fd_sc_hd__or4_1 _3622_ (.A(_1533_),
    .B(_1565_),
    .C(_1601_),
    .D(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__or4_1 _3623_ (.A(_1984_),
    .B(_0370_),
    .C(_0793_),
    .D(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__or4_2 _3624_ (.A(_0788_),
    .B(_0790_),
    .C(_0791_),
    .D(_0796_),
    .X(_0797_));
 sky130_fd_sc_hd__o41a_1 _3625_ (.A1(_0720_),
    .A2(_0779_),
    .A3(_0784_),
    .A4(_0797_),
    .B1(_1493_),
    .X(_0798_));
 sky130_fd_sc_hd__a221o_4 _3626_ (.A1(net34),
    .A2(_0753_),
    .B1(_0775_),
    .B2(net21),
    .C1(_0798_),
    .X(_0799_));
 sky130_fd_sc_hd__or4_2 _3627_ (.A(_1880_),
    .B(_0228_),
    .C(_0316_),
    .D(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__or4_1 _3628_ (.A(_1331_),
    .B(_1388_),
    .C(_1618_),
    .D(_1680_),
    .X(_0801_));
 sky130_fd_sc_hd__a41o_2 _3629_ (.A1(net113),
    .A2(net106),
    .A3(net91),
    .A4(net149),
    .B1(_1359_),
    .X(_0802_));
 sky130_fd_sc_hd__or4b_1 _3630_ (.A(_0499_),
    .B(_0757_),
    .C(_0801_),
    .D_N(_0802_),
    .X(_0804_));
 sky130_fd_sc_hd__o31a_2 _3631_ (.A1(_1601_),
    .A2(_0481_),
    .A3(_0804_),
    .B1(net34),
    .X(_0805_));
 sky130_fd_sc_hd__a211o_2 _3632_ (.A1(_0957_),
    .A2(_1138_),
    .B1(_1354_),
    .C1(_1357_),
    .X(_0806_));
 sky130_fd_sc_hd__a21oi_1 _3633_ (.A1(net101),
    .A2(net93),
    .B1(net102),
    .Y(_0807_));
 sky130_fd_sc_hd__a31o_4 _3634_ (.A1(net108),
    .A2(net101),
    .A3(net92),
    .B1(net103),
    .X(_0808_));
 sky130_fd_sc_hd__or4b_4 _3635_ (.A(_0782_),
    .B(_0783_),
    .C(_0806_),
    .D_N(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__or2_2 _3636_ (.A(_1495_),
    .B(_1881_),
    .X(_0810_));
 sky130_fd_sc_hd__and3_1 _3637_ (.A(net226),
    .B(net219),
    .C(net203),
    .X(_0811_));
 sky130_fd_sc_hd__or4_1 _3638_ (.A(_1921_),
    .B(_0262_),
    .C(_0810_),
    .D(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__or3_1 _3639_ (.A(_1485_),
    .B(_1494_),
    .C(_0776_),
    .X(_0813_));
 sky130_fd_sc_hd__o31a_1 _3640_ (.A1(_0809_),
    .A2(_0812_),
    .A3(_0813_),
    .B1(net24),
    .X(_0815_));
 sky130_fd_sc_hd__or4_4 _3641_ (.A(_1607_),
    .B(_1705_),
    .C(_0474_),
    .D(_0499_),
    .X(_0816_));
 sky130_fd_sc_hd__or4_1 _3642_ (.A(_1355_),
    .B(_1850_),
    .C(_0783_),
    .D(_0810_),
    .X(_0817_));
 sky130_fd_sc_hd__nor2_1 _3643_ (.A(_1379_),
    .B(_1682_),
    .Y(_0818_));
 sky130_fd_sc_hd__or4_1 _3644_ (.A(_1347_),
    .B(_1379_),
    .C(_1595_),
    .D(_1682_),
    .X(_0819_));
 sky130_fd_sc_hd__o31a_2 _3645_ (.A1(_0816_),
    .A2(_0817_),
    .A3(_0819_),
    .B1(net59),
    .X(_0820_));
 sky130_fd_sc_hd__or4_2 _3646_ (.A(_0348_),
    .B(_0805_),
    .C(_0815_),
    .D(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__a211o_1 _3647_ (.A1(net62),
    .A2(_1920_),
    .B1(_0237_),
    .C1(_0317_),
    .X(_0822_));
 sky130_fd_sc_hd__or4_2 _3648_ (.A(_1893_),
    .B(_1979_),
    .C(_0821_),
    .D(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__or3_2 _3649_ (.A(_1410_),
    .B(_1442_),
    .C(_0782_),
    .X(_0824_));
 sky130_fd_sc_hd__or3_4 _3650_ (.A(_1640_),
    .B(net16),
    .C(net14),
    .X(_0826_));
 sky130_fd_sc_hd__and3_1 _3651_ (.A(net264),
    .B(_1045_),
    .C(net89),
    .X(_0827_));
 sky130_fd_sc_hd__a22o_1 _3652_ (.A1(_1146_),
    .A2(_1205_),
    .B1(net89),
    .B2(net243),
    .X(_0828_));
 sky130_fd_sc_hd__or4_1 _3653_ (.A(_1636_),
    .B(_0702_),
    .C(_0827_),
    .D(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__or3_1 _3654_ (.A(_1628_),
    .B(_1630_),
    .C(_1692_),
    .X(_0830_));
 sky130_fd_sc_hd__or4_4 _3655_ (.A(_0824_),
    .B(_0826_),
    .C(_0829_),
    .D(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__o31a_1 _3656_ (.A1(_0654_),
    .A2(_0696_),
    .A3(_0831_),
    .B1(net23),
    .X(_0832_));
 sky130_fd_sc_hd__or4_2 _3657_ (.A(_1360_),
    .B(_1463_),
    .C(_1525_),
    .D(_1851_),
    .X(_0833_));
 sky130_fd_sc_hd__or4_1 _3658_ (.A(_1750_),
    .B(_0525_),
    .C(_0663_),
    .D(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__o31a_1 _3659_ (.A1(_0631_),
    .A2(_0758_),
    .A3(_0834_),
    .B1(_1427_),
    .X(_0835_));
 sky130_fd_sc_hd__nor2_1 _3660_ (.A(_0078_),
    .B(_0493_),
    .Y(_0837_));
 sky130_fd_sc_hd__or3b_1 _3661_ (.A(_1607_),
    .B(_1705_),
    .C_N(_0818_),
    .X(_0838_));
 sky130_fd_sc_hd__o41a_1 _3662_ (.A1(net197),
    .A2(net183),
    .A3(net154),
    .A4(net151),
    .B1(_0957_),
    .X(_0839_));
 sky130_fd_sc_hd__or2_1 _3663_ (.A(_1742_),
    .B(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__or4b_2 _3664_ (.A(_1766_),
    .B(_0078_),
    .C(_0493_),
    .D_N(_0808_),
    .X(_0841_));
 sky130_fd_sc_hd__o41a_1 _3665_ (.A1(_1285_),
    .A2(_0838_),
    .A3(_0840_),
    .A4(_0841_),
    .B1(net52),
    .X(_0842_));
 sky130_fd_sc_hd__or3_1 _3666_ (.A(_1377_),
    .B(_1495_),
    .C(_1680_),
    .X(_0843_));
 sky130_fd_sc_hd__or3_1 _3667_ (.A(_1565_),
    .B(_1575_),
    .C(_1595_),
    .X(_0844_));
 sky130_fd_sc_hd__or4_1 _3668_ (.A(_1344_),
    .B(_0839_),
    .C(_0843_),
    .D(_0844_),
    .X(_0845_));
 sky130_fd_sc_hd__or4_1 _3669_ (.A(_1577_),
    .B(_1579_),
    .C(_1762_),
    .D(_1950_),
    .X(_0846_));
 sky130_fd_sc_hd__o31a_1 _3670_ (.A1(_0816_),
    .A2(_0845_),
    .A3(_0846_),
    .B1(net47),
    .X(_0848_));
 sky130_fd_sc_hd__or3_1 _3671_ (.A(_1342_),
    .B(_1544_),
    .C(_1549_),
    .X(_0849_));
 sky130_fd_sc_hd__or3_1 _3672_ (.A(_1368_),
    .B(_1397_),
    .C(_0689_),
    .X(_0850_));
 sky130_fd_sc_hd__o41a_1 _3673_ (.A1(net177),
    .A2(net168),
    .A3(net141),
    .A4(net134),
    .B1(net84),
    .X(_0851_));
 sky130_fd_sc_hd__or4_1 _3674_ (.A(_0481_),
    .B(_0849_),
    .C(_0850_),
    .D(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__o31a_1 _3675_ (.A1(_0479_),
    .A2(_0631_),
    .A3(_0852_),
    .B1(_1372_),
    .X(_0853_));
 sky130_fd_sc_hd__or4_1 _3676_ (.A(_1806_),
    .B(_0360_),
    .C(_0363_),
    .D(_0630_),
    .X(_0854_));
 sky130_fd_sc_hd__or3_1 _3677_ (.A(_1397_),
    .B(_1527_),
    .C(_1795_),
    .X(_0855_));
 sky130_fd_sc_hd__or4_1 _3678_ (.A(_1308_),
    .B(_1430_),
    .C(_1745_),
    .D(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__o31a_1 _3679_ (.A1(_0758_),
    .A2(_0854_),
    .A3(_0856_),
    .B1(net43),
    .X(_0857_));
 sky130_fd_sc_hd__or3_1 _3680_ (.A(_1575_),
    .B(_0480_),
    .C(_0629_),
    .X(_0859_));
 sky130_fd_sc_hd__nand2_1 _3681_ (.A(_0802_),
    .B(_0818_),
    .Y(_0860_));
 sky130_fd_sc_hd__o41a_1 _3682_ (.A1(_0816_),
    .A2(_0840_),
    .A3(_0859_),
    .A4(_0860_),
    .B1(net55),
    .X(_0861_));
 sky130_fd_sc_hd__or4_1 _3683_ (.A(_0848_),
    .B(_0853_),
    .C(_0857_),
    .D(_0861_),
    .X(_0862_));
 sky130_fd_sc_hd__or4_4 _3684_ (.A(_0832_),
    .B(_0835_),
    .C(_0842_),
    .D(_0862_),
    .X(_0863_));
 sky130_fd_sc_hd__or3_4 _3685_ (.A(_0141_),
    .B(_0422_),
    .C(_0493_),
    .X(_0864_));
 sky130_fd_sc_hd__o41a_1 _3686_ (.A1(_1881_),
    .A2(_2009_),
    .A3(_0447_),
    .A4(_0864_),
    .B1(net31),
    .X(_0865_));
 sky130_fd_sc_hd__or4_1 _3687_ (.A(_1391_),
    .B(_1432_),
    .C(_1434_),
    .D(_1569_),
    .X(_0866_));
 sky130_fd_sc_hd__or4_1 _3688_ (.A(_1368_),
    .B(_1394_),
    .C(_1454_),
    .D(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__o41a_1 _3689_ (.A1(_1549_),
    .A2(_1745_),
    .A3(_0755_),
    .A4(_0867_),
    .B1(net60),
    .X(_0868_));
 sky130_fd_sc_hd__or4_1 _3690_ (.A(_1691_),
    .B(_1701_),
    .C(_1707_),
    .D(_1714_),
    .X(_0870_));
 sky130_fd_sc_hd__o21a_1 _3691_ (.A1(_0688_),
    .A2(_0870_),
    .B1(net33),
    .X(_0871_));
 sky130_fd_sc_hd__a2111o_1 _3692_ (.A1(net125),
    .A2(net152),
    .B1(_1406_),
    .C1(_1432_),
    .D1(_1568_),
    .X(_0872_));
 sky130_fd_sc_hd__o41a_1 _3693_ (.A1(_1472_),
    .A2(_1628_),
    .A3(_0785_),
    .A4(_0872_),
    .B1(net26),
    .X(_0873_));
 sky130_fd_sc_hd__or4_1 _3694_ (.A(_0865_),
    .B(_0868_),
    .C(_0871_),
    .D(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__or4_1 _3695_ (.A(_1301_),
    .B(_1469_),
    .C(_1756_),
    .D(_0782_),
    .X(_0875_));
 sky130_fd_sc_hd__or3_1 _3696_ (.A(_1243_),
    .B(_1623_),
    .C(_1629_),
    .X(_0876_));
 sky130_fd_sc_hd__o31a_1 _3697_ (.A1(_0596_),
    .A2(_0875_),
    .A3(_0876_),
    .B1(net55),
    .X(_0877_));
 sky130_fd_sc_hd__a211o_1 _3698_ (.A1(_1288_),
    .A2(net147),
    .B1(_1331_),
    .C1(_1763_),
    .X(_0878_));
 sky130_fd_sc_hd__or3_2 _3699_ (.A(_1281_),
    .B(_1764_),
    .C(_0590_),
    .X(_0879_));
 sky130_fd_sc_hd__o41a_1 _3700_ (.A1(_1422_),
    .A2(_1634_),
    .A3(_0878_),
    .A4(_0879_),
    .B1(net23),
    .X(_0881_));
 sky130_fd_sc_hd__or3_1 _3701_ (.A(_1568_),
    .B(_1684_),
    .C(_1802_),
    .X(_0882_));
 sky130_fd_sc_hd__or4_2 _3702_ (.A(_1254_),
    .B(_1564_),
    .C(_1591_),
    .D(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__o31a_1 _3703_ (.A1(_1735_),
    .A2(_0724_),
    .A3(_0883_),
    .B1(net49),
    .X(_0884_));
 sky130_fd_sc_hd__o31a_1 _3704_ (.A1(_1669_),
    .A2(_1824_),
    .A3(_1844_),
    .B1(net62),
    .X(_0885_));
 sky130_fd_sc_hd__or4_1 _3705_ (.A(_0877_),
    .B(_0881_),
    .C(_0884_),
    .D(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__or3_1 _3706_ (.A(_1577_),
    .B(_1762_),
    .C(_1768_),
    .X(_0887_));
 sky130_fd_sc_hd__or4b_1 _3707_ (.A(_1485_),
    .B(_1501_),
    .C(_1575_),
    .D_N(_1659_),
    .X(_0888_));
 sky130_fd_sc_hd__or4_1 _3708_ (.A(_1489_),
    .B(_1656_),
    .C(_0085_),
    .D(_0887_),
    .X(_0889_));
 sky130_fd_sc_hd__o21a_1 _3709_ (.A1(_0888_),
    .A2(_0889_),
    .B1(net19),
    .X(_0890_));
 sky130_fd_sc_hd__or2_1 _3710_ (.A(_1724_),
    .B(_1745_),
    .X(_0892_));
 sky130_fd_sc_hd__or4_2 _3711_ (.A(_1308_),
    .B(_1466_),
    .C(_1613_),
    .D(_1646_),
    .X(_0893_));
 sky130_fd_sc_hd__or4_1 _3712_ (.A(_1444_),
    .B(_1471_),
    .C(_1726_),
    .D(_0425_),
    .X(_0894_));
 sky130_fd_sc_hd__o31a_1 _3713_ (.A1(_0892_),
    .A2(_0893_),
    .A3(_0894_),
    .B1(net37),
    .X(_0895_));
 sky130_fd_sc_hd__o41a_1 _3714_ (.A1(net243),
    .A2(net195),
    .A3(_1230_),
    .A4(net147),
    .B1(net84),
    .X(_0896_));
 sky130_fd_sc_hd__or4_4 _3715_ (.A(_1345_),
    .B(_0478_),
    .C(_0480_),
    .D(_0630_),
    .X(_0897_));
 sky130_fd_sc_hd__o21a_1 _3716_ (.A1(_0896_),
    .A2(_0897_),
    .B1(net52),
    .X(_0898_));
 sky130_fd_sc_hd__or4_1 _3717_ (.A(_1280_),
    .B(_1283_),
    .C(_1309_),
    .D(_1881_),
    .X(_0899_));
 sky130_fd_sc_hd__or4_1 _3718_ (.A(_1291_),
    .B(_1296_),
    .C(_1490_),
    .D(_1736_),
    .X(_0900_));
 sky130_fd_sc_hd__o21a_1 _3719_ (.A1(_0899_),
    .A2(_0900_),
    .B1(net66),
    .X(_0901_));
 sky130_fd_sc_hd__or4_1 _3720_ (.A(_0890_),
    .B(_0895_),
    .C(_0898_),
    .D(_0901_),
    .X(_0903_));
 sky130_fd_sc_hd__or4_1 _3721_ (.A(_1888_),
    .B(_0874_),
    .C(_0886_),
    .D(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__a22o_1 _3722_ (.A1(net65),
    .A2(_1746_),
    .B1(_0807_),
    .B2(_1372_),
    .X(_0905_));
 sky130_fd_sc_hd__o21a_1 _3723_ (.A1(_1319_),
    .A2(_1428_),
    .B1(net40),
    .X(_0906_));
 sky130_fd_sc_hd__a211o_1 _3724_ (.A1(net60),
    .A2(_1395_),
    .B1(_0905_),
    .C1(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__or2_1 _3725_ (.A(_1747_),
    .B(_0078_),
    .X(_0908_));
 sky130_fd_sc_hd__a22o_1 _3726_ (.A1(net75),
    .A2(net31),
    .B1(_0908_),
    .B2(_1372_),
    .X(_0909_));
 sky130_fd_sc_hd__or3b_1 _3727_ (.A(net76),
    .B(_1487_),
    .C_N(_1645_),
    .X(_0910_));
 sky130_fd_sc_hd__o31a_1 _3728_ (.A1(_1445_),
    .A2(_1764_),
    .A3(_0910_),
    .B1(net40),
    .X(_0911_));
 sky130_fd_sc_hd__o31a_1 _3729_ (.A1(_1365_),
    .A2(_1368_),
    .A3(_1555_),
    .B1(net20),
    .X(_0912_));
 sky130_fd_sc_hd__or4_1 _3730_ (.A(_0907_),
    .B(_0909_),
    .C(_0911_),
    .D(_0912_),
    .X(_0914_));
 sky130_fd_sc_hd__and2b_1 _3731_ (.A_N(_0808_),
    .B(_1451_),
    .X(_0915_));
 sky130_fd_sc_hd__o21a_1 _3732_ (.A1(_1345_),
    .A2(_1356_),
    .B1(net20),
    .X(_0916_));
 sky130_fd_sc_hd__o41a_1 _3733_ (.A1(_1378_),
    .A2(_1390_),
    .A3(_1428_),
    .A4(_0757_),
    .B1(net55),
    .X(_0917_));
 sky130_fd_sc_hd__o21a_1 _3734_ (.A1(_1254_),
    .A2(_1844_),
    .B1(net33),
    .X(_0918_));
 sky130_fd_sc_hd__o41a_2 _3735_ (.A1(_1374_),
    .A2(_2016_),
    .A3(_0476_),
    .A4(_0521_),
    .B1(net47),
    .X(_0919_));
 sky130_fd_sc_hd__o31a_1 _3736_ (.A1(_1258_),
    .A2(_1328_),
    .A3(_1479_),
    .B1(net35),
    .X(_0920_));
 sky130_fd_sc_hd__or4_1 _3737_ (.A(_0917_),
    .B(_0918_),
    .C(_0919_),
    .D(_0920_),
    .X(_0921_));
 sky130_fd_sc_hd__a2111o_1 _3738_ (.A1(net52),
    .A2(_1947_),
    .B1(_0915_),
    .C1(_0916_),
    .D1(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__or4b_1 _3739_ (.A(_0074_),
    .B(_0177_),
    .C(_0235_),
    .D_N(_0413_),
    .X(_0923_));
 sky130_fd_sc_hd__or4_1 _3740_ (.A(_1903_),
    .B(_1980_),
    .C(_0068_),
    .D(_0182_),
    .X(_0925_));
 sky130_fd_sc_hd__or3_1 _3741_ (.A(_1901_),
    .B(_2031_),
    .C(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__or4_1 _3742_ (.A(_0914_),
    .B(_0922_),
    .C(_0923_),
    .D(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__or4_1 _3743_ (.A(_0823_),
    .B(_0863_),
    .C(_0904_),
    .D(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__or4b_1 _3744_ (.A(_1679_),
    .B(_0593_),
    .C(_1699_),
    .D_N(_0505_),
    .X(_0929_));
 sky130_fd_sc_hd__or3_1 _3745_ (.A(_1610_),
    .B(_1792_),
    .C(_0416_),
    .X(_0930_));
 sky130_fd_sc_hd__or4_1 _3746_ (.A(_1397_),
    .B(_1590_),
    .C(_1596_),
    .D(_1736_),
    .X(_0931_));
 sky130_fd_sc_hd__or4_1 _3747_ (.A(_0745_),
    .B(_0929_),
    .C(_0930_),
    .D(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__or4_1 _3748_ (.A(_1717_),
    .B(net13),
    .C(_0243_),
    .D(_0447_),
    .X(_0933_));
 sky130_fd_sc_hd__or3b_1 _3749_ (.A(_1731_),
    .B(_2016_),
    .C_N(_1659_),
    .X(_0934_));
 sky130_fd_sc_hd__or4_1 _3750_ (.A(_0468_),
    .B(_0642_),
    .C(_0933_),
    .D(_0934_),
    .X(_0936_));
 sky130_fd_sc_hd__or4b_2 _3751_ (.A(_0088_),
    .B(_0141_),
    .C(_0521_),
    .D_N(_0802_),
    .X(_0937_));
 sky130_fd_sc_hd__or4_1 _3752_ (.A(_1413_),
    .B(_1418_),
    .C(_1678_),
    .D(_1868_),
    .X(_0938_));
 sky130_fd_sc_hd__or4_2 _3753_ (.A(_0540_),
    .B(_0754_),
    .C(_0937_),
    .D(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__or3_1 _3754_ (.A(_0932_),
    .B(_0936_),
    .C(_0939_),
    .X(_0940_));
 sky130_fd_sc_hd__or3b_1 _3755_ (.A(_1615_),
    .B(_1688_),
    .C_N(_0808_),
    .X(_0941_));
 sky130_fd_sc_hd__or4_1 _3756_ (.A(_1502_),
    .B(_1637_),
    .C(_0507_),
    .D(_0941_),
    .X(_0942_));
 sky130_fd_sc_hd__nand2b_1 _3757_ (.A_N(_1643_),
    .B(_0722_),
    .Y(_0943_));
 sky130_fd_sc_hd__a21o_1 _3758_ (.A1(net125),
    .A2(_1269_),
    .B1(_1722_),
    .X(_0944_));
 sky130_fd_sc_hd__or4_2 _3759_ (.A(_1373_),
    .B(_1592_),
    .C(_1610_),
    .D(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__or3_1 _3760_ (.A(_1674_),
    .B(_1678_),
    .C(_1691_),
    .X(_0947_));
 sky130_fd_sc_hd__or2_1 _3761_ (.A(_1296_),
    .B(_1423_),
    .X(_0948_));
 sky130_fd_sc_hd__or4_2 _3762_ (.A(_1508_),
    .B(_1582_),
    .C(_1724_),
    .D(_0948_),
    .X(_0949_));
 sky130_fd_sc_hd__or4_1 _3763_ (.A(_0943_),
    .B(_0945_),
    .C(_0947_),
    .D(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__or4_1 _3764_ (.A(_1281_),
    .B(_1284_),
    .C(_1764_),
    .D(_0493_),
    .X(_0951_));
 sky130_fd_sc_hd__or4_2 _3765_ (.A(_1545_),
    .B(_1951_),
    .C(_0449_),
    .D(_0483_),
    .X(_0952_));
 sky130_fd_sc_hd__or4_1 _3766_ (.A(_0426_),
    .B(_0520_),
    .C(_0951_),
    .D(_0952_),
    .X(_0953_));
 sky130_fd_sc_hd__or4_1 _3767_ (.A(_0088_),
    .B(_0287_),
    .C(_0366_),
    .D(_0701_),
    .X(_0954_));
 sky130_fd_sc_hd__or4_1 _3768_ (.A(_1672_),
    .B(_1765_),
    .C(_0078_),
    .D(_0107_),
    .X(_0955_));
 sky130_fd_sc_hd__a21o_1 _3769_ (.A1(net98),
    .A2(net152),
    .B1(_0084_),
    .X(_0956_));
 sky130_fd_sc_hd__or4_1 _3770_ (.A(net15),
    .B(_1923_),
    .C(_0515_),
    .D(_0956_),
    .X(_0958_));
 sky130_fd_sc_hd__or4_1 _3771_ (.A(_1771_),
    .B(_0954_),
    .C(_0955_),
    .D(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__or4_2 _3772_ (.A(_0942_),
    .B(_0950_),
    .C(_0953_),
    .D(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__a22o_1 _3773_ (.A1(net59),
    .A2(_0940_),
    .B1(_0960_),
    .B2(net47),
    .X(_0961_));
 sky130_fd_sc_hd__or4_1 _3774_ (.A(_0454_),
    .B(_0629_),
    .C(_0662_),
    .D(_0782_),
    .X(_0962_));
 sky130_fd_sc_hd__or3_1 _3775_ (.A(_1654_),
    .B(_1872_),
    .C(_0527_),
    .X(_0963_));
 sky130_fd_sc_hd__or4_1 _3776_ (.A(_1772_),
    .B(_2014_),
    .C(_0962_),
    .D(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__or4_1 _3777_ (.A(net70),
    .B(_1570_),
    .C(_1742_),
    .D(_0453_),
    .X(_0965_));
 sky130_fd_sc_hd__or3_1 _3778_ (.A(_0558_),
    .B(_0806_),
    .C(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__or4_1 _3779_ (.A(_1280_),
    .B(_1575_),
    .C(_1639_),
    .D(_1762_),
    .X(_0967_));
 sky130_fd_sc_hd__or4_1 _3780_ (.A(_1290_),
    .B(net94),
    .C(_1394_),
    .D(_1395_),
    .X(_0969_));
 sky130_fd_sc_hd__or4_2 _3781_ (.A(_1430_),
    .B(_1586_),
    .C(_0967_),
    .D(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__or4_2 _3782_ (.A(_1284_),
    .B(_0483_),
    .C(_0493_),
    .D(_0692_),
    .X(_0971_));
 sky130_fd_sc_hd__or4_1 _3783_ (.A(_0625_),
    .B(_0966_),
    .C(_0970_),
    .D(_0971_),
    .X(_0972_));
 sky130_fd_sc_hd__o31a_1 _3784_ (.A1(_0566_),
    .A2(_0964_),
    .A3(_0972_),
    .B1(net37),
    .X(_0973_));
 sky130_fd_sc_hd__or4_1 _3785_ (.A(_1276_),
    .B(_1455_),
    .C(net73),
    .D(net27),
    .X(_0974_));
 sky130_fd_sc_hd__or3_1 _3786_ (.A(_1423_),
    .B(_1500_),
    .C(_0433_),
    .X(_0975_));
 sky130_fd_sc_hd__or4_1 _3787_ (.A(_1538_),
    .B(_1739_),
    .C(_0974_),
    .D(_0975_),
    .X(_0976_));
 sky130_fd_sc_hd__or3_1 _3788_ (.A(_1243_),
    .B(_1624_),
    .C(_0430_),
    .X(_0977_));
 sky130_fd_sc_hd__or3_1 _3789_ (.A(_0568_),
    .B(_0777_),
    .C(_0977_),
    .X(_0978_));
 sky130_fd_sc_hd__or4_1 _3790_ (.A(_0425_),
    .B(_0588_),
    .C(_0595_),
    .D(_0755_),
    .X(_0980_));
 sky130_fd_sc_hd__or4_2 _3791_ (.A(_1391_),
    .B(_1513_),
    .C(_1584_),
    .D(_1641_),
    .X(_0981_));
 sky130_fd_sc_hd__or4_1 _3792_ (.A(_1512_),
    .B(net16),
    .C(_1867_),
    .D(_0446_),
    .X(_0982_));
 sky130_fd_sc_hd__a2111o_1 _3793_ (.A1(net243),
    .A2(_1089_),
    .B1(_1222_),
    .C1(_1509_),
    .D1(_1709_),
    .X(_0983_));
 sky130_fd_sc_hd__or3b_1 _3794_ (.A(_1660_),
    .B(_1419_),
    .C_N(_1659_),
    .X(_0984_));
 sky130_fd_sc_hd__or4_1 _3795_ (.A(_0981_),
    .B(_0982_),
    .C(_0983_),
    .D(_0984_),
    .X(_0985_));
 sky130_fd_sc_hd__or3_1 _3796_ (.A(_0448_),
    .B(_0541_),
    .C(_0824_),
    .X(_0986_));
 sky130_fd_sc_hd__or4_1 _3797_ (.A(_0978_),
    .B(_0980_),
    .C(_0985_),
    .D(_0986_),
    .X(_0987_));
 sky130_fd_sc_hd__o31a_1 _3798_ (.A1(_0424_),
    .A2(_0976_),
    .A3(_0987_),
    .B1(net52),
    .X(_0988_));
 sky130_fd_sc_hd__or4_1 _3799_ (.A(_1310_),
    .B(_1447_),
    .C(_0419_),
    .D(_0421_),
    .X(_0989_));
 sky130_fd_sc_hd__or4_1 _3800_ (.A(_1410_),
    .B(_1442_),
    .C(_1643_),
    .D(_0782_),
    .X(_0991_));
 sky130_fd_sc_hd__or4_1 _3801_ (.A(_1636_),
    .B(_1716_),
    .C(_0078_),
    .D(_0373_),
    .X(_0992_));
 sky130_fd_sc_hd__or2_1 _3802_ (.A(_0633_),
    .B(_0951_),
    .X(_0993_));
 sky130_fd_sc_hd__or2_1 _3803_ (.A(_0443_),
    .B(_0991_),
    .X(_0994_));
 sky130_fd_sc_hd__or3_1 _3804_ (.A(_1548_),
    .B(_1687_),
    .C(_1739_),
    .X(_0995_));
 sky130_fd_sc_hd__a211o_1 _3805_ (.A1(_1146_),
    .A2(net89),
    .B1(_1489_),
    .C1(_1745_),
    .X(_0996_));
 sky130_fd_sc_hd__or3_1 _3806_ (.A(_1222_),
    .B(_1257_),
    .C(_1923_),
    .X(_0997_));
 sky130_fd_sc_hd__or4_1 _3807_ (.A(_0538_),
    .B(_0995_),
    .C(_0996_),
    .D(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__or4_1 _3808_ (.A(_1657_),
    .B(_1765_),
    .C(_1824_),
    .D(_0514_),
    .X(_0999_));
 sky130_fd_sc_hd__or4_1 _3809_ (.A(_0526_),
    .B(_0989_),
    .C(_0992_),
    .D(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__or4_4 _3810_ (.A(_0993_),
    .B(_0994_),
    .C(_0998_),
    .D(_1000_),
    .X(_1002_));
 sky130_fd_sc_hd__a2111o_2 _3811_ (.A1(net32),
    .A2(_1002_),
    .B1(_0167_),
    .C1(_0152_),
    .D1(_0066_),
    .X(_1003_));
 sky130_fd_sc_hd__or4_2 _3812_ (.A(_0961_),
    .B(_0973_),
    .C(_0988_),
    .D(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__or4_2 _3813_ (.A(_1377_),
    .B(_1767_),
    .C(_1868_),
    .D(net67),
    .X(_1005_));
 sky130_fd_sc_hd__or4_4 _3814_ (.A(_1803_),
    .B(_1804_),
    .C(_1860_),
    .D(_1955_),
    .X(_1006_));
 sky130_fd_sc_hd__or4_1 _3815_ (.A(_1812_),
    .B(_1814_),
    .C(_1829_),
    .D(_0280_),
    .X(_1007_));
 sky130_fd_sc_hd__or4_1 _3816_ (.A(_1651_),
    .B(_1673_),
    .C(_1755_),
    .D(_1787_),
    .X(_1008_));
 sky130_fd_sc_hd__or4_1 _3817_ (.A(_1429_),
    .B(_1436_),
    .C(_1465_),
    .D(_0086_),
    .X(_1009_));
 sky130_fd_sc_hd__a221o_1 _3818_ (.A1(net129),
    .A2(net193),
    .B1(net138),
    .B2(net119),
    .C1(net71),
    .X(_1010_));
 sky130_fd_sc_hd__a2111o_1 _3819_ (.A1(net123),
    .A2(net138),
    .B1(_1354_),
    .C1(_1494_),
    .D1(net73),
    .X(_1011_));
 sky130_fd_sc_hd__a211o_1 _3820_ (.A1(net182),
    .A2(net88),
    .B1(_1010_),
    .C1(_1011_),
    .X(_1013_));
 sky130_fd_sc_hd__or4_4 _3821_ (.A(_1007_),
    .B(_1008_),
    .C(_1009_),
    .D(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__or4_4 _3822_ (.A(_1806_),
    .B(_0206_),
    .C(_0432_),
    .D(_0702_),
    .X(_1015_));
 sky130_fd_sc_hd__or3_1 _3823_ (.A(_0480_),
    .B(_0623_),
    .C(_1005_),
    .X(_1016_));
 sky130_fd_sc_hd__or4_1 _3824_ (.A(_0584_),
    .B(_0631_),
    .C(_1015_),
    .D(_1016_),
    .X(_1017_));
 sky130_fd_sc_hd__or4_1 _3825_ (.A(_1569_),
    .B(_1570_),
    .C(_0421_),
    .D(_0453_),
    .X(_1018_));
 sky130_fd_sc_hd__or4_1 _3826_ (.A(_0478_),
    .B(_0502_),
    .C(_0632_),
    .D(_0756_),
    .X(_1019_));
 sky130_fd_sc_hd__or4_1 _3827_ (.A(_0558_),
    .B(_0586_),
    .C(_1018_),
    .D(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__a2111o_1 _3828_ (.A1(net105),
    .A2(net138),
    .B1(_1363_),
    .C1(net69),
    .D1(net94),
    .X(_1021_));
 sky130_fd_sc_hd__a2111o_4 _3829_ (.A1(net202),
    .A2(net88),
    .B1(_1525_),
    .C1(_1021_),
    .D1(_1290_),
    .X(_1022_));
 sky130_fd_sc_hd__or3_1 _3830_ (.A(_1396_),
    .B(_1458_),
    .C(_1461_),
    .X(_1024_));
 sky130_fd_sc_hd__or4_1 _3831_ (.A(_0697_),
    .B(_1006_),
    .C(_1022_),
    .D(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__or4_4 _3832_ (.A(_1014_),
    .B(_1017_),
    .C(_1020_),
    .D(_1025_),
    .X(_1026_));
 sky130_fd_sc_hd__o41a_2 _3833_ (.A1(_0427_),
    .A2(_0471_),
    .A3(_0991_),
    .A4(_1026_),
    .B1(net66),
    .X(_1027_));
 sky130_fd_sc_hd__or3_1 _3834_ (.A(_1590_),
    .B(_1983_),
    .C(_0578_),
    .X(_1028_));
 sky130_fd_sc_hd__or3_1 _3835_ (.A(net76),
    .B(_1417_),
    .C(net69),
    .X(_1029_));
 sky130_fd_sc_hd__or4_1 _3836_ (.A(_1468_),
    .B(_1637_),
    .C(_1678_),
    .D(_1782_),
    .X(_1030_));
 sky130_fd_sc_hd__or4_1 _3837_ (.A(_1661_),
    .B(_0416_),
    .C(_0644_),
    .D(_0727_),
    .X(_1031_));
 sky130_fd_sc_hd__or3_1 _3838_ (.A(_0580_),
    .B(_0609_),
    .C(_0746_),
    .X(_1032_));
 sky130_fd_sc_hd__or4_2 _3839_ (.A(_1297_),
    .B(_1812_),
    .C(_1992_),
    .D(_0527_),
    .X(_1033_));
 sky130_fd_sc_hd__o31a_1 _3840_ (.A1(net168),
    .A2(net141),
    .A3(net135),
    .B1(_1205_),
    .X(_1035_));
 sky130_fd_sc_hd__or4_1 _3841_ (.A(_1923_),
    .B(_1926_),
    .C(_1029_),
    .D(_1035_),
    .X(_1036_));
 sky130_fd_sc_hd__or4_2 _3842_ (.A(_1771_),
    .B(_0723_),
    .C(_1033_),
    .D(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__or4_1 _3843_ (.A(net70),
    .B(_1690_),
    .C(_1696_),
    .D(_1713_),
    .X(_1038_));
 sky130_fd_sc_hd__or4_1 _3844_ (.A(_1576_),
    .B(_0086_),
    .C(_1030_),
    .D(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__or4_4 _3845_ (.A(_0935_),
    .B(_1463_),
    .C(_1613_),
    .D(_1744_),
    .X(_1040_));
 sky130_fd_sc_hd__or4_1 _3846_ (.A(_1585_),
    .B(_1725_),
    .C(_1743_),
    .D(_1040_),
    .X(_1041_));
 sky130_fd_sc_hd__or4_1 _3847_ (.A(_1032_),
    .B(_1037_),
    .C(_1039_),
    .D(_1041_),
    .X(_1042_));
 sky130_fd_sc_hd__or4_1 _3848_ (.A(_0779_),
    .B(_1028_),
    .C(_1031_),
    .D(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__a2111o_2 _3849_ (.A1(_1372_),
    .A2(_1043_),
    .B1(_1027_),
    .C1(_0410_),
    .D1(_0139_),
    .X(_1044_));
 sky130_fd_sc_hd__or4_2 _3850_ (.A(_1347_),
    .B(_1428_),
    .C(_1971_),
    .D(_0629_),
    .X(_1046_));
 sky130_fd_sc_hd__or4_1 _3851_ (.A(_1346_),
    .B(_1355_),
    .C(_1682_),
    .D(_1697_),
    .X(_1047_));
 sky130_fd_sc_hd__a211o_1 _3852_ (.A1(_1294_),
    .A2(net81),
    .B1(_1494_),
    .C1(_1578_),
    .X(_1048_));
 sky130_fd_sc_hd__or4_1 _3853_ (.A(net82),
    .B(_1584_),
    .C(_1885_),
    .D(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__or4_2 _3854_ (.A(_1500_),
    .B(_1586_),
    .C(_1679_),
    .D(_1699_),
    .X(_1050_));
 sky130_fd_sc_hd__or4_4 _3855_ (.A(_0851_),
    .B(_1047_),
    .C(_1049_),
    .D(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__o31a_1 _3856_ (.A1(_0446_),
    .A2(_1046_),
    .A3(_1051_),
    .B1(net62),
    .X(_1052_));
 sky130_fd_sc_hd__or3_1 _3857_ (.A(_1895_),
    .B(_1897_),
    .C(_0178_),
    .X(_1053_));
 sky130_fd_sc_hd__or4_1 _3858_ (.A(_1319_),
    .B(_1435_),
    .C(_1568_),
    .D(_1606_),
    .X(_1054_));
 sky130_fd_sc_hd__or2_1 _3859_ (.A(_1258_),
    .B(_0782_),
    .X(_1055_));
 sky130_fd_sc_hd__or4_1 _3860_ (.A(_1350_),
    .B(_1618_),
    .C(_1054_),
    .D(_1055_),
    .X(_1057_));
 sky130_fd_sc_hd__or4_1 _3861_ (.A(_1410_),
    .B(_1641_),
    .C(_0496_),
    .D(_0896_),
    .X(_1058_));
 sky130_fd_sc_hd__or4_1 _3862_ (.A(_1280_),
    .B(_0179_),
    .C(_0474_),
    .D(_0785_),
    .X(_1059_));
 sky130_fd_sc_hd__or3_4 _3863_ (.A(_1433_),
    .B(_1519_),
    .C(_1764_),
    .X(_1060_));
 sky130_fd_sc_hd__or4_1 _3864_ (.A(_1896_),
    .B(_1058_),
    .C(_1059_),
    .D(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__o31a_1 _3865_ (.A1(_1053_),
    .A2(_1057_),
    .A3(_1061_),
    .B1(net19),
    .X(_1062_));
 sky130_fd_sc_hd__or3_2 _3866_ (.A(_1254_),
    .B(_1309_),
    .C(_1552_),
    .X(_1063_));
 sky130_fd_sc_hd__or3_1 _3867_ (.A(_1757_),
    .B(_0826_),
    .C(_1063_),
    .X(_1064_));
 sky130_fd_sc_hd__or3_1 _3868_ (.A(_1646_),
    .B(net15),
    .C(_0359_),
    .X(_1065_));
 sky130_fd_sc_hd__a22o_1 _3869_ (.A1(net155),
    .A2(net89),
    .B1(net81),
    .B2(net244),
    .X(_1066_));
 sky130_fd_sc_hd__or4_1 _3870_ (.A(_1305_),
    .B(_1921_),
    .C(_0077_),
    .D(_1066_),
    .X(_1068_));
 sky130_fd_sc_hd__or4_1 _3871_ (.A(_2014_),
    .B(_0280_),
    .C(_1065_),
    .D(_1068_),
    .X(_1069_));
 sky130_fd_sc_hd__o31a_1 _3872_ (.A1(_0661_),
    .A2(_1064_),
    .A3(_1069_),
    .B1(net31),
    .X(_1070_));
 sky130_fd_sc_hd__or4_2 _3873_ (.A(_1447_),
    .B(_1731_),
    .C(_0445_),
    .D(_0755_),
    .X(_1071_));
 sky130_fd_sc_hd__or4_1 _3874_ (.A(_0470_),
    .B(_0521_),
    .C(_0828_),
    .D(_0956_),
    .X(_1072_));
 sky130_fd_sc_hd__or4_1 _3875_ (.A(_1291_),
    .B(_1644_),
    .C(_1691_),
    .D(_2016_),
    .X(_1073_));
 sky130_fd_sc_hd__or3_1 _3876_ (.A(_1419_),
    .B(_1439_),
    .C(_1442_),
    .X(_1074_));
 sky130_fd_sc_hd__or4_1 _3877_ (.A(_1479_),
    .B(_1653_),
    .C(_1733_),
    .D(_0544_),
    .X(_1075_));
 sky130_fd_sc_hd__or4_2 _3878_ (.A(_0579_),
    .B(_1073_),
    .C(_1074_),
    .D(_1075_),
    .X(_1076_));
 sky130_fd_sc_hd__or4_1 _3879_ (.A(_1678_),
    .B(_1729_),
    .C(_0287_),
    .D(_0692_),
    .X(_1077_));
 sky130_fd_sc_hd__or3_1 _3880_ (.A(_1615_),
    .B(_1688_),
    .C(_1770_),
    .X(_1079_));
 sky130_fd_sc_hd__or3_2 _3881_ (.A(_1072_),
    .B(_1077_),
    .C(_1079_),
    .X(_1080_));
 sky130_fd_sc_hd__or4_4 _3882_ (.A(_0952_),
    .B(_1071_),
    .C(_1076_),
    .D(_1080_),
    .X(_1081_));
 sky130_fd_sc_hd__a2111o_1 _3883_ (.A1(net19),
    .A2(_1081_),
    .B1(_1070_),
    .C1(_1062_),
    .D1(_1052_),
    .X(_1082_));
 sky130_fd_sc_hd__or2_1 _3884_ (.A(_1407_),
    .B(_1418_),
    .X(_1083_));
 sky130_fd_sc_hd__or4_1 _3885_ (.A(_1274_),
    .B(_1537_),
    .C(_1550_),
    .D(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__or3_2 _3886_ (.A(_1564_),
    .B(_1610_),
    .C(_0537_),
    .X(_1085_));
 sky130_fd_sc_hd__or4_1 _3887_ (.A(_1955_),
    .B(_0086_),
    .C(_1084_),
    .D(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__or3_1 _3888_ (.A(_1767_),
    .B(net68),
    .C(_0453_),
    .X(_1087_));
 sky130_fd_sc_hd__or4_1 _3889_ (.A(_1802_),
    .B(_0497_),
    .C(_0509_),
    .D(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__or3_1 _3890_ (.A(_1526_),
    .B(_1795_),
    .C(_0435_),
    .X(_1090_));
 sky130_fd_sc_hd__or3_1 _3891_ (.A(_1514_),
    .B(_0309_),
    .C(_1090_),
    .X(_1091_));
 sky130_fd_sc_hd__or4_2 _3892_ (.A(_0524_),
    .B(_1086_),
    .C(_1088_),
    .D(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__a2111o_1 _3893_ (.A1(net55),
    .A2(_1092_),
    .B1(_0230_),
    .C1(_0090_),
    .D1(_0073_),
    .X(_1093_));
 sky130_fd_sc_hd__or4b_2 _3894_ (.A(_1420_),
    .B(_1651_),
    .C(_0522_),
    .D_N(_1659_),
    .X(_1094_));
 sky130_fd_sc_hd__or4_1 _3895_ (.A(_1366_),
    .B(_1434_),
    .C(_1576_),
    .D(_1755_),
    .X(_1095_));
 sky130_fd_sc_hd__or3_1 _3896_ (.A(_0690_),
    .B(_1071_),
    .C(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__a2111o_1 _3897_ (.A1(net129),
    .A2(net183),
    .B1(_1316_),
    .C1(_0494_),
    .D1(_0593_),
    .X(_1097_));
 sky130_fd_sc_hd__or4_2 _3898_ (.A(_1807_),
    .B(_0576_),
    .C(_1085_),
    .D(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__or4_1 _3899_ (.A(_1607_),
    .B(_1618_),
    .C(_1794_),
    .D(_0698_),
    .X(_1099_));
 sky130_fd_sc_hd__or4_2 _3900_ (.A(_0935_),
    .B(_1271_),
    .C(_1342_),
    .D(_1363_),
    .X(_1101_));
 sky130_fd_sc_hd__or4_1 _3901_ (.A(_1590_),
    .B(_1743_),
    .C(_0085_),
    .D(_0544_),
    .X(_1102_));
 sky130_fd_sc_hd__or4_1 _3902_ (.A(_1094_),
    .B(_1099_),
    .C(_1101_),
    .D(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__o31a_1 _3903_ (.A1(_1096_),
    .A2(_1098_),
    .A3(_1103_),
    .B1(net37),
    .X(_1104_));
 sky130_fd_sc_hd__or2_1 _3904_ (.A(_0504_),
    .B(_0608_),
    .X(_1105_));
 sky130_fd_sc_hd__or4_1 _3905_ (.A(_1446_),
    .B(_1835_),
    .C(_0088_),
    .D(_0786_),
    .X(_1106_));
 sky130_fd_sc_hd__or4_1 _3906_ (.A(_0589_),
    .B(_1028_),
    .C(_1105_),
    .D(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__or4b_1 _3907_ (.A(_1453_),
    .B(_0077_),
    .C(_0824_),
    .D_N(_0837_),
    .X(_1108_));
 sky130_fd_sc_hd__or4_1 _3908_ (.A(_1257_),
    .B(_1531_),
    .C(_1570_),
    .D(_1628_),
    .X(_1109_));
 sky130_fd_sc_hd__or4_1 _3909_ (.A(_1629_),
    .B(_1712_),
    .C(_0425_),
    .D(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__or3_1 _3910_ (.A(_1243_),
    .B(_1654_),
    .C(_0432_),
    .X(_1112_));
 sky130_fd_sc_hd__or4_2 _3911_ (.A(_1222_),
    .B(_1473_),
    .C(_1690_),
    .D(_1112_),
    .X(_1113_));
 sky130_fd_sc_hd__or3_1 _3912_ (.A(_1108_),
    .B(_1110_),
    .C(_1113_),
    .X(_1114_));
 sky130_fd_sc_hd__a221o_2 _3913_ (.A1(net52),
    .A2(_1107_),
    .B1(_1114_),
    .B2(net59),
    .C1(_1104_),
    .X(_1115_));
 sky130_fd_sc_hd__or4_1 _3914_ (.A(_1970_),
    .B(_1082_),
    .C(_1093_),
    .D(_1115_),
    .X(_1116_));
 sky130_fd_sc_hd__or4_4 _3915_ (.A(_0928_),
    .B(_1004_),
    .C(_1044_),
    .D(_1116_),
    .X(_1117_));
 sky130_fd_sc_hd__nor4_2 _3916_ (.A(_1780_),
    .B(_0744_),
    .C(_0800_),
    .D(_1117_),
    .Y(_0000_));
 sky130_fd_sc_hd__and3_1 _3917_ (.A(\vgatest.vcounter[3] ),
    .B(\vgatest.vcounter[2] ),
    .C(\vgatest.vcounter[0] ),
    .X(_1118_));
 sky130_fd_sc_hd__and4_4 _3918_ (.A(\vgatest.vcounter[5] ),
    .B(_0094_),
    .C(_0149_),
    .D(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__and2_1 _3919_ (.A(\vgatest.hcounter[0] ),
    .B(\vgatest.hcounter[1] ),
    .X(_1120_));
 sky130_fd_sc_hd__and3_4 _3920_ (.A(\vgatest.hcounter[0] ),
    .B(\vgatest.hcounter[1] ),
    .C(\vgatest.hcounter[2] ),
    .X(_1122_));
 sky130_fd_sc_hd__and3b_1 _3921_ (.A_N(\vgatest.hcounter[6] ),
    .B(\vgatest.hcounter[7] ),
    .C(\vgatest.hcounter[5] ),
    .X(_1123_));
 sky130_fd_sc_hd__nor2_1 _3922_ (.A(\vgatest.hcounter[3] ),
    .B(\vgatest.hcounter[4] ),
    .Y(_1124_));
 sky130_fd_sc_hd__and4b_1 _3923_ (.A_N(_0202_),
    .B(_1122_),
    .C(_1123_),
    .D(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__clkinv_2 _3924_ (.A(net275),
    .Y(_1126_));
 sky130_fd_sc_hd__and2_2 _3925_ (.A(_1119_),
    .B(net274),
    .X(_1127_));
 sky130_fd_sc_hd__and3_2 _3926_ (.A(\vgatest.framecounter[0] ),
    .B(_1119_),
    .C(net274),
    .X(_1128_));
 sky130_fd_sc_hd__nor2_1 _3927_ (.A(net277),
    .B(_1128_),
    .Y(_1129_));
 sky130_fd_sc_hd__o21a_1 _3928_ (.A1(\vgatest.framecounter[0] ),
    .A2(_1127_),
    .B1(_1129_),
    .X(_0001_));
 sky130_fd_sc_hd__and2_2 _3929_ (.A(\vgatest.framecounter[1] ),
    .B(_1128_),
    .X(_1130_));
 sky130_fd_sc_hd__nor2_1 _3930_ (.A(net277),
    .B(_1130_),
    .Y(_1132_));
 sky130_fd_sc_hd__o21a_1 _3931_ (.A1(\vgatest.framecounter[1] ),
    .A2(_1128_),
    .B1(_1132_),
    .X(_0002_));
 sky130_fd_sc_hd__a21oi_1 _3932_ (.A1(\vgatest.framecounter[2] ),
    .A2(_1130_),
    .B1(net277),
    .Y(_1133_));
 sky130_fd_sc_hd__o21a_1 _3933_ (.A1(\vgatest.framecounter[2] ),
    .A2(_1130_),
    .B1(_1133_),
    .X(_0003_));
 sky130_fd_sc_hd__a21oi_1 _3934_ (.A1(\vgatest.framecounter[2] ),
    .A2(_1130_),
    .B1(\vgatest.framecounter[3] ),
    .Y(_1134_));
 sky130_fd_sc_hd__and3_1 _3935_ (.A(\vgatest.framecounter[3] ),
    .B(\vgatest.framecounter[2] ),
    .C(_1130_),
    .X(_1135_));
 sky130_fd_sc_hd__nor3_1 _3936_ (.A(net277),
    .B(_1134_),
    .C(_1135_),
    .Y(_0004_));
 sky130_fd_sc_hd__and2_1 _3937_ (.A(\vgatest.framecounter[4] ),
    .B(_1135_),
    .X(_1136_));
 sky130_fd_sc_hd__nor2_1 _3938_ (.A(net277),
    .B(_1136_),
    .Y(_1137_));
 sky130_fd_sc_hd__o21a_1 _3939_ (.A1(\vgatest.framecounter[4] ),
    .A2(_1135_),
    .B1(_1137_),
    .X(_0005_));
 sky130_fd_sc_hd__a21oi_1 _3940_ (.A1(\vgatest.framecounter[5] ),
    .A2(_1136_),
    .B1(net277),
    .Y(_1139_));
 sky130_fd_sc_hd__o21a_1 _3941_ (.A1(\vgatest.framecounter[5] ),
    .A2(_1136_),
    .B1(_1139_),
    .X(_0006_));
 sky130_fd_sc_hd__a21oi_1 _3942_ (.A1(\vgatest.vcounter[0] ),
    .A2(net274),
    .B1(net277),
    .Y(_1140_));
 sky130_fd_sc_hd__o21a_1 _3943_ (.A1(\vgatest.vcounter[0] ),
    .A2(net274),
    .B1(_1140_),
    .X(_0007_));
 sky130_fd_sc_hd__and2_4 _3944_ (.A(\vgatest.vcounter[1] ),
    .B(\vgatest.vcounter[0] ),
    .X(_1141_));
 sky130_fd_sc_hd__nor2_4 _3945_ (.A(_1119_),
    .B(_1126_),
    .Y(_1142_));
 sky130_fd_sc_hd__or2_4 _3946_ (.A(_1119_),
    .B(_1126_),
    .X(_1143_));
 sky130_fd_sc_hd__o32a_1 _3947_ (.A1(_0138_),
    .A2(_1141_),
    .A3(_1143_),
    .B1(net275),
    .B2(_0094_),
    .X(_1144_));
 sky130_fd_sc_hd__nor2_1 _3948_ (.A(net278),
    .B(_1144_),
    .Y(_0008_));
 sky130_fd_sc_hd__nor2_1 _3949_ (.A(net277),
    .B(net274),
    .Y(_1145_));
 sky130_fd_sc_hd__or2_1 _3950_ (.A(\vgatest.vcounter[2] ),
    .B(_1141_),
    .X(_1147_));
 sky130_fd_sc_hd__and3_2 _3951_ (.A(\vgatest.vcounter[2] ),
    .B(\vgatest.vcounter[1] ),
    .C(\vgatest.vcounter[0] ),
    .X(_1148_));
 sky130_fd_sc_hd__inv_2 _3952_ (.A(_1148_),
    .Y(_1149_));
 sky130_fd_sc_hd__nor2_8 _3953_ (.A(net278),
    .B(_1143_),
    .Y(_1150_));
 sky130_fd_sc_hd__a32o_1 _3954_ (.A1(_1147_),
    .A2(_1149_),
    .A3(_1150_),
    .B1(net268),
    .B2(\vgatest.vcounter[2] ),
    .X(_0009_));
 sky130_fd_sc_hd__nor2_1 _3955_ (.A(\vgatest.vcounter[3] ),
    .B(_1148_),
    .Y(_1151_));
 sky130_fd_sc_hd__a21oi_1 _3956_ (.A1(\vgatest.vcounter[1] ),
    .A2(_1118_),
    .B1(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hd__a22o_1 _3957_ (.A1(\vgatest.vcounter[3] ),
    .A2(net269),
    .B1(_1150_),
    .B2(_1152_),
    .X(_0010_));
 sky130_fd_sc_hd__and3_2 _3958_ (.A(\vgatest.vcounter[4] ),
    .B(\vgatest.vcounter[3] ),
    .C(_1148_),
    .X(_1153_));
 sky130_fd_sc_hd__a21o_1 _3959_ (.A1(\vgatest.vcounter[3] ),
    .A2(_1148_),
    .B1(\vgatest.vcounter[4] ),
    .X(_1154_));
 sky130_fd_sc_hd__and2b_1 _3960_ (.A_N(_1153_),
    .B(_1154_),
    .X(_1156_));
 sky130_fd_sc_hd__a22o_1 _3961_ (.A1(\vgatest.vcounter[4] ),
    .A2(net269),
    .B1(_1150_),
    .B2(_1156_),
    .X(_0011_));
 sky130_fd_sc_hd__nand3_1 _3962_ (.A(\vgatest.vcounter[5] ),
    .B(net274),
    .C(_1153_),
    .Y(_1157_));
 sky130_fd_sc_hd__nor2_4 _3963_ (.A(net277),
    .B(_1127_),
    .Y(_1158_));
 sky130_fd_sc_hd__a21o_1 _3964_ (.A1(net274),
    .A2(_1153_),
    .B1(\vgatest.vcounter[5] ),
    .X(_1159_));
 sky130_fd_sc_hd__and3_1 _3965_ (.A(_1157_),
    .B(_1158_),
    .C(_1159_),
    .X(_0012_));
 sky130_fd_sc_hd__and3_1 _3966_ (.A(\vgatest.vcounter[6] ),
    .B(\vgatest.vcounter[5] ),
    .C(_1153_),
    .X(_1160_));
 sky130_fd_sc_hd__a21o_1 _3967_ (.A1(net274),
    .A2(_1160_),
    .B1(net278),
    .X(_1161_));
 sky130_fd_sc_hd__a21oi_1 _3968_ (.A1(_0083_),
    .A2(_1157_),
    .B1(_1161_),
    .Y(_0013_));
 sky130_fd_sc_hd__and2_1 _3969_ (.A(\vgatest.vcounter[7] ),
    .B(_1160_),
    .X(_1162_));
 sky130_fd_sc_hd__a21o_1 _3970_ (.A1(_1142_),
    .A2(_1160_),
    .B1(\vgatest.vcounter[7] ),
    .X(_1164_));
 sky130_fd_sc_hd__nand2_1 _3971_ (.A(net275),
    .B(_1162_),
    .Y(_1165_));
 sky130_fd_sc_hd__and3_1 _3972_ (.A(_1158_),
    .B(_1164_),
    .C(_1165_),
    .X(_0014_));
 sky130_fd_sc_hd__a21o_1 _3973_ (.A1(_1142_),
    .A2(_1162_),
    .B1(\vgatest.vcounter[8] ),
    .X(_1166_));
 sky130_fd_sc_hd__o211ai_1 _3974_ (.A1(_1143_),
    .A2(_1162_),
    .B1(\vgatest.vcounter[8] ),
    .C1(net274),
    .Y(_1167_));
 sky130_fd_sc_hd__and3_1 _3975_ (.A(_0116_),
    .B(_1166_),
    .C(_1167_),
    .X(_0015_));
 sky130_fd_sc_hd__o311a_2 _3976_ (.A1(\vgatest.vcounter[6] ),
    .A2(\vgatest.vcounter[5] ),
    .A3(\vgatest.vcounter[4] ),
    .B1(\vgatest.vcounter[7] ),
    .C1(\vgatest.vcounter[8] ),
    .X(_1168_));
 sky130_fd_sc_hd__a2111o_4 _3977_ (.A1(\vgatest.hcounter[8] ),
    .A2(\vgatest.hcounter[9] ),
    .B1(net278),
    .C1(_0191_),
    .D1(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__mux4_2 _3978_ (.A0(\vgatest.bitmap.res[0] ),
    .A1(\vgatest.bitmap.res[1] ),
    .A2(\vgatest.bitmap.res[2] ),
    .A3(\vgatest.bitmap.res[3] ),
    .S0(\vgatest.hcounter[2] ),
    .S1(\vgatest.hcounter[3] ),
    .X(_1170_));
 sky130_fd_sc_hd__nand2_4 _3979_ (.A(_0127_),
    .B(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__o21ai_1 _3980_ (.A1(\vgatest.framecounter[2] ),
    .A2(\vgatest.hcounter[0] ),
    .B1(net1),
    .Y(_1173_));
 sky130_fd_sc_hd__a21o_1 _3981_ (.A1(\vgatest.framecounter[2] ),
    .A2(\vgatest.hcounter[0] ),
    .B1(_1173_),
    .X(_1174_));
 sky130_fd_sc_hd__a21oi_1 _3982_ (.A1(_1171_),
    .A2(_1174_),
    .B1(_1169_),
    .Y(_0016_));
 sky130_fd_sc_hd__nand2_2 _3983_ (.A(\vgatest.framecounter[3] ),
    .B(\vgatest.hcounter[1] ),
    .Y(_1175_));
 sky130_fd_sc_hd__or2_1 _3984_ (.A(\vgatest.framecounter[3] ),
    .B(\vgatest.hcounter[1] ),
    .X(_1176_));
 sky130_fd_sc_hd__and2_2 _3985_ (.A(_1175_),
    .B(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__a21oi_1 _3986_ (.A1(\vgatest.framecounter[2] ),
    .A2(\vgatest.hcounter[0] ),
    .B1(_1177_),
    .Y(_1178_));
 sky130_fd_sc_hd__nand3_4 _3987_ (.A(\vgatest.framecounter[2] ),
    .B(\vgatest.hcounter[0] ),
    .C(_1177_),
    .Y(_1179_));
 sky130_fd_sc_hd__or3b_1 _3988_ (.A(_0127_),
    .B(_1178_),
    .C_N(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__a21oi_1 _3989_ (.A1(_1171_),
    .A2(_1180_),
    .B1(_1169_),
    .Y(_0017_));
 sky130_fd_sc_hd__and2_2 _3990_ (.A(\vgatest.framecounter[4] ),
    .B(\vgatest.hcounter[2] ),
    .X(_1182_));
 sky130_fd_sc_hd__nor2_2 _3991_ (.A(\vgatest.framecounter[4] ),
    .B(\vgatest.hcounter[2] ),
    .Y(_1183_));
 sky130_fd_sc_hd__a211oi_4 _3992_ (.A1(_1175_),
    .A2(_1179_),
    .B1(_1182_),
    .C1(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hd__o211a_1 _3993_ (.A1(_1182_),
    .A2(_1183_),
    .B1(_1175_),
    .C1(_1179_),
    .X(_1185_));
 sky130_fd_sc_hd__o31a_1 _3994_ (.A1(_0127_),
    .A2(_1184_),
    .A3(_1185_),
    .B1(_1171_),
    .X(_1186_));
 sky130_fd_sc_hd__nor2_1 _3995_ (.A(_1169_),
    .B(_1186_),
    .Y(_0018_));
 sky130_fd_sc_hd__xor2_2 _3996_ (.A(\vgatest.framecounter[5] ),
    .B(\vgatest.hcounter[3] ),
    .X(_1187_));
 sky130_fd_sc_hd__nor3_1 _3997_ (.A(_1182_),
    .B(_1184_),
    .C(_1187_),
    .Y(_1188_));
 sky130_fd_sc_hd__o21a_1 _3998_ (.A1(_1182_),
    .A2(_1184_),
    .B1(_1187_),
    .X(_1189_));
 sky130_fd_sc_hd__o31a_1 _3999_ (.A1(_0127_),
    .A2(_1188_),
    .A3(_1189_),
    .B1(_1171_),
    .X(_1190_));
 sky130_fd_sc_hd__nor2_1 _4000_ (.A(_1169_),
    .B(_1190_),
    .Y(_0019_));
 sky130_fd_sc_hd__nand2_1 _4001_ (.A(\vgatest.vcounter[0] ),
    .B(net1),
    .Y(_1192_));
 sky130_fd_sc_hd__a21oi_1 _4002_ (.A1(_1171_),
    .A2(_1192_),
    .B1(_1169_),
    .Y(_0020_));
 sky130_fd_sc_hd__nand2_1 _4003_ (.A(\vgatest.vcounter[1] ),
    .B(net1),
    .Y(_1193_));
 sky130_fd_sc_hd__a21oi_1 _4004_ (.A1(_1171_),
    .A2(_1193_),
    .B1(_1169_),
    .Y(_0021_));
 sky130_fd_sc_hd__nand2_1 _4005_ (.A(\vgatest.vcounter[2] ),
    .B(net1),
    .Y(_1194_));
 sky130_fd_sc_hd__a21oi_1 _4006_ (.A1(_1171_),
    .A2(_1194_),
    .B1(_1169_),
    .Y(_0022_));
 sky130_fd_sc_hd__nand2_1 _4007_ (.A(\vgatest.vcounter[3] ),
    .B(net1),
    .Y(_1195_));
 sky130_fd_sc_hd__a21oi_1 _4008_ (.A1(_1171_),
    .A2(_1195_),
    .B1(_1169_),
    .Y(_0023_));
 sky130_fd_sc_hd__and3_2 _4009_ (.A(\vgatest.bitmapColAddr[2] ),
    .B(\vgatest.vcounter[1] ),
    .C(\vgatest.vcounter[0] ),
    .X(_1196_));
 sky130_fd_sc_hd__a2bb2o_1 _4010_ (.A1_N(_1196_),
    .A2_N(_1143_),
    .B1(_1126_),
    .B2(\vgatest.bitmapColAddr[2] ),
    .X(_1198_));
 sky130_fd_sc_hd__o211a_1 _4011_ (.A1(\vgatest.bitmapColAddr[2] ),
    .A2(_1141_),
    .B1(_1198_),
    .C1(_0116_),
    .X(_0024_));
 sky130_fd_sc_hd__nand2_1 _4012_ (.A(\vgatest.bitmapColAddr[3] ),
    .B(_1196_),
    .Y(_1199_));
 sky130_fd_sc_hd__or2_1 _4013_ (.A(\vgatest.bitmapColAddr[3] ),
    .B(_1196_),
    .X(_1200_));
 sky130_fd_sc_hd__a32o_1 _4014_ (.A1(_1150_),
    .A2(_1199_),
    .A3(_1200_),
    .B1(net268),
    .B2(\vgatest.bitmapColAddr[3] ),
    .X(_0025_));
 sky130_fd_sc_hd__nand4_1 _4015_ (.A(\vgatest.bitmapColAddr[4] ),
    .B(net275),
    .C(_1141_),
    .D(_1199_),
    .Y(_1201_));
 sky130_fd_sc_hd__a31o_1 _4016_ (.A1(net275),
    .A2(_1141_),
    .A3(_1199_),
    .B1(\vgatest.bitmapColAddr[4] ),
    .X(_1202_));
 sky130_fd_sc_hd__and3_1 _4017_ (.A(_1158_),
    .B(_1201_),
    .C(_1202_),
    .X(_0026_));
 sky130_fd_sc_hd__a22o_2 _4018_ (.A1(\vgatest.bitmapColAddr[4] ),
    .A2(_1141_),
    .B1(_1196_),
    .B2(\vgatest.bitmapColAddr[3] ),
    .X(_1203_));
 sky130_fd_sc_hd__and3_1 _4019_ (.A(\vgatest.bitmapColAddr[5] ),
    .B(\vgatest.vcounter[1] ),
    .C(\vgatest.vcounter[0] ),
    .X(_1204_));
 sky130_fd_sc_hd__nor2_1 _4020_ (.A(\vgatest.bitmapColAddr[5] ),
    .B(_1141_),
    .Y(_1206_));
 sky130_fd_sc_hd__or2_1 _4021_ (.A(_1204_),
    .B(_1206_),
    .X(_1207_));
 sky130_fd_sc_hd__xnor2_1 _4022_ (.A(_1203_),
    .B(_1207_),
    .Y(_1208_));
 sky130_fd_sc_hd__a22o_1 _4023_ (.A1(\vgatest.bitmapColAddr[5] ),
    .A2(net269),
    .B1(_1150_),
    .B2(_1208_),
    .X(_0027_));
 sky130_fd_sc_hd__o21a_1 _4024_ (.A1(_1203_),
    .A2(_1204_),
    .B1(\vgatest.bitmapColAddr[6] ),
    .X(_1209_));
 sky130_fd_sc_hd__o31ai_1 _4025_ (.A1(\vgatest.bitmapColAddr[6] ),
    .A2(_1203_),
    .A3(_1204_),
    .B1(_1150_),
    .Y(_1210_));
 sky130_fd_sc_hd__a2bb2o_1 _4026_ (.A1_N(_1209_),
    .A2_N(_1210_),
    .B1(\vgatest.bitmapColAddr[6] ),
    .B2(net268),
    .X(_0028_));
 sky130_fd_sc_hd__xnor2_1 _4027_ (.A(\vgatest.bitmapColAddr[7] ),
    .B(_1141_),
    .Y(_1211_));
 sky130_fd_sc_hd__xnor2_1 _4028_ (.A(_1209_),
    .B(_1211_),
    .Y(_1212_));
 sky130_fd_sc_hd__a22o_1 _4029_ (.A1(\vgatest.bitmapColAddr[7] ),
    .A2(net268),
    .B1(_1150_),
    .B2(_1212_),
    .X(_0029_));
 sky130_fd_sc_hd__a21o_2 _4030_ (.A1(\vgatest.bitmapColAddr[7] ),
    .A2(_1141_),
    .B1(_1209_),
    .X(_1214_));
 sky130_fd_sc_hd__and2_1 _4031_ (.A(\vgatest.bitmapColAddr[8] ),
    .B(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__nor2_1 _4032_ (.A(_1143_),
    .B(_1215_),
    .Y(_1216_));
 sky130_fd_sc_hd__a21o_1 _4033_ (.A1(_1142_),
    .A2(_1214_),
    .B1(\vgatest.bitmapColAddr[8] ),
    .X(_1217_));
 sky130_fd_sc_hd__nand2_1 _4034_ (.A(net275),
    .B(_1215_),
    .Y(_1218_));
 sky130_fd_sc_hd__and3_1 _4035_ (.A(_1158_),
    .B(_1217_),
    .C(_1218_),
    .X(_0030_));
 sky130_fd_sc_hd__a31o_1 _4036_ (.A1(\vgatest.bitmapColAddr[8] ),
    .A2(_1142_),
    .A3(_1214_),
    .B1(\vgatest.bitmapColAddr[9] ),
    .X(_1219_));
 sky130_fd_sc_hd__o311a_1 _4037_ (.A1(_0072_),
    .A2(_1126_),
    .A3(_1216_),
    .B1(_1219_),
    .C1(_0116_),
    .X(_0031_));
 sky130_fd_sc_hd__and3_2 _4038_ (.A(\vgatest.bitmapColAddr[10] ),
    .B(\vgatest.bitmapColAddr[9] ),
    .C(_1215_),
    .X(_1220_));
 sky130_fd_sc_hd__inv_2 _4039_ (.A(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__a31o_1 _4040_ (.A1(\vgatest.bitmapColAddr[9] ),
    .A2(\vgatest.bitmapColAddr[8] ),
    .A3(_1214_),
    .B1(\vgatest.bitmapColAddr[10] ),
    .X(_1223_));
 sky130_fd_sc_hd__a32o_1 _4041_ (.A1(_1150_),
    .A2(_1221_),
    .A3(_1223_),
    .B1(net268),
    .B2(\vgatest.bitmapColAddr[10] ),
    .X(_0032_));
 sky130_fd_sc_hd__nand2_1 _4042_ (.A(net276),
    .B(net269),
    .Y(_1224_));
 sky130_fd_sc_hd__and2_2 _4043_ (.A(net276),
    .B(_1220_),
    .X(_1225_));
 sky130_fd_sc_hd__o21ai_1 _4044_ (.A1(\vgatest.bitmapColAddr[11] ),
    .A2(_1220_),
    .B1(_1150_),
    .Y(_1226_));
 sky130_fd_sc_hd__o21ai_1 _4045_ (.A1(_1225_),
    .A2(_1226_),
    .B1(_1224_),
    .Y(_0033_));
 sky130_fd_sc_hd__nand2_1 _4046_ (.A(\vgatest.bitmapColAddr[12] ),
    .B(_1225_),
    .Y(_1227_));
 sky130_fd_sc_hd__or2_1 _4047_ (.A(\vgatest.bitmapColAddr[12] ),
    .B(_1225_),
    .X(_1228_));
 sky130_fd_sc_hd__a32o_1 _4048_ (.A1(_1150_),
    .A2(_1227_),
    .A3(_1228_),
    .B1(net269),
    .B2(\vgatest.bitmapColAddr[12] ),
    .X(_0034_));
 sky130_fd_sc_hd__nor2_1 _4049_ (.A(_2037_),
    .B(_1227_),
    .Y(_1229_));
 sky130_fd_sc_hd__a31o_1 _4050_ (.A1(\vgatest.bitmapColAddr[12] ),
    .A2(_1142_),
    .A3(_1225_),
    .B1(\vgatest.bitmapColAddr[13] ),
    .X(_1231_));
 sky130_fd_sc_hd__nand2_1 _4051_ (.A(_1142_),
    .B(_1229_),
    .Y(_1232_));
 sky130_fd_sc_hd__and3_1 _4052_ (.A(_1158_),
    .B(_1231_),
    .C(_1232_),
    .X(_0035_));
 sky130_fd_sc_hd__o211a_1 _4053_ (.A1(_1143_),
    .A2(_1229_),
    .B1(\vgatest.bitmapColAddr[14] ),
    .C1(net274),
    .X(_1233_));
 sky130_fd_sc_hd__a211oi_1 _4054_ (.A1(_2026_),
    .A2(_1232_),
    .B1(_1233_),
    .C1(net277),
    .Y(_0036_));
 sky130_fd_sc_hd__nor2_1 _4055_ (.A(\vgatest.hcounter[0] ),
    .B(net278),
    .Y(_0037_));
 sky130_fd_sc_hd__o21ai_1 _4056_ (.A1(\vgatest.hcounter[0] ),
    .A2(\vgatest.hcounter[1] ),
    .B1(net269),
    .Y(_1234_));
 sky130_fd_sc_hd__nor2_1 _4057_ (.A(_1120_),
    .B(_1234_),
    .Y(_0038_));
 sky130_fd_sc_hd__nor2_1 _4058_ (.A(net278),
    .B(_1122_),
    .Y(_1235_));
 sky130_fd_sc_hd__o21a_1 _4059_ (.A1(\vgatest.hcounter[2] ),
    .A2(_1120_),
    .B1(_1235_),
    .X(_0039_));
 sky130_fd_sc_hd__o21ai_1 _4060_ (.A1(\vgatest.hcounter[3] ),
    .A2(_1122_),
    .B1(net269),
    .Y(_1237_));
 sky130_fd_sc_hd__a21oi_1 _4061_ (.A1(\vgatest.hcounter[3] ),
    .A2(_1122_),
    .B1(_1237_),
    .Y(_0040_));
 sky130_fd_sc_hd__nand3_1 _4062_ (.A(\vgatest.hcounter[3] ),
    .B(\vgatest.hcounter[4] ),
    .C(_1122_),
    .Y(_1238_));
 sky130_fd_sc_hd__a21o_1 _4063_ (.A1(\vgatest.hcounter[3] ),
    .A2(_1122_),
    .B1(\vgatest.hcounter[4] ),
    .X(_1239_));
 sky130_fd_sc_hd__and3_1 _4064_ (.A(net268),
    .B(_1238_),
    .C(_1239_),
    .X(_0041_));
 sky130_fd_sc_hd__and4_2 _4065_ (.A(\vgatest.hcounter[3] ),
    .B(\vgatest.hcounter[4] ),
    .C(\vgatest.hcounter[5] ),
    .D(_1122_),
    .X(_1240_));
 sky130_fd_sc_hd__a2111oi_1 _4066_ (.A1(_0105_),
    .A2(_1238_),
    .B1(_1240_),
    .C1(net278),
    .D1(net275),
    .Y(_0042_));
 sky130_fd_sc_hd__and2_1 _4067_ (.A(\vgatest.hcounter[6] ),
    .B(_1240_),
    .X(_1241_));
 sky130_fd_sc_hd__o21ai_1 _4068_ (.A1(\vgatest.hcounter[6] ),
    .A2(_1240_),
    .B1(net268),
    .Y(_1242_));
 sky130_fd_sc_hd__nor2_1 _4069_ (.A(_1241_),
    .B(_1242_),
    .Y(_0043_));
 sky130_fd_sc_hd__and3_1 _4070_ (.A(\vgatest.hcounter[6] ),
    .B(\vgatest.hcounter[7] ),
    .C(_1240_),
    .X(_1244_));
 sky130_fd_sc_hd__o21ai_1 _4071_ (.A1(\vgatest.hcounter[7] ),
    .A2(_1241_),
    .B1(net268),
    .Y(_1245_));
 sky130_fd_sc_hd__nor2_1 _4072_ (.A(_1244_),
    .B(_1245_),
    .Y(_0044_));
 sky130_fd_sc_hd__and2_1 _4073_ (.A(\vgatest.hcounter[8] ),
    .B(_1244_),
    .X(_1246_));
 sky130_fd_sc_hd__o21ai_1 _4074_ (.A1(\vgatest.hcounter[8] ),
    .A2(_1244_),
    .B1(net268),
    .Y(_1247_));
 sky130_fd_sc_hd__nor2_1 _4075_ (.A(_1246_),
    .B(_1247_),
    .Y(_0045_));
 sky130_fd_sc_hd__a21boi_1 _4076_ (.A1(\vgatest.hcounter[9] ),
    .A2(_1246_),
    .B1_N(net268),
    .Y(_1248_));
 sky130_fd_sc_hd__o21a_1 _4077_ (.A1(\vgatest.hcounter[9] ),
    .A2(_1246_),
    .B1(_1248_),
    .X(_0046_));
 sky130_fd_sc_hd__dlxtn_1 _4078_ (.D(_0047_),
    .GATE_N(_0000_),
    .Q(\vgatest.bitmap.res[0] ));
 sky130_fd_sc_hd__dlxtn_1 _4079_ (.D(_0048_),
    .GATE_N(_0000_),
    .Q(\vgatest.bitmap.res[1] ));
 sky130_fd_sc_hd__dlxtn_1 _4080_ (.D(_0049_),
    .GATE_N(_0000_),
    .Q(\vgatest.bitmap.res[2] ));
 sky130_fd_sc_hd__dlxtn_1 _4081_ (.D(_0050_),
    .GATE_N(_0000_),
    .Q(\vgatest.bitmap.res[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4082_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0001_),
    .Q(\vgatest.framecounter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4083_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0002_),
    .Q(\vgatest.framecounter[1] ));
 sky130_fd_sc_hd__dfxtp_4 _4084_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0003_),
    .Q(\vgatest.framecounter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4085_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0004_),
    .Q(\vgatest.framecounter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4086_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0005_),
    .Q(\vgatest.framecounter[4] ));
 sky130_fd_sc_hd__dfxtp_2 _4087_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0006_),
    .Q(\vgatest.framecounter[5] ));
 sky130_fd_sc_hd__dfxtp_4 _4088_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0007_),
    .Q(\vgatest.vcounter[0] ));
 sky130_fd_sc_hd__dfxtp_4 _4089_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0008_),
    .Q(\vgatest.vcounter[1] ));
 sky130_fd_sc_hd__dfxtp_2 _4090_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0009_),
    .Q(\vgatest.vcounter[2] ));
 sky130_fd_sc_hd__dfxtp_2 _4091_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0010_),
    .Q(\vgatest.vcounter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4092_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0011_),
    .Q(\vgatest.vcounter[4] ));
 sky130_fd_sc_hd__dfxtp_2 _4093_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0012_),
    .Q(\vgatest.vcounter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4094_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0013_),
    .Q(\vgatest.vcounter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4095_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0014_),
    .Q(\vgatest.vcounter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4096_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0015_),
    .Q(\vgatest.vcounter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4097_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0016_),
    .Q(net3));
 sky130_fd_sc_hd__dfxtp_1 _4098_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0017_),
    .Q(net4));
 sky130_fd_sc_hd__dfxtp_1 _4099_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0018_),
    .Q(net5));
 sky130_fd_sc_hd__dfxtp_1 _4100_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0019_),
    .Q(net6));
 sky130_fd_sc_hd__dfxtp_1 _4101_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0020_),
    .Q(net7));
 sky130_fd_sc_hd__dfxtp_1 _4102_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0021_),
    .Q(net8));
 sky130_fd_sc_hd__dfxtp_1 _4103_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0022_),
    .Q(net9));
 sky130_fd_sc_hd__dfxtp_1 _4104_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0023_),
    .Q(net10));
 sky130_fd_sc_hd__dfxtp_4 _4105_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0024_),
    .Q(\vgatest.bitmapColAddr[2] ));
 sky130_fd_sc_hd__dfxtp_4 _4106_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0025_),
    .Q(\vgatest.bitmapColAddr[3] ));
 sky130_fd_sc_hd__dfxtp_4 _4107_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0026_),
    .Q(\vgatest.bitmapColAddr[4] ));
 sky130_fd_sc_hd__dfxtp_4 _4108_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0027_),
    .Q(\vgatest.bitmapColAddr[5] ));
 sky130_fd_sc_hd__dfxtp_4 _4109_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0028_),
    .Q(\vgatest.bitmapColAddr[6] ));
 sky130_fd_sc_hd__dfxtp_4 _4110_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0029_),
    .Q(\vgatest.bitmapColAddr[7] ));
 sky130_fd_sc_hd__dfxtp_4 _4111_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0030_),
    .Q(\vgatest.bitmapColAddr[8] ));
 sky130_fd_sc_hd__dfxtp_4 _4112_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0031_),
    .Q(\vgatest.bitmapColAddr[9] ));
 sky130_fd_sc_hd__dfxtp_4 _4113_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0032_),
    .Q(\vgatest.bitmapColAddr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4114_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0033_),
    .Q(\vgatest.bitmapColAddr[11] ));
 sky130_fd_sc_hd__dfxtp_4 _4115_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0034_),
    .Q(\vgatest.bitmapColAddr[12] ));
 sky130_fd_sc_hd__dfxtp_2 _4116_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0035_),
    .Q(\vgatest.bitmapColAddr[13] ));
 sky130_fd_sc_hd__dfxtp_4 _4117_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0036_),
    .Q(\vgatest.bitmapColAddr[14] ));
 sky130_fd_sc_hd__dfxtp_4 _4118_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0037_),
    .Q(\vgatest.hcounter[0] ));
 sky130_fd_sc_hd__dfxtp_2 _4119_ (.CLK(clknet_2_1__leaf_clk),
    .D(_0038_),
    .Q(\vgatest.hcounter[1] ));
 sky130_fd_sc_hd__dfxtp_4 _4120_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0039_),
    .Q(\vgatest.hcounter[2] ));
 sky130_fd_sc_hd__dfxtp_4 _4121_ (.CLK(clknet_2_0__leaf_clk),
    .D(_0040_),
    .Q(\vgatest.hcounter[3] ));
 sky130_fd_sc_hd__dfxtp_4 _4122_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0041_),
    .Q(\vgatest.hcounter[4] ));
 sky130_fd_sc_hd__dfxtp_4 _4123_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0042_),
    .Q(\vgatest.hcounter[5] ));
 sky130_fd_sc_hd__dfxtp_4 _4124_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0043_),
    .Q(\vgatest.hcounter[6] ));
 sky130_fd_sc_hd__dfxtp_4 _4125_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0044_),
    .Q(\vgatest.hcounter[7] ));
 sky130_fd_sc_hd__dfxtp_4 _4126_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0045_),
    .Q(\vgatest.hcounter[8] ));
 sky130_fd_sc_hd__dfxtp_4 _4127_ (.CLK(clknet_2_2__leaf_clk),
    .D(_0046_),
    .Q(\vgatest.hcounter[9] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__buf_12 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__buf_12 fanout101 (.A(_1256_),
    .X(net101));
 sky130_fd_sc_hd__buf_12 fanout102 (.A(_1253_),
    .X(net102));
 sky130_fd_sc_hd__buf_12 fanout103 (.A(net104),
    .X(net103));
 sky130_fd_sc_hd__buf_12 fanout104 (.A(_1253_),
    .X(net104));
 sky130_fd_sc_hd__buf_12 fanout105 (.A(_1252_),
    .X(net105));
 sky130_fd_sc_hd__buf_12 fanout106 (.A(net108),
    .X(net106));
 sky130_fd_sc_hd__buf_12 fanout107 (.A(_1251_),
    .X(net107));
 sky130_fd_sc_hd__buf_6 fanout108 (.A(_1251_),
    .X(net108));
 sky130_fd_sc_hd__buf_12 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__buf_12 fanout110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__buf_12 fanout111 (.A(_1213_),
    .X(net111));
 sky130_fd_sc_hd__buf_12 fanout112 (.A(_1205_),
    .X(net112));
 sky130_fd_sc_hd__buf_12 fanout113 (.A(net115),
    .X(net113));
 sky130_fd_sc_hd__buf_12 fanout114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__buf_12 fanout115 (.A(_1155_),
    .X(net115));
 sky130_fd_sc_hd__buf_12 fanout116 (.A(net118),
    .X(net116));
 sky130_fd_sc_hd__buf_12 fanout117 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__buf_12 fanout118 (.A(_1100_),
    .X(net118));
 sky130_fd_sc_hd__buf_8 fanout119 (.A(net120),
    .X(net119));
 sky130_fd_sc_hd__buf_12 fanout120 (.A(_1089_),
    .X(net120));
 sky130_fd_sc_hd__buf_12 fanout121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__buf_12 fanout122 (.A(_1023_),
    .X(net122));
 sky130_fd_sc_hd__buf_8 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__buf_12 fanout124 (.A(_1012_),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_16 fanout125 (.A(_1012_),
    .X(net125));
 sky130_fd_sc_hd__buf_12 fanout126 (.A(net128),
    .X(net126));
 sky130_fd_sc_hd__buf_12 fanout127 (.A(net128),
    .X(net127));
 sky130_fd_sc_hd__buf_12 fanout128 (.A(_0924_),
    .X(net128));
 sky130_fd_sc_hd__buf_12 fanout129 (.A(_0913_),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_16 fanout13 (.A(_1926_),
    .X(net13));
 sky130_fd_sc_hd__buf_12 fanout130 (.A(_1330_),
    .X(net130));
 sky130_fd_sc_hd__buf_6 fanout131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__buf_12 fanout132 (.A(_1330_),
    .X(net132));
 sky130_fd_sc_hd__buf_8 fanout133 (.A(_1329_),
    .X(net133));
 sky130_fd_sc_hd__buf_6 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__buf_6 fanout135 (.A(_1329_),
    .X(net135));
 sky130_fd_sc_hd__buf_12 fanout136 (.A(net137),
    .X(net136));
 sky130_fd_sc_hd__buf_12 fanout137 (.A(_1327_),
    .X(net137));
 sky130_fd_sc_hd__buf_8 fanout138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_16 fanout139 (.A(_1326_),
    .X(net139));
 sky130_fd_sc_hd__buf_8 fanout14 (.A(_1824_),
    .X(net14));
 sky130_fd_sc_hd__buf_8 fanout140 (.A(net141),
    .X(net140));
 sky130_fd_sc_hd__buf_6 fanout141 (.A(_1326_),
    .X(net141));
 sky130_fd_sc_hd__buf_12 fanout142 (.A(_1307_),
    .X(net142));
 sky130_fd_sc_hd__buf_12 fanout143 (.A(_1307_),
    .X(net143));
 sky130_fd_sc_hd__buf_12 fanout144 (.A(net147),
    .X(net144));
 sky130_fd_sc_hd__buf_4 fanout145 (.A(net147),
    .X(net145));
 sky130_fd_sc_hd__buf_12 fanout146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__buf_12 fanout147 (.A(_1306_),
    .X(net147));
 sky130_fd_sc_hd__buf_12 fanout148 (.A(net149),
    .X(net148));
 sky130_fd_sc_hd__buf_12 fanout149 (.A(_1303_),
    .X(net149));
 sky130_fd_sc_hd__buf_12 fanout15 (.A(_1733_),
    .X(net15));
 sky130_fd_sc_hd__buf_12 fanout150 (.A(_1303_),
    .X(net150));
 sky130_fd_sc_hd__buf_6 fanout151 (.A(net153),
    .X(net151));
 sky130_fd_sc_hd__buf_12 fanout152 (.A(net153),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_16 fanout153 (.A(_1302_),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_16 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__buf_12 fanout155 (.A(_1294_),
    .X(net155));
 sky130_fd_sc_hd__buf_4 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__buf_4 fanout157 (.A(net161),
    .X(net157));
 sky130_fd_sc_hd__buf_4 fanout158 (.A(net160),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 fanout159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__buf_12 fanout16 (.A(_1657_),
    .X(net16));
 sky130_fd_sc_hd__buf_2 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_4 fanout161 (.A(net164),
    .X(net161));
 sky130_fd_sc_hd__buf_4 fanout162 (.A(net164),
    .X(net162));
 sky130_fd_sc_hd__buf_6 fanout163 (.A(net164),
    .X(net163));
 sky130_fd_sc_hd__buf_12 fanout164 (.A(_1286_),
    .X(net164));
 sky130_fd_sc_hd__buf_12 fanout165 (.A(_1278_),
    .X(net165));
 sky130_fd_sc_hd__buf_12 fanout166 (.A(net167),
    .X(net166));
 sky130_fd_sc_hd__buf_12 fanout167 (.A(_1278_),
    .X(net167));
 sky130_fd_sc_hd__buf_6 fanout168 (.A(_1277_),
    .X(net168));
 sky130_fd_sc_hd__buf_8 fanout169 (.A(_1277_),
    .X(net169));
 sky130_fd_sc_hd__buf_6 fanout17 (.A(_1605_),
    .X(net17));
 sky130_fd_sc_hd__buf_12 fanout170 (.A(net171),
    .X(net170));
 sky130_fd_sc_hd__buf_12 fanout171 (.A(_1270_),
    .X(net171));
 sky130_fd_sc_hd__buf_6 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__buf_12 fanout173 (.A(_1269_),
    .X(net173));
 sky130_fd_sc_hd__buf_12 fanout174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__buf_12 fanout175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__buf_12 fanout176 (.A(_1266_),
    .X(net176));
 sky130_fd_sc_hd__buf_8 fanout177 (.A(_1265_),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_4 fanout178 (.A(net179),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_16 fanout179 (.A(_1265_),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_4 fanout18 (.A(_1605_),
    .X(net18));
 sky130_fd_sc_hd__buf_8 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__buf_12 fanout181 (.A(_1255_),
    .X(net181));
 sky130_fd_sc_hd__buf_6 fanout182 (.A(net183),
    .X(net182));
 sky130_fd_sc_hd__buf_12 fanout183 (.A(net184),
    .X(net183));
 sky130_fd_sc_hd__buf_12 fanout184 (.A(_1250_),
    .X(net184));
 sky130_fd_sc_hd__buf_12 fanout185 (.A(net186),
    .X(net185));
 sky130_fd_sc_hd__buf_12 fanout186 (.A(_1236_),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_16 fanout187 (.A(net189),
    .X(net187));
 sky130_fd_sc_hd__buf_4 fanout188 (.A(net189),
    .X(net188));
 sky130_fd_sc_hd__buf_12 fanout189 (.A(_1230_),
    .X(net189));
 sky130_fd_sc_hd__buf_6 fanout19 (.A(_1605_),
    .X(net19));
 sky130_fd_sc_hd__buf_12 fanout190 (.A(net192),
    .X(net190));
 sky130_fd_sc_hd__buf_12 fanout191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__buf_12 fanout192 (.A(_1197_),
    .X(net192));
 sky130_fd_sc_hd__buf_6 fanout193 (.A(net195),
    .X(net193));
 sky130_fd_sc_hd__buf_8 fanout194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__buf_12 fanout195 (.A(_1191_),
    .X(net195));
 sky130_fd_sc_hd__buf_8 fanout196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__buf_12 fanout197 (.A(net198),
    .X(net197));
 sky130_fd_sc_hd__buf_12 fanout198 (.A(_1146_),
    .X(net198));
 sky130_fd_sc_hd__buf_12 fanout199 (.A(_1078_),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_4 fanout20 (.A(_1605_),
    .X(net20));
 sky130_fd_sc_hd__buf_12 fanout200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__buf_12 fanout201 (.A(_1078_),
    .X(net201));
 sky130_fd_sc_hd__buf_8 fanout202 (.A(_1067_),
    .X(net202));
 sky130_fd_sc_hd__buf_4 fanout203 (.A(_1067_),
    .X(net203));
 sky130_fd_sc_hd__buf_8 fanout204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__buf_6 fanout205 (.A(_1067_),
    .X(net205));
 sky130_fd_sc_hd__buf_12 fanout206 (.A(net208),
    .X(net206));
 sky130_fd_sc_hd__buf_12 fanout207 (.A(net208),
    .X(net207));
 sky130_fd_sc_hd__buf_12 fanout208 (.A(_1001_),
    .X(net208));
 sky130_fd_sc_hd__buf_6 fanout209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_16 fanout21 (.A(net23),
    .X(net21));
 sky130_fd_sc_hd__buf_6 fanout210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__buf_12 fanout211 (.A(_0990_),
    .X(net211));
 sky130_fd_sc_hd__buf_4 fanout212 (.A(net215),
    .X(net212));
 sky130_fd_sc_hd__buf_4 fanout213 (.A(net215),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 fanout214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__buf_4 fanout215 (.A(net218),
    .X(net215));
 sky130_fd_sc_hd__buf_4 fanout216 (.A(net217),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_8 fanout217 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__buf_4 fanout218 (.A(net219),
    .X(net218));
 sky130_fd_sc_hd__buf_8 fanout219 (.A(_0946_),
    .X(net219));
 sky130_fd_sc_hd__buf_8 fanout22 (.A(net23),
    .X(net22));
 sky130_fd_sc_hd__buf_6 fanout220 (.A(_0946_),
    .X(net220));
 sky130_fd_sc_hd__buf_4 fanout221 (.A(net222),
    .X(net221));
 sky130_fd_sc_hd__buf_4 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_8 fanout223 (.A(net225),
    .X(net223));
 sky130_fd_sc_hd__buf_4 fanout224 (.A(net225),
    .X(net224));
 sky130_fd_sc_hd__buf_4 fanout225 (.A(net226),
    .X(net225));
 sky130_fd_sc_hd__buf_8 fanout226 (.A(net229),
    .X(net226));
 sky130_fd_sc_hd__buf_6 fanout227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__buf_8 fanout228 (.A(net229),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_8 fanout229 (.A(_0902_),
    .X(net229));
 sky130_fd_sc_hd__buf_12 fanout23 (.A(_1588_),
    .X(net23));
 sky130_fd_sc_hd__buf_4 fanout230 (.A(net231),
    .X(net230));
 sky130_fd_sc_hd__buf_4 fanout231 (.A(net235),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_8 fanout232 (.A(net235),
    .X(net232));
 sky130_fd_sc_hd__buf_4 fanout233 (.A(net234),
    .X(net233));
 sky130_fd_sc_hd__buf_2 fanout234 (.A(net235),
    .X(net234));
 sky130_fd_sc_hd__buf_6 fanout235 (.A(net236),
    .X(net235));
 sky130_fd_sc_hd__buf_12 fanout236 (.A(net239),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_8 fanout237 (.A(net239),
    .X(net237));
 sky130_fd_sc_hd__buf_6 fanout238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__buf_12 fanout239 (.A(_0891_),
    .X(net239));
 sky130_fd_sc_hd__buf_8 fanout24 (.A(net26),
    .X(net24));
 sky130_fd_sc_hd__buf_12 fanout240 (.A(net241),
    .X(net240));
 sky130_fd_sc_hd__buf_12 fanout241 (.A(_0770_),
    .X(net241));
 sky130_fd_sc_hd__buf_12 fanout242 (.A(net244),
    .X(net242));
 sky130_fd_sc_hd__buf_8 fanout243 (.A(net244),
    .X(net243));
 sky130_fd_sc_hd__buf_12 fanout244 (.A(_0759_),
    .X(net244));
 sky130_fd_sc_hd__buf_4 fanout245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_4 fanout246 (.A(net248),
    .X(net246));
 sky130_fd_sc_hd__buf_4 fanout247 (.A(net248),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_8 fanout248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__buf_6 fanout249 (.A(net250),
    .X(net249));
 sky130_fd_sc_hd__buf_4 fanout25 (.A(net26),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_16 fanout250 (.A(net254),
    .X(net250));
 sky130_fd_sc_hd__buf_6 fanout251 (.A(net253),
    .X(net251));
 sky130_fd_sc_hd__buf_4 fanout252 (.A(net253),
    .X(net252));
 sky130_fd_sc_hd__buf_6 fanout253 (.A(net254),
    .X(net253));
 sky130_fd_sc_hd__buf_6 fanout254 (.A(_0869_),
    .X(net254));
 sky130_fd_sc_hd__buf_4 fanout255 (.A(net256),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_4 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__buf_4 fanout257 (.A(net260),
    .X(net257));
 sky130_fd_sc_hd__buf_4 fanout258 (.A(net259),
    .X(net258));
 sky130_fd_sc_hd__buf_2 fanout259 (.A(net260),
    .X(net259));
 sky130_fd_sc_hd__buf_8 fanout26 (.A(_1573_),
    .X(net26));
 sky130_fd_sc_hd__buf_6 fanout260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_16 fanout261 (.A(_0858_),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_8 fanout262 (.A(net263),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_16 fanout263 (.A(_0858_),
    .X(net263));
 sky130_fd_sc_hd__buf_6 fanout264 (.A(_0748_),
    .X(net264));
 sky130_fd_sc_hd__buf_2 fanout265 (.A(_0748_),
    .X(net265));
 sky130_fd_sc_hd__buf_4 fanout266 (.A(net267),
    .X(net266));
 sky130_fd_sc_hd__buf_4 fanout267 (.A(_0737_),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_8 fanout268 (.A(net269),
    .X(net268));
 sky130_fd_sc_hd__buf_6 fanout269 (.A(_1145_),
    .X(net269));
 sky130_fd_sc_hd__buf_6 fanout27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 fanout270 (.A(net271),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_4 fanout271 (.A(_0715_),
    .X(net271));
 sky130_fd_sc_hd__buf_6 fanout272 (.A(_0704_),
    .X(net272));
 sky130_fd_sc_hd__buf_2 fanout273 (.A(_0704_),
    .X(net273));
 sky130_fd_sc_hd__buf_4 fanout274 (.A(net275),
    .X(net274));
 sky130_fd_sc_hd__buf_4 fanout275 (.A(_1125_),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_4 fanout276 (.A(\vgatest.bitmapColAddr[11] ),
    .X(net276));
 sky130_fd_sc_hd__buf_6 fanout277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_16 fanout278 (.A(net2),
    .X(net278));
 sky130_fd_sc_hd__buf_4 fanout28 (.A(_1534_),
    .X(net28));
 sky130_fd_sc_hd__buf_8 fanout29 (.A(_1521_),
    .X(net29));
 sky130_fd_sc_hd__buf_6 fanout30 (.A(_1521_),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_16 fanout31 (.A(_1521_),
    .X(net31));
 sky130_fd_sc_hd__buf_6 fanout32 (.A(net34),
    .X(net32));
 sky130_fd_sc_hd__buf_8 fanout33 (.A(net34),
    .X(net33));
 sky130_fd_sc_hd__buf_12 fanout34 (.A(_1505_),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_16 fanout35 (.A(_1493_),
    .X(net35));
 sky130_fd_sc_hd__buf_12 fanout36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__buf_12 fanout37 (.A(_1483_),
    .X(net37));
 sky130_fd_sc_hd__buf_6 fanout38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__buf_8 fanout39 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__buf_12 fanout40 (.A(_1451_),
    .X(net40));
 sky130_fd_sc_hd__buf_6 fanout41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__buf_6 fanout42 (.A(_1427_),
    .X(net42));
 sky130_fd_sc_hd__buf_12 fanout43 (.A(_1403_),
    .X(net43));
 sky130_fd_sc_hd__buf_8 fanout44 (.A(net47),
    .X(net44));
 sky130_fd_sc_hd__buf_8 fanout45 (.A(net47),
    .X(net45));
 sky130_fd_sc_hd__buf_6 fanout46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__buf_12 fanout47 (.A(_1387_),
    .X(net47));
 sky130_fd_sc_hd__buf_8 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__buf_12 fanout49 (.A(_1372_),
    .X(net49));
 sky130_fd_sc_hd__buf_6 fanout50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__buf_8 fanout51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__buf_12 fanout52 (.A(_1353_),
    .X(net52));
 sky130_fd_sc_hd__buf_8 fanout53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_16 fanout54 (.A(net56),
    .X(net54));
 sky130_fd_sc_hd__buf_12 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__buf_6 fanout56 (.A(_1338_),
    .X(net56));
 sky130_fd_sc_hd__buf_8 fanout57 (.A(net60),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_8 fanout58 (.A(net60),
    .X(net58));
 sky130_fd_sc_hd__buf_12 fanout59 (.A(net60),
    .X(net59));
 sky130_fd_sc_hd__buf_8 fanout60 (.A(_1314_),
    .X(net60));
 sky130_fd_sc_hd__buf_6 fanout61 (.A(net62),
    .X(net61));
 sky130_fd_sc_hd__buf_6 fanout62 (.A(_1263_),
    .X(net62));
 sky130_fd_sc_hd__buf_8 fanout63 (.A(_1263_),
    .X(net63));
 sky130_fd_sc_hd__buf_6 fanout64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__buf_8 fanout65 (.A(net66),
    .X(net65));
 sky130_fd_sc_hd__buf_12 fanout66 (.A(_0627_),
    .X(net66));
 sky130_fd_sc_hd__buf_8 fanout67 (.A(_1957_),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_16 fanout68 (.A(_1868_),
    .X(net68));
 sky130_fd_sc_hd__buf_12 fanout69 (.A(_1785_),
    .X(net69));
 sky130_fd_sc_hd__buf_12 fanout70 (.A(_1569_),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_16 fanout71 (.A(_1513_),
    .X(net71));
 sky130_fd_sc_hd__buf_8 fanout72 (.A(_1512_),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_16 fanout73 (.A(_1507_),
    .X(net73));
 sky130_fd_sc_hd__buf_12 fanout74 (.A(_1441_),
    .X(net74));
 sky130_fd_sc_hd__buf_12 fanout75 (.A(_1438_),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_16 fanout76 (.A(_1413_),
    .X(net76));
 sky130_fd_sc_hd__buf_12 fanout77 (.A(net79),
    .X(net77));
 sky130_fd_sc_hd__buf_8 fanout78 (.A(net79),
    .X(net78));
 sky130_fd_sc_hd__buf_12 fanout79 (.A(_1409_),
    .X(net79));
 sky130_fd_sc_hd__buf_12 fanout80 (.A(_1409_),
    .X(net80));
 sky130_fd_sc_hd__buf_12 fanout81 (.A(_1408_),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_16 fanout82 (.A(_1328_),
    .X(net82));
 sky130_fd_sc_hd__buf_6 fanout83 (.A(net84),
    .X(net83));
 sky130_fd_sc_hd__buf_12 fanout84 (.A(_1317_),
    .X(net84));
 sky130_fd_sc_hd__buf_12 fanout85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__buf_12 fanout86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__buf_12 fanout87 (.A(_1300_),
    .X(net87));
 sky130_fd_sc_hd__buf_8 fanout88 (.A(net90),
    .X(net88));
 sky130_fd_sc_hd__buf_12 fanout89 (.A(net90),
    .X(net89));
 sky130_fd_sc_hd__buf_8 fanout90 (.A(_1299_),
    .X(net90));
 sky130_fd_sc_hd__buf_12 fanout91 (.A(net93),
    .X(net91));
 sky130_fd_sc_hd__buf_12 fanout92 (.A(net93),
    .X(net92));
 sky130_fd_sc_hd__buf_12 fanout93 (.A(_1295_),
    .X(net93));
 sky130_fd_sc_hd__buf_8 fanout94 (.A(_1293_),
    .X(net94));
 sky130_fd_sc_hd__buf_12 fanout95 (.A(_1273_),
    .X(net95));
 sky130_fd_sc_hd__buf_12 fanout96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__buf_12 fanout97 (.A(_1273_),
    .X(net97));
 sky130_fd_sc_hd__buf_12 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__buf_12 fanout99 (.A(_1272_),
    .X(net99));
 sky130_fd_sc_hd__buf_6 input1 (.A(io_in),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(rst),
    .X(net2));
 sky130_fd_sc_hd__buf_4 output10 (.A(net10),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_4 output11 (.A(net11),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_4 output12 (.A(net12),
    .X(io_out[9]));
 sky130_fd_sc_hd__buf_4 output3 (.A(net3),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_4 output4 (.A(net4),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_4 output5 (.A(net5),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_4 output6 (.A(net6),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_4 output7 (.A(net7),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_4 output8 (.A(net8),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_4 output9 (.A(net9),
    .X(io_out[6]));
endmodule

