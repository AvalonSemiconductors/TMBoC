magic
tech sky130B
magscale 1 2
timestamp 1682097309
<< viali >>
rect 9689 37281 9723 37315
rect 12173 37281 12207 37315
rect 26525 37281 26559 37315
rect 28641 37281 28675 37315
rect 32597 37281 32631 37315
rect 33609 37281 33643 37315
rect 1869 37213 1903 37247
rect 5089 37213 5123 37247
rect 7941 37213 7975 37247
rect 11805 37213 11839 37247
rect 15209 37213 15243 37247
rect 18245 37213 18279 37247
rect 22109 37213 22143 37247
rect 25145 37213 25179 37247
rect 26433 37213 26467 37247
rect 26617 37213 26651 37247
rect 28457 37213 28491 37247
rect 32413 37213 32447 37247
rect 33793 37213 33827 37247
rect 36461 37213 36495 37247
rect 37657 37213 37691 37247
rect 2697 37145 2731 37179
rect 5825 37145 5859 37179
rect 8493 37145 8527 37179
rect 9505 37145 9539 37179
rect 15761 37145 15795 37179
rect 18613 37145 18647 37179
rect 22845 37145 22879 37179
rect 25513 37145 25547 37179
rect 36737 37145 36771 37179
rect 38025 37145 38059 37179
rect 9137 37077 9171 37111
rect 9597 37077 9631 37111
rect 33977 37077 34011 37111
rect 6561 36873 6595 36907
rect 9321 36873 9355 36907
rect 4712 36805 4746 36839
rect 8208 36805 8242 36839
rect 26341 36805 26375 36839
rect 34498 36805 34532 36839
rect 36737 36805 36771 36839
rect 4445 36737 4479 36771
rect 6929 36737 6963 36771
rect 12081 36737 12115 36771
rect 12348 36737 12382 36771
rect 14289 36737 14323 36771
rect 16865 36737 16899 36771
rect 17785 36737 17819 36771
rect 22017 36737 22051 36771
rect 22273 36737 22307 36771
rect 23949 36737 23983 36771
rect 26249 36737 26283 36771
rect 27537 36737 27571 36771
rect 27804 36737 27838 36771
rect 29469 36737 29503 36771
rect 29736 36737 29770 36771
rect 32321 36737 32355 36771
rect 32577 36737 32611 36771
rect 36461 36737 36495 36771
rect 37841 36737 37875 36771
rect 7021 36669 7055 36703
rect 7205 36669 7239 36703
rect 7941 36669 7975 36703
rect 14565 36669 14599 36703
rect 18061 36669 18095 36703
rect 20269 36669 20303 36703
rect 21005 36669 21039 36703
rect 24225 36669 24259 36703
rect 34253 36669 34287 36703
rect 38117 36669 38151 36703
rect 5825 36601 5859 36635
rect 16037 36601 16071 36635
rect 13461 36533 13495 36567
rect 16957 36533 16991 36567
rect 19533 36533 19567 36567
rect 23397 36533 23431 36567
rect 25697 36533 25731 36567
rect 28917 36533 28951 36567
rect 30849 36533 30883 36567
rect 33701 36533 33735 36567
rect 35633 36533 35667 36567
rect 12633 36329 12667 36363
rect 15301 36329 15335 36363
rect 19533 36329 19567 36363
rect 27445 36329 27479 36363
rect 28181 36329 28215 36363
rect 30113 36329 30147 36363
rect 31585 36329 31619 36363
rect 32689 36329 32723 36363
rect 33609 36329 33643 36363
rect 9229 36261 9263 36295
rect 25145 36261 25179 36295
rect 5641 36193 5675 36227
rect 5825 36193 5859 36227
rect 9597 36193 9631 36227
rect 13093 36193 13127 36227
rect 13277 36193 13311 36227
rect 15853 36193 15887 36227
rect 23949 36193 23983 36227
rect 25237 36193 25271 36227
rect 26065 36193 26099 36227
rect 31217 36193 31251 36227
rect 34897 36193 34931 36227
rect 6377 36125 6411 36159
rect 10517 36125 10551 36159
rect 13001 36125 13035 36159
rect 15209 36125 15243 36159
rect 16221 36125 16255 36159
rect 18429 36125 18463 36159
rect 19441 36125 19475 36159
rect 20269 36125 20303 36159
rect 24685 36125 24719 36159
rect 24777 36125 24811 36159
rect 26341 36125 26375 36159
rect 28365 36125 28399 36159
rect 28641 36125 28675 36159
rect 29745 36125 29779 36159
rect 30021 36125 30055 36159
rect 31309 36125 31343 36159
rect 32597 36125 32631 36159
rect 32781 36125 32815 36159
rect 33425 36125 33459 36159
rect 36829 36125 36863 36159
rect 5549 36057 5583 36091
rect 6644 36057 6678 36091
rect 9781 36057 9815 36091
rect 10784 36057 10818 36091
rect 18705 36057 18739 36091
rect 20545 36057 20579 36091
rect 21465 36057 21499 36091
rect 23765 36057 23799 36091
rect 28549 36057 28583 36091
rect 33241 36057 33275 36091
rect 35142 36057 35176 36091
rect 37096 36057 37130 36091
rect 5181 35989 5215 36023
rect 7757 35989 7791 36023
rect 9689 35989 9723 36023
rect 11897 35989 11931 36023
rect 17647 35989 17681 36023
rect 22477 35989 22511 36023
rect 25513 35989 25547 36023
rect 30297 35989 30331 36023
rect 36277 35989 36311 36023
rect 38209 35989 38243 36023
rect 7113 35785 7147 35819
rect 7573 35785 7607 35819
rect 11713 35785 11747 35819
rect 12173 35785 12207 35819
rect 22017 35785 22051 35819
rect 22477 35785 22511 35819
rect 26525 35785 26559 35819
rect 33701 35785 33735 35819
rect 36829 35785 36863 35819
rect 37473 35785 37507 35819
rect 7481 35717 7515 35751
rect 26341 35717 26375 35751
rect 9965 35649 9999 35683
rect 12081 35649 12115 35683
rect 13369 35649 13403 35683
rect 16865 35649 16899 35683
rect 17693 35649 17727 35683
rect 18797 35649 18831 35683
rect 19809 35649 19843 35683
rect 19993 35649 20027 35683
rect 20453 35649 20487 35683
rect 22385 35649 22419 35683
rect 23213 35649 23247 35683
rect 23397 35649 23431 35683
rect 24961 35649 24995 35683
rect 26617 35649 26651 35683
rect 27261 35649 27295 35683
rect 28641 35649 28675 35683
rect 28908 35649 28942 35683
rect 32781 35649 32815 35683
rect 32965 35649 32999 35683
rect 33057 35649 33091 35683
rect 33609 35649 33643 35683
rect 33793 35649 33827 35683
rect 36737 35649 36771 35683
rect 37841 35649 37875 35683
rect 7665 35581 7699 35615
rect 10057 35581 10091 35615
rect 10149 35581 10183 35615
rect 12265 35581 12299 35615
rect 13645 35581 13679 35615
rect 17969 35581 18003 35615
rect 19073 35581 19107 35615
rect 20729 35581 20763 35615
rect 22661 35581 22695 35615
rect 23673 35581 23707 35615
rect 24869 35581 24903 35615
rect 25421 35581 25455 35615
rect 27537 35581 27571 35615
rect 37933 35581 37967 35615
rect 38025 35581 38059 35615
rect 26341 35513 26375 35547
rect 32781 35513 32815 35547
rect 9597 35445 9631 35479
rect 15117 35445 15151 35479
rect 16957 35445 16991 35479
rect 19809 35445 19843 35479
rect 25329 35445 25363 35479
rect 25697 35445 25731 35479
rect 30021 35445 30055 35479
rect 10517 35241 10551 35275
rect 14841 35241 14875 35275
rect 17141 35241 17175 35275
rect 20913 35241 20947 35275
rect 23581 35241 23615 35275
rect 29009 35241 29043 35275
rect 31309 35241 31343 35275
rect 32413 35241 32447 35275
rect 33057 35241 33091 35275
rect 33241 35241 33275 35275
rect 11345 35173 11379 35207
rect 18889 35173 18923 35207
rect 5733 35105 5767 35139
rect 12725 35105 12759 35139
rect 15393 35105 15427 35139
rect 20269 35105 20303 35139
rect 22385 35105 22419 35139
rect 23673 35105 23707 35139
rect 29101 35105 29135 35139
rect 36277 35105 36311 35139
rect 9137 35037 9171 35071
rect 12817 35037 12851 35071
rect 13001 35037 13035 35071
rect 14749 35037 14783 35071
rect 18245 35037 18279 35071
rect 19809 35037 19843 35071
rect 20111 35037 20145 35071
rect 22109 35037 22143 35071
rect 23121 35037 23155 35071
rect 23213 35037 23247 35071
rect 27353 35037 27387 35071
rect 27446 35037 27480 35071
rect 28825 35037 28859 35071
rect 28917 35037 28951 35071
rect 30665 35037 30699 35071
rect 30758 35037 30792 35071
rect 31033 35037 31067 35071
rect 31171 35037 31205 35071
rect 31769 35037 31803 35071
rect 31917 35037 31951 35071
rect 32234 35037 32268 35071
rect 5457 34969 5491 35003
rect 9404 34969 9438 35003
rect 11621 34969 11655 35003
rect 11805 34969 11839 35003
rect 11897 34969 11931 35003
rect 13461 34969 13495 35003
rect 15669 34969 15703 35003
rect 18613 34969 18647 35003
rect 18730 34969 18764 35003
rect 19901 34969 19935 35003
rect 19993 34969 20027 35003
rect 20729 34969 20763 35003
rect 25145 34969 25179 35003
rect 30941 34969 30975 35003
rect 32045 34969 32079 35003
rect 32137 34969 32171 35003
rect 32873 34969 32907 35003
rect 36522 34969 36556 35003
rect 5089 34901 5123 34935
rect 5549 34901 5583 34935
rect 18521 34901 18555 34935
rect 19625 34901 19659 34935
rect 20913 34901 20947 34935
rect 21097 34901 21131 34935
rect 23949 34901 23983 34935
rect 26433 34901 26467 34935
rect 27721 34901 27755 34935
rect 33073 34901 33107 34935
rect 37657 34901 37691 34935
rect 5733 34697 5767 34731
rect 9597 34697 9631 34731
rect 10057 34697 10091 34731
rect 20453 34697 20487 34731
rect 36185 34697 36219 34731
rect 9965 34629 9999 34663
rect 34406 34629 34440 34663
rect 4353 34561 4387 34595
rect 4620 34561 4654 34595
rect 7573 34561 7607 34595
rect 7665 34561 7699 34595
rect 7849 34561 7883 34595
rect 17693 34561 17727 34595
rect 18245 34561 18279 34595
rect 18889 34561 18923 34595
rect 19257 34561 19291 34595
rect 20269 34561 20303 34595
rect 21189 34561 21223 34595
rect 21281 34561 21315 34595
rect 21465 34561 21499 34595
rect 22017 34561 22051 34595
rect 23489 34561 23523 34595
rect 25053 34561 25087 34595
rect 27169 34561 27203 34595
rect 27353 34561 27387 34595
rect 28365 34561 28399 34595
rect 29101 34561 29135 34595
rect 33057 34561 33091 34595
rect 34161 34561 34195 34595
rect 36553 34561 36587 34595
rect 37841 34561 37875 34595
rect 8309 34493 8343 34527
rect 10149 34493 10183 34527
rect 20085 34493 20119 34527
rect 22569 34493 22603 34527
rect 23673 34493 23707 34527
rect 25881 34493 25915 34527
rect 28457 34493 28491 34527
rect 33149 34493 33183 34527
rect 33425 34493 33459 34527
rect 36645 34493 36679 34527
rect 36829 34493 36863 34527
rect 38117 34493 38151 34527
rect 22477 34425 22511 34459
rect 18153 34357 18187 34391
rect 22385 34357 22419 34391
rect 22661 34357 22695 34391
rect 27445 34357 27479 34391
rect 29193 34357 29227 34391
rect 35541 34357 35575 34391
rect 10701 34153 10735 34187
rect 25789 34153 25823 34187
rect 26249 34153 26283 34187
rect 30389 34153 30423 34187
rect 31861 34153 31895 34187
rect 11161 34085 11195 34119
rect 26709 34085 26743 34119
rect 5825 34017 5859 34051
rect 5917 34017 5951 34051
rect 8217 34017 8251 34051
rect 9873 34017 9907 34051
rect 10885 34017 10919 34051
rect 21189 34017 21223 34051
rect 25881 34017 25915 34051
rect 28917 34017 28951 34051
rect 29101 34017 29135 34051
rect 5733 33949 5767 33983
rect 7757 33949 7791 33983
rect 8125 33949 8159 33983
rect 10701 33949 10735 33983
rect 10977 33949 11011 33983
rect 11897 33949 11931 33983
rect 12081 33949 12115 33983
rect 15301 33949 15335 33983
rect 15485 33949 15519 33983
rect 16773 33949 16807 33983
rect 16957 33949 16991 33983
rect 19441 33949 19475 33983
rect 19625 33949 19659 33983
rect 20085 33949 20119 33983
rect 20269 33949 20303 33983
rect 21281 33949 21315 33983
rect 22385 33949 22419 33983
rect 22477 33949 22511 33983
rect 22569 33949 22603 33983
rect 22753 33949 22787 33983
rect 23581 33949 23615 33983
rect 23857 33949 23891 33983
rect 24777 33949 24811 33983
rect 24961 33949 24995 33983
rect 25145 33949 25179 33983
rect 26065 33949 26099 33983
rect 26985 33949 27019 33983
rect 27537 33949 27571 33983
rect 29193 33949 29227 33983
rect 29745 33949 29779 33983
rect 29893 33949 29927 33983
rect 30210 33949 30244 33983
rect 31217 33949 31251 33983
rect 31310 33949 31344 33983
rect 31682 33949 31716 33983
rect 37841 33949 37875 33983
rect 9137 33881 9171 33915
rect 17417 33881 17451 33915
rect 18153 33881 18187 33915
rect 21557 33881 21591 33915
rect 21649 33881 21683 33915
rect 22109 33881 22143 33915
rect 25789 33881 25823 33915
rect 26709 33881 26743 33915
rect 26893 33881 26927 33915
rect 27905 33881 27939 33915
rect 30021 33881 30055 33915
rect 30113 33881 30147 33915
rect 31493 33881 31527 33915
rect 31585 33881 31619 33915
rect 38117 33881 38151 33915
rect 5365 33813 5399 33847
rect 11989 33813 12023 33847
rect 15393 33813 15427 33847
rect 16957 33813 16991 33847
rect 19533 33813 19567 33847
rect 20177 33813 20211 33847
rect 21005 33813 21039 33847
rect 28733 33813 28767 33847
rect 13553 33609 13587 33643
rect 14657 33609 14691 33643
rect 16037 33609 16071 33643
rect 19073 33609 19107 33643
rect 20453 33609 20487 33643
rect 21373 33609 21407 33643
rect 25513 33609 25547 33643
rect 31677 33609 31711 33643
rect 36093 33609 36127 33643
rect 28917 33541 28951 33575
rect 31309 33541 31343 33575
rect 31401 33541 31435 33575
rect 33149 33541 33183 33575
rect 33241 33541 33275 33575
rect 34709 33541 34743 33575
rect 5365 33473 5399 33507
rect 5457 33473 5491 33507
rect 5917 33473 5951 33507
rect 7021 33473 7055 33507
rect 8125 33473 8159 33507
rect 8309 33473 8343 33507
rect 10241 33473 10275 33507
rect 10517 33473 10551 33507
rect 12081 33473 12115 33507
rect 12265 33473 12299 33507
rect 13185 33473 13219 33507
rect 13277 33473 13311 33507
rect 13369 33473 13403 33507
rect 14013 33473 14047 33507
rect 14473 33473 14507 33507
rect 15393 33473 15427 33507
rect 15853 33473 15887 33507
rect 17417 33473 17451 33507
rect 19257 33473 19291 33507
rect 19349 33473 19383 33507
rect 19533 33473 19567 33507
rect 19625 33473 19659 33507
rect 20269 33473 20303 33507
rect 20545 33473 20579 33507
rect 21281 33473 21315 33507
rect 22477 33473 22511 33507
rect 22753 33473 22787 33507
rect 24225 33473 24259 33507
rect 24869 33473 24903 33507
rect 26249 33473 26283 33507
rect 26433 33473 26467 33507
rect 27537 33473 27571 33507
rect 28733 33473 28767 33507
rect 29745 33473 29779 33507
rect 31033 33473 31067 33507
rect 31126 33473 31160 33507
rect 31498 33473 31532 33507
rect 32873 33473 32907 33507
rect 32966 33473 33000 33507
rect 33379 33473 33413 33507
rect 34437 33473 34471 33507
rect 34575 33473 34609 33507
rect 34805 33473 34839 33507
rect 35449 33473 35483 33507
rect 35542 33473 35576 33507
rect 35725 33473 35759 33507
rect 35817 33473 35851 33507
rect 35914 33473 35948 33507
rect 37841 33473 37875 33507
rect 7297 33405 7331 33439
rect 14381 33405 14415 33439
rect 15669 33405 15703 33439
rect 17325 33405 17359 33439
rect 17877 33405 17911 33439
rect 22569 33405 22603 33439
rect 22937 33405 22971 33439
rect 23673 33405 23707 33439
rect 24041 33405 24075 33439
rect 24133 33405 24167 33439
rect 25237 33405 25271 33439
rect 27813 33405 27847 33439
rect 29009 33405 29043 33439
rect 30021 33405 30055 33439
rect 37933 33405 37967 33439
rect 38025 33405 38059 33439
rect 12081 33337 12115 33371
rect 26525 33337 26559 33371
rect 34989 33337 35023 33371
rect 8401 33269 8435 33303
rect 10057 33269 10091 33303
rect 14105 33269 14139 33303
rect 15485 33269 15519 33303
rect 17785 33269 17819 33303
rect 18153 33269 18187 33303
rect 20085 33269 20119 33303
rect 25007 33269 25041 33303
rect 25145 33269 25179 33303
rect 33517 33269 33551 33303
rect 37473 33269 37507 33303
rect 6837 33065 6871 33099
rect 10885 33065 10919 33099
rect 12081 33065 12115 33099
rect 15853 33065 15887 33099
rect 16037 33065 16071 33099
rect 17601 33065 17635 33099
rect 17785 33065 17819 33099
rect 18337 33065 18371 33099
rect 25237 33065 25271 33099
rect 30389 33065 30423 33099
rect 31493 33065 31527 33099
rect 32505 33065 32539 33099
rect 36369 33065 36403 33099
rect 7757 32997 7791 33031
rect 8309 32997 8343 33031
rect 11345 32997 11379 33031
rect 22753 32997 22787 33031
rect 25421 32997 25455 33031
rect 8493 32929 8527 32963
rect 10057 32929 10091 32963
rect 10977 32929 11011 32963
rect 12449 32929 12483 32963
rect 15025 32929 15059 32963
rect 15761 32929 15795 32963
rect 17509 32929 17543 32963
rect 18521 32929 18555 32963
rect 21005 32929 21039 32963
rect 24777 32929 24811 32963
rect 27445 32929 27479 32963
rect 28733 32929 28767 32963
rect 36829 32929 36863 32963
rect 4445 32861 4479 32895
rect 4537 32861 4571 32895
rect 5181 32861 5215 32895
rect 5273 32861 5307 32895
rect 6745 32861 6779 32895
rect 6929 32861 6963 32895
rect 7389 32861 7423 32895
rect 7573 32861 7607 32895
rect 8217 32861 8251 32895
rect 9689 32861 9723 32895
rect 9873 32861 9907 32895
rect 9965 32861 9999 32895
rect 10241 32861 10275 32895
rect 11161 32861 11195 32895
rect 12265 32861 12299 32895
rect 12357 32861 12391 32895
rect 12541 32861 12575 32895
rect 13553 32861 13587 32895
rect 13737 32861 13771 32895
rect 15669 32861 15703 32895
rect 17601 32861 17635 32895
rect 18245 32861 18279 32895
rect 19717 32861 19751 32895
rect 19901 32861 19935 32895
rect 20545 32861 20579 32895
rect 20637 32861 20671 32895
rect 21925 32861 21959 32895
rect 22017 32861 22051 32895
rect 22661 32861 22695 32895
rect 22937 32861 22971 32895
rect 24869 32861 24903 32895
rect 25237 32861 25271 32895
rect 26157 32861 26191 32895
rect 26801 32861 26835 32895
rect 27905 32861 27939 32895
rect 28273 32861 28307 32895
rect 28825 32861 28859 32895
rect 29745 32861 29779 32895
rect 29893 32861 29927 32895
rect 30113 32861 30147 32895
rect 30210 32861 30244 32895
rect 30849 32861 30883 32895
rect 30942 32861 30976 32895
rect 31314 32861 31348 32895
rect 31953 32861 31987 32895
rect 32229 32861 32263 32895
rect 32321 32861 32355 32895
rect 35725 32861 35759 32895
rect 35818 32861 35852 32895
rect 36001 32861 36035 32895
rect 36190 32861 36224 32895
rect 37096 32861 37130 32895
rect 4721 32793 4755 32827
rect 5733 32793 5767 32827
rect 10885 32793 10919 32827
rect 14289 32793 14323 32827
rect 17325 32793 17359 32827
rect 20913 32793 20947 32827
rect 22201 32793 22235 32827
rect 30021 32793 30055 32827
rect 31125 32793 31159 32827
rect 31217 32793 31251 32827
rect 32137 32793 32171 32827
rect 36093 32793 36127 32827
rect 8493 32725 8527 32759
rect 10425 32725 10459 32759
rect 13737 32725 13771 32759
rect 18521 32725 18555 32759
rect 19809 32725 19843 32759
rect 20361 32725 20395 32759
rect 21925 32725 21959 32759
rect 23121 32725 23155 32759
rect 38209 32725 38243 32759
rect 9137 32521 9171 32555
rect 9597 32521 9631 32555
rect 12173 32521 12207 32555
rect 13185 32521 13219 32555
rect 14657 32521 14691 32555
rect 20729 32521 20763 32555
rect 25973 32521 26007 32555
rect 30849 32521 30883 32555
rect 35449 32521 35483 32555
rect 6561 32453 6595 32487
rect 8217 32453 8251 32487
rect 8401 32453 8435 32487
rect 11805 32453 11839 32487
rect 11989 32453 12023 32487
rect 14197 32453 14231 32487
rect 16865 32453 16899 32487
rect 30481 32453 30515 32487
rect 30570 32453 30604 32487
rect 35081 32453 35115 32487
rect 35173 32453 35207 32487
rect 4629 32385 4663 32419
rect 5549 32385 5583 32419
rect 6009 32385 6043 32419
rect 6745 32385 6779 32419
rect 9413 32385 9447 32419
rect 9505 32385 9539 32419
rect 9873 32385 9907 32419
rect 10333 32385 10367 32419
rect 12081 32385 12115 32419
rect 12817 32385 12851 32419
rect 14473 32385 14507 32419
rect 15301 32385 15335 32419
rect 16037 32385 16071 32419
rect 17325 32385 17359 32419
rect 17969 32385 18003 32419
rect 18153 32385 18187 32419
rect 20545 32385 20579 32419
rect 21281 32385 21315 32419
rect 21465 32385 21499 32419
rect 22017 32385 22051 32419
rect 22293 32385 22327 32419
rect 23121 32385 23155 32419
rect 23305 32385 23339 32419
rect 24133 32385 24167 32419
rect 24225 32385 24259 32419
rect 24409 32385 24443 32419
rect 25881 32385 25915 32419
rect 26341 32385 26375 32419
rect 27169 32385 27203 32419
rect 27353 32385 27387 32419
rect 28457 32385 28491 32419
rect 28825 32385 28859 32419
rect 28917 32385 28951 32419
rect 30205 32385 30239 32419
rect 30298 32385 30332 32419
rect 30670 32385 30704 32419
rect 33037 32385 33071 32419
rect 34897 32385 34931 32419
rect 35265 32385 35299 32419
rect 37841 32385 37875 32419
rect 4445 32317 4479 32351
rect 5641 32317 5675 32351
rect 10517 32317 10551 32351
rect 12357 32317 12391 32351
rect 12909 32317 12943 32351
rect 14381 32317 14415 32351
rect 15117 32317 15151 32351
rect 15393 32317 15427 32351
rect 15485 32317 15519 32351
rect 17233 32317 17267 32351
rect 20361 32317 20395 32351
rect 22385 32317 22419 32351
rect 24869 32317 24903 32351
rect 28365 32317 28399 32351
rect 32781 32317 32815 32351
rect 38117 32317 38151 32351
rect 4813 32249 4847 32283
rect 8585 32249 8619 32283
rect 6837 32181 6871 32215
rect 9781 32181 9815 32215
rect 12817 32181 12851 32215
rect 14197 32181 14231 32215
rect 16221 32181 16255 32215
rect 16957 32181 16991 32215
rect 17509 32181 17543 32215
rect 18061 32181 18095 32215
rect 21281 32181 21315 32215
rect 23397 32181 23431 32215
rect 27169 32181 27203 32215
rect 27905 32181 27939 32215
rect 34161 32181 34195 32215
rect 6469 31977 6503 32011
rect 9229 31977 9263 32011
rect 10149 31977 10183 32011
rect 11529 31977 11563 32011
rect 12541 31977 12575 32011
rect 14933 31977 14967 32011
rect 15117 31977 15151 32011
rect 15577 31977 15611 32011
rect 19625 31977 19659 32011
rect 19809 31977 19843 32011
rect 24777 31977 24811 32011
rect 25789 31977 25823 32011
rect 29745 31977 29779 32011
rect 32781 31977 32815 32011
rect 35909 31977 35943 32011
rect 4261 31909 4295 31943
rect 6837 31909 6871 31943
rect 18889 31909 18923 31943
rect 29009 31909 29043 31943
rect 32045 31909 32079 31943
rect 9597 31841 9631 31875
rect 21649 31841 21683 31875
rect 26709 31841 26743 31875
rect 27629 31841 27663 31875
rect 36369 31841 36403 31875
rect 4077 31773 4111 31807
rect 4261 31773 4295 31807
rect 4813 31773 4847 31807
rect 4925 31773 4959 31807
rect 5365 31773 5399 31807
rect 6653 31773 6687 31807
rect 6745 31773 6779 31807
rect 6929 31773 6963 31807
rect 7941 31773 7975 31807
rect 8033 31773 8067 31807
rect 8217 31773 8251 31807
rect 8309 31773 8343 31807
rect 9413 31773 9447 31807
rect 9689 31773 9723 31807
rect 10333 31773 10367 31807
rect 10609 31773 10643 31807
rect 11713 31773 11747 31807
rect 11805 31773 11839 31807
rect 11989 31773 12023 31807
rect 12081 31773 12115 31807
rect 12541 31773 12575 31807
rect 12633 31773 12667 31807
rect 14657 31773 14691 31807
rect 14841 31773 14875 31807
rect 14933 31773 14967 31807
rect 15577 31773 15611 31807
rect 15669 31773 15703 31807
rect 16957 31773 16991 31807
rect 17325 31773 17359 31807
rect 17417 31773 17451 31807
rect 18521 31773 18555 31807
rect 18705 31773 18739 31807
rect 19441 31773 19475 31807
rect 19625 31773 19659 31807
rect 21281 31773 21315 31807
rect 21557 31773 21591 31807
rect 22937 31773 22971 31807
rect 24685 31773 24719 31807
rect 24961 31773 24995 31807
rect 25605 31773 25639 31807
rect 25789 31773 25823 31807
rect 26893 31773 26927 31807
rect 28181 31773 28215 31807
rect 28641 31773 28675 31807
rect 29745 31773 29779 31807
rect 29929 31773 29963 31807
rect 32229 31773 32263 31807
rect 32321 31773 32355 31807
rect 32781 31773 32815 31807
rect 32965 31773 32999 31807
rect 35265 31773 35299 31807
rect 35358 31773 35392 31807
rect 35541 31773 35575 31807
rect 35633 31773 35667 31807
rect 35771 31773 35805 31807
rect 36636 31773 36670 31807
rect 23305 31705 23339 31739
rect 32045 31705 32079 31739
rect 7757 31637 7791 31671
rect 10517 31637 10551 31671
rect 12909 31637 12943 31671
rect 15945 31637 15979 31671
rect 21281 31637 21315 31671
rect 25973 31637 26007 31671
rect 27077 31637 27111 31671
rect 37749 31637 37783 31671
rect 7205 31433 7239 31467
rect 12173 31433 12207 31467
rect 12817 31433 12851 31467
rect 14749 31433 14783 31467
rect 17509 31433 17543 31467
rect 18889 31433 18923 31467
rect 22293 31433 22327 31467
rect 28641 31433 28675 31467
rect 31309 31433 31343 31467
rect 32505 31433 32539 31467
rect 32689 31433 32723 31467
rect 35081 31433 35115 31467
rect 37473 31433 37507 31467
rect 37933 31433 37967 31467
rect 8217 31365 8251 31399
rect 14013 31365 14047 31399
rect 16865 31365 16899 31399
rect 31033 31365 31067 31399
rect 32321 31365 32355 31399
rect 34713 31365 34747 31399
rect 34805 31365 34839 31399
rect 5365 31297 5399 31331
rect 5549 31297 5583 31331
rect 7389 31297 7423 31331
rect 7665 31297 7699 31331
rect 10149 31297 10183 31331
rect 10425 31297 10459 31331
rect 11805 31297 11839 31331
rect 11989 31297 12023 31331
rect 12633 31297 12667 31331
rect 12909 31297 12943 31331
rect 14289 31297 14323 31331
rect 14565 31297 14599 31331
rect 15301 31297 15335 31331
rect 17325 31297 17359 31331
rect 18245 31297 18279 31331
rect 18521 31297 18555 31331
rect 18705 31297 18739 31331
rect 19625 31297 19659 31331
rect 19717 31297 19751 31331
rect 20453 31297 20487 31331
rect 21281 31297 21315 31331
rect 21465 31297 21499 31331
rect 22293 31297 22327 31331
rect 22569 31297 22603 31331
rect 23673 31297 23707 31331
rect 23949 31297 23983 31331
rect 25697 31297 25731 31331
rect 25789 31297 25823 31331
rect 25881 31297 25915 31331
rect 26041 31297 26075 31331
rect 27445 31297 27479 31331
rect 28549 31297 28583 31331
rect 28733 31297 28767 31331
rect 29377 31297 29411 31331
rect 29561 31297 29595 31331
rect 30665 31297 30699 31331
rect 30758 31297 30792 31331
rect 30941 31297 30975 31331
rect 31171 31297 31205 31331
rect 34529 31297 34563 31331
rect 34897 31297 34931 31331
rect 37841 31297 37875 31331
rect 7481 31229 7515 31263
rect 9045 31229 9079 31263
rect 10241 31229 10275 31263
rect 14473 31229 14507 31263
rect 15485 31229 15519 31263
rect 17233 31229 17267 31263
rect 19441 31229 19475 31263
rect 19809 31229 19843 31263
rect 19901 31229 19935 31263
rect 20729 31229 20763 31263
rect 24409 31229 24443 31263
rect 27721 31229 27755 31263
rect 38025 31229 38059 31263
rect 7573 31161 7607 31195
rect 12633 31161 12667 31195
rect 23765 31161 23799 31195
rect 29653 31161 29687 31195
rect 5641 31093 5675 31127
rect 10425 31093 10459 31127
rect 10609 31093 10643 31127
rect 14289 31093 14323 31127
rect 17325 31093 17359 31127
rect 18337 31093 18371 31127
rect 21281 31093 21315 31127
rect 25421 31093 25455 31127
rect 32505 31093 32539 31127
rect 6561 30889 6595 30923
rect 7021 30889 7055 30923
rect 7941 30889 7975 30923
rect 11437 30889 11471 30923
rect 12725 30889 12759 30923
rect 13553 30889 13587 30923
rect 17877 30889 17911 30923
rect 19717 30889 19751 30923
rect 20453 30889 20487 30923
rect 28273 30889 28307 30923
rect 26249 30821 26283 30855
rect 28917 30821 28951 30855
rect 31401 30821 31435 30855
rect 6653 30753 6687 30787
rect 8401 30753 8435 30787
rect 10333 30753 10367 30787
rect 13645 30753 13679 30787
rect 17785 30753 17819 30787
rect 19533 30753 19567 30787
rect 20637 30753 20671 30787
rect 28181 30753 28215 30787
rect 32413 30753 32447 30787
rect 32689 30753 32723 30787
rect 5089 30685 5123 30719
rect 5825 30685 5859 30719
rect 6009 30685 6043 30719
rect 6837 30685 6871 30719
rect 8125 30685 8159 30719
rect 8309 30685 8343 30719
rect 9781 30685 9815 30719
rect 9965 30685 9999 30719
rect 11713 30685 11747 30719
rect 12081 30685 12115 30719
rect 12173 30685 12207 30719
rect 12725 30685 12759 30719
rect 12909 30685 12943 30719
rect 13369 30685 13403 30719
rect 13461 30685 13495 30719
rect 15117 30685 15151 30719
rect 15301 30685 15335 30719
rect 15393 30685 15427 30719
rect 15485 30685 15519 30719
rect 15669 30685 15703 30719
rect 16405 30685 16439 30719
rect 16589 30685 16623 30719
rect 17877 30685 17911 30719
rect 19717 30685 19751 30719
rect 20361 30685 20395 30719
rect 22293 30685 22327 30719
rect 22661 30685 22695 30719
rect 23305 30685 23339 30719
rect 23397 30685 23431 30719
rect 23581 30685 23615 30719
rect 24961 30685 24995 30719
rect 25145 30685 25179 30719
rect 25329 30685 25363 30719
rect 25421 30685 25455 30719
rect 25881 30685 25915 30719
rect 26709 30685 26743 30719
rect 26893 30685 26927 30719
rect 27353 30685 27387 30719
rect 27537 30685 27571 30719
rect 28089 30685 28123 30719
rect 28917 30685 28951 30719
rect 29101 30685 29135 30719
rect 29745 30685 29779 30719
rect 30757 30685 30791 30719
rect 30850 30685 30884 30719
rect 31263 30685 31297 30719
rect 32321 30685 32355 30719
rect 35081 30685 35115 30719
rect 35357 30685 35391 30719
rect 35449 30685 35483 30719
rect 36737 30685 36771 30719
rect 4905 30617 4939 30651
rect 5273 30617 5307 30651
rect 6101 30617 6135 30651
rect 6561 30617 6595 30651
rect 11897 30617 11931 30651
rect 16773 30617 16807 30651
rect 17601 30617 17635 30651
rect 19441 30617 19475 30651
rect 22845 30617 22879 30651
rect 26065 30617 26099 30651
rect 29929 30617 29963 30651
rect 30113 30617 30147 30651
rect 31033 30617 31067 30651
rect 31125 30617 31159 30651
rect 35265 30617 35299 30651
rect 37013 30617 37047 30651
rect 37749 30617 37783 30651
rect 11805 30549 11839 30583
rect 15853 30549 15887 30583
rect 18061 30549 18095 30583
rect 19901 30549 19935 30583
rect 20637 30549 20671 30583
rect 23765 30549 23799 30583
rect 26801 30549 26835 30583
rect 27445 30549 27479 30583
rect 28457 30549 28491 30583
rect 35633 30549 35667 30583
rect 38025 30549 38059 30583
rect 15117 30345 15151 30379
rect 30389 30345 30423 30379
rect 35173 30345 35207 30379
rect 36461 30345 36495 30379
rect 37841 30345 37875 30379
rect 10517 30277 10551 30311
rect 12449 30277 12483 30311
rect 13829 30277 13863 30311
rect 20269 30277 20303 30311
rect 24317 30277 24351 30311
rect 31401 30277 31435 30311
rect 34060 30277 34094 30311
rect 36185 30277 36219 30311
rect 37933 30277 37967 30311
rect 2881 30209 2915 30243
rect 3148 30209 3182 30243
rect 5181 30209 5215 30243
rect 6745 30209 6779 30243
rect 7021 30209 7055 30243
rect 8677 30209 8711 30243
rect 9045 30209 9079 30243
rect 9965 30209 9999 30243
rect 10149 30209 10183 30243
rect 12081 30209 12115 30243
rect 12265 30209 12299 30243
rect 12909 30209 12943 30243
rect 14013 30209 14047 30243
rect 14105 30209 14139 30243
rect 14749 30209 14783 30243
rect 15209 30209 15243 30243
rect 15669 30209 15703 30243
rect 17417 30209 17451 30243
rect 18245 30209 18279 30243
rect 18429 30209 18463 30243
rect 20453 30209 20487 30243
rect 22661 30209 22695 30243
rect 24501 30209 24535 30243
rect 26065 30209 26099 30243
rect 26433 30209 26467 30243
rect 26525 30209 26559 30243
rect 27169 30209 27203 30243
rect 27629 30209 27663 30243
rect 28365 30209 28399 30243
rect 28512 30209 28546 30243
rect 29745 30209 29779 30243
rect 29838 30209 29872 30243
rect 30021 30209 30055 30243
rect 30113 30209 30147 30243
rect 30251 30209 30285 30243
rect 30757 30209 30791 30243
rect 31125 30209 31159 30243
rect 31273 30209 31307 30243
rect 31493 30209 31527 30243
rect 31590 30209 31624 30243
rect 35817 30209 35851 30243
rect 35910 30209 35944 30243
rect 36093 30209 36127 30243
rect 36282 30209 36316 30243
rect 5365 30141 5399 30175
rect 6561 30141 6595 30175
rect 6837 30141 6871 30175
rect 13185 30141 13219 30175
rect 15761 30141 15795 30175
rect 17509 30141 17543 30175
rect 23029 30141 23063 30175
rect 23213 30141 23247 30175
rect 24685 30141 24719 30175
rect 26157 30141 26191 30175
rect 27721 30141 27755 30175
rect 28733 30141 28767 30175
rect 33793 30141 33827 30175
rect 38025 30141 38059 30175
rect 6929 30073 6963 30107
rect 14289 30073 14323 30107
rect 17785 30073 17819 30107
rect 22799 30073 22833 30107
rect 22937 30073 22971 30107
rect 4261 30005 4295 30039
rect 8217 30005 8251 30039
rect 13829 30005 13863 30039
rect 14887 30005 14921 30039
rect 15025 30005 15059 30039
rect 15669 30005 15703 30039
rect 16037 30005 16071 30039
rect 17417 30005 17451 30039
rect 18245 30005 18279 30039
rect 20637 30005 20671 30039
rect 25513 30005 25547 30039
rect 28641 30005 28675 30039
rect 29009 30005 29043 30039
rect 31769 30005 31803 30039
rect 37473 30005 37507 30039
rect 3985 29801 4019 29835
rect 10425 29801 10459 29835
rect 11805 29801 11839 29835
rect 11989 29801 12023 29835
rect 12449 29801 12483 29835
rect 15945 29801 15979 29835
rect 17325 29801 17359 29835
rect 17785 29801 17819 29835
rect 20269 29801 20303 29835
rect 22293 29801 22327 29835
rect 23397 29801 23431 29835
rect 25973 29801 26007 29835
rect 30481 29801 30515 29835
rect 38209 29801 38243 29835
rect 11437 29733 11471 29767
rect 12817 29733 12851 29767
rect 21281 29733 21315 29767
rect 22845 29733 22879 29767
rect 32413 29733 32447 29767
rect 4537 29665 4571 29699
rect 5641 29665 5675 29699
rect 15025 29665 15059 29699
rect 17417 29665 17451 29699
rect 21465 29665 21499 29699
rect 22477 29665 22511 29699
rect 27353 29665 27387 29699
rect 31861 29665 31895 29699
rect 36829 29665 36863 29699
rect 3249 29597 3283 29631
rect 3433 29597 3467 29631
rect 4353 29597 4387 29631
rect 5365 29597 5399 29631
rect 5549 29597 5583 29631
rect 6101 29597 6135 29631
rect 6285 29597 6319 29631
rect 7021 29597 7055 29631
rect 7297 29597 7331 29631
rect 7573 29597 7607 29631
rect 7757 29597 7791 29631
rect 12449 29597 12483 29631
rect 12541 29597 12575 29631
rect 13277 29597 13311 29631
rect 13461 29597 13495 29631
rect 15853 29597 15887 29631
rect 16589 29597 16623 29631
rect 16773 29597 16807 29631
rect 17601 29597 17635 29631
rect 20453 29597 20487 29631
rect 20637 29597 20671 29631
rect 20729 29597 20763 29631
rect 21189 29597 21223 29631
rect 22206 29597 22240 29631
rect 22661 29597 22695 29631
rect 23305 29597 23339 29631
rect 23489 29597 23523 29631
rect 24593 29597 24627 29631
rect 24777 29597 24811 29631
rect 26893 29597 26927 29631
rect 27077 29597 27111 29631
rect 28273 29597 28307 29631
rect 29837 29597 29871 29631
rect 29985 29597 30019 29631
rect 30113 29597 30147 29631
rect 30343 29597 30377 29631
rect 32413 29597 32447 29631
rect 32689 29597 32723 29631
rect 33149 29597 33183 29631
rect 33333 29597 33367 29631
rect 35265 29597 35299 29631
rect 35541 29597 35575 29631
rect 35633 29597 35667 29631
rect 37096 29597 37130 29631
rect 9137 29529 9171 29563
rect 11805 29529 11839 29563
rect 14289 29529 14323 29563
rect 17325 29529 17359 29563
rect 25789 29529 25823 29563
rect 28549 29529 28583 29563
rect 30205 29529 30239 29563
rect 31033 29529 31067 29563
rect 35449 29529 35483 29563
rect 3341 29461 3375 29495
rect 4445 29461 4479 29495
rect 5181 29461 5215 29495
rect 6193 29461 6227 29495
rect 7297 29461 7331 29495
rect 13369 29461 13403 29495
rect 16681 29461 16715 29495
rect 21465 29461 21499 29495
rect 24685 29461 24719 29495
rect 25989 29461 26023 29495
rect 26157 29461 26191 29495
rect 32597 29461 32631 29495
rect 33241 29461 33275 29495
rect 35817 29461 35851 29495
rect 10517 29257 10551 29291
rect 11805 29257 11839 29291
rect 15853 29257 15887 29291
rect 23397 29257 23431 29291
rect 24961 29257 24995 29291
rect 26341 29257 26375 29291
rect 32505 29257 32539 29291
rect 32689 29257 32723 29291
rect 36369 29257 36403 29291
rect 4261 29189 4295 29223
rect 4353 29189 4387 29223
rect 7665 29189 7699 29223
rect 8861 29189 8895 29223
rect 19533 29189 19567 29223
rect 27721 29189 27755 29223
rect 29377 29189 29411 29223
rect 32321 29189 32355 29223
rect 33578 29189 33612 29223
rect 36093 29189 36127 29223
rect 4077 29121 4111 29155
rect 4445 29121 4479 29155
rect 5089 29121 5123 29155
rect 5273 29121 5307 29155
rect 7297 29121 7331 29155
rect 9137 29121 9171 29155
rect 10057 29121 10091 29155
rect 10333 29121 10367 29155
rect 11713 29121 11747 29155
rect 11897 29121 11931 29155
rect 12817 29121 12851 29155
rect 13645 29121 13679 29155
rect 16037 29121 16071 29155
rect 16865 29121 16899 29155
rect 17049 29121 17083 29155
rect 17969 29121 18003 29155
rect 19349 29121 19383 29155
rect 19717 29121 19751 29155
rect 20269 29121 20303 29155
rect 20361 29121 20395 29155
rect 20729 29121 20763 29155
rect 22569 29121 22603 29155
rect 22753 29121 22787 29155
rect 23581 29121 23615 29155
rect 23765 29121 23799 29155
rect 25145 29121 25179 29155
rect 25329 29121 25363 29155
rect 25421 29121 25455 29155
rect 25973 29121 26007 29155
rect 27353 29121 27387 29155
rect 27537 29121 27571 29155
rect 28181 29121 28215 29155
rect 28365 29121 28399 29155
rect 28457 29121 28491 29155
rect 28549 29121 28583 29155
rect 29653 29121 29687 29155
rect 30389 29121 30423 29155
rect 30941 29121 30975 29155
rect 35725 29121 35759 29155
rect 35818 29121 35852 29155
rect 36001 29121 36035 29155
rect 36231 29121 36265 29155
rect 37473 29121 37507 29155
rect 9045 29053 9079 29087
rect 10149 29053 10183 29087
rect 12909 29053 12943 29087
rect 14381 29053 14415 29087
rect 16221 29053 16255 29087
rect 16313 29053 16347 29087
rect 17417 29053 17451 29087
rect 18521 29053 18555 29087
rect 18797 29053 18831 29087
rect 23673 29053 23707 29087
rect 23857 29053 23891 29087
rect 25237 29053 25271 29087
rect 26065 29053 26099 29087
rect 29561 29053 29595 29087
rect 30757 29053 30791 29087
rect 33333 29053 33367 29087
rect 37749 29053 37783 29087
rect 4629 28985 4663 29019
rect 9321 28985 9355 29019
rect 13185 28985 13219 29019
rect 18429 28985 18463 29019
rect 20913 28985 20947 29019
rect 22937 28985 22971 29019
rect 27353 28985 27387 29019
rect 28733 28985 28767 29019
rect 29837 28985 29871 29019
rect 34713 28985 34747 29019
rect 5457 28917 5491 28951
rect 8861 28917 8895 28951
rect 10057 28917 10091 28951
rect 12817 28917 12851 28951
rect 18337 28917 18371 28951
rect 20729 28917 20763 28951
rect 26157 28917 26191 28951
rect 29377 28917 29411 28951
rect 32505 28917 32539 28951
rect 4629 28713 4663 28747
rect 11069 28713 11103 28747
rect 11989 28713 12023 28747
rect 14841 28713 14875 28747
rect 16129 28713 16163 28747
rect 17877 28713 17911 28747
rect 23305 28713 23339 28747
rect 24961 28713 24995 28747
rect 11253 28645 11287 28679
rect 16405 28645 16439 28679
rect 23397 28645 23431 28679
rect 25053 28645 25087 28679
rect 31953 28645 31987 28679
rect 16497 28577 16531 28611
rect 21281 28577 21315 28611
rect 25145 28577 25179 28611
rect 30481 28577 30515 28611
rect 32689 28577 32723 28611
rect 33149 28577 33183 28611
rect 35725 28577 35759 28611
rect 36829 28577 36863 28611
rect 4537 28509 4571 28543
rect 5181 28509 5215 28543
rect 5365 28509 5399 28543
rect 5549 28509 5583 28543
rect 8309 28509 8343 28543
rect 8401 28509 8435 28543
rect 9137 28509 9171 28543
rect 9597 28509 9631 28543
rect 12725 28509 12759 28543
rect 12909 28509 12943 28543
rect 14289 28509 14323 28543
rect 14473 28509 14507 28543
rect 14657 28509 14691 28543
rect 16313 28509 16347 28543
rect 16589 28509 16623 28543
rect 16773 28509 16807 28543
rect 17785 28509 17819 28543
rect 17969 28509 18003 28543
rect 19717 28509 19751 28543
rect 19809 28509 19843 28543
rect 19901 28509 19935 28543
rect 20085 28509 20119 28543
rect 21005 28509 21039 28543
rect 23121 28509 23155 28543
rect 23213 28509 23247 28543
rect 23581 28509 23615 28543
rect 24593 28509 24627 28543
rect 27261 28509 27295 28543
rect 27997 28509 28031 28543
rect 28365 28509 28399 28543
rect 30205 28509 30239 28543
rect 31309 28509 31343 28543
rect 31402 28509 31436 28543
rect 31585 28509 31619 28543
rect 31774 28509 31808 28543
rect 32781 28509 32815 28543
rect 5457 28441 5491 28475
rect 6653 28441 6687 28475
rect 6837 28441 6871 28475
rect 7021 28441 7055 28475
rect 10885 28441 10919 28475
rect 11805 28441 11839 28475
rect 11989 28441 12023 28475
rect 14565 28441 14599 28475
rect 21490 28441 21524 28475
rect 28181 28441 28215 28475
rect 28273 28441 28307 28475
rect 31677 28441 31711 28475
rect 34897 28441 34931 28475
rect 37096 28441 37130 28475
rect 5733 28373 5767 28407
rect 8309 28373 8343 28407
rect 9229 28373 9263 28407
rect 11069 28373 11103 28407
rect 12173 28373 12207 28407
rect 12817 28373 12851 28407
rect 19441 28373 19475 28407
rect 21373 28373 21407 28407
rect 21649 28373 21683 28407
rect 22845 28373 22879 28407
rect 25421 28373 25455 28407
rect 27445 28373 27479 28407
rect 28549 28373 28583 28407
rect 38209 28373 38243 28407
rect 11069 28169 11103 28203
rect 16957 28169 16991 28203
rect 24133 28169 24167 28203
rect 25605 28169 25639 28203
rect 30757 28169 30791 28203
rect 36277 28169 36311 28203
rect 37473 28169 37507 28203
rect 37933 28169 37967 28203
rect 7297 28101 7331 28135
rect 14197 28101 14231 28135
rect 22569 28101 22603 28135
rect 23673 28101 23707 28135
rect 27169 28101 27203 28135
rect 28457 28101 28491 28135
rect 28549 28101 28583 28135
rect 30389 28101 30423 28135
rect 34130 28101 34164 28135
rect 37841 28101 37875 28135
rect 4905 28033 4939 28067
rect 5181 28033 5215 28067
rect 8309 28033 8343 28067
rect 8585 28033 8619 28067
rect 9137 28033 9171 28067
rect 9413 28033 9447 28067
rect 9965 28033 9999 28067
rect 10241 28033 10275 28067
rect 10977 28033 11011 28067
rect 11161 28033 11195 28067
rect 12725 28033 12759 28067
rect 13185 28033 13219 28067
rect 13461 28033 13495 28067
rect 14013 28033 14047 28067
rect 14289 28033 14323 28067
rect 14381 28033 14415 28067
rect 16865 28033 16899 28067
rect 17049 28033 17083 28067
rect 18889 28033 18923 28067
rect 19073 28033 19107 28067
rect 20085 28033 20119 28067
rect 22109 28033 22143 28067
rect 24593 28033 24627 28067
rect 25513 28033 25547 28067
rect 25697 28033 25731 28067
rect 27629 28033 27663 28067
rect 28273 28033 28307 28067
rect 28693 28033 28727 28067
rect 30113 28033 30147 28067
rect 30206 28033 30240 28067
rect 30481 28033 30515 28067
rect 30578 28033 30612 28067
rect 33885 28033 33919 28067
rect 36093 28033 36127 28067
rect 5089 27965 5123 27999
rect 6929 27965 6963 27999
rect 10149 27965 10183 27999
rect 20177 27965 20211 27999
rect 22477 27965 22511 27999
rect 24777 27965 24811 27999
rect 27445 27965 27479 27999
rect 38025 27965 38059 27999
rect 7481 27897 7515 27931
rect 8401 27897 8435 27931
rect 10425 27897 10459 27931
rect 19165 27897 19199 27931
rect 24041 27897 24075 27931
rect 4997 27829 5031 27863
rect 5365 27829 5399 27863
rect 7297 27829 7331 27863
rect 9229 27829 9263 27863
rect 10241 27829 10275 27863
rect 14565 27829 14599 27863
rect 20085 27829 20119 27863
rect 20453 27829 20487 27863
rect 27445 27829 27479 27863
rect 27813 27829 27847 27863
rect 28825 27829 28859 27863
rect 35265 27829 35299 27863
rect 13277 27625 13311 27659
rect 31493 27625 31527 27659
rect 4261 27557 4295 27591
rect 7021 27557 7055 27591
rect 9965 27557 9999 27591
rect 13737 27557 13771 27591
rect 15669 27557 15703 27591
rect 17325 27557 17359 27591
rect 24041 27557 24075 27591
rect 4353 27489 4387 27523
rect 5365 27489 5399 27523
rect 8033 27489 8067 27523
rect 8125 27489 8159 27523
rect 8217 27489 8251 27523
rect 18245 27489 18279 27523
rect 26249 27489 26283 27523
rect 29929 27489 29963 27523
rect 4169 27421 4203 27455
rect 4445 27421 4479 27455
rect 4629 27421 4663 27455
rect 5089 27421 5123 27455
rect 5273 27421 5307 27455
rect 5457 27421 5491 27455
rect 5641 27421 5675 27455
rect 6745 27421 6779 27455
rect 7021 27421 7055 27455
rect 8309 27421 8343 27455
rect 10425 27421 10459 27455
rect 11161 27421 11195 27455
rect 11345 27421 11379 27455
rect 13185 27421 13219 27455
rect 13553 27421 13587 27455
rect 14289 27421 14323 27455
rect 14556 27421 14590 27455
rect 17509 27421 17543 27455
rect 17601 27421 17635 27455
rect 18153 27421 18187 27455
rect 19441 27421 19475 27455
rect 20177 27421 20211 27455
rect 21097 27421 21131 27455
rect 22753 27421 22787 27455
rect 23489 27421 23523 27455
rect 26525 27421 26559 27455
rect 26614 27415 26648 27449
rect 26709 27421 26743 27455
rect 26893 27421 26927 27455
rect 27629 27421 27663 27455
rect 27721 27421 27755 27455
rect 27813 27421 27847 27455
rect 27997 27421 28031 27455
rect 28825 27421 28859 27455
rect 30021 27421 30055 27455
rect 30389 27421 30423 27455
rect 30849 27421 30883 27455
rect 30942 27421 30976 27455
rect 31125 27421 31159 27455
rect 31314 27421 31348 27455
rect 31953 27421 31987 27455
rect 32321 27421 32355 27455
rect 32965 27421 32999 27455
rect 33149 27421 33183 27455
rect 36921 27421 36955 27455
rect 37841 27421 37875 27455
rect 9597 27353 9631 27387
rect 9781 27353 9815 27387
rect 19993 27353 20027 27387
rect 21649 27353 21683 27387
rect 23213 27353 23247 27387
rect 28641 27353 28675 27387
rect 29193 27353 29227 27387
rect 30297 27353 30331 27387
rect 31217 27353 31251 27387
rect 32137 27353 32171 27387
rect 32229 27353 32263 27387
rect 37197 27353 37231 27387
rect 38117 27353 38151 27387
rect 3985 27285 4019 27319
rect 5825 27285 5859 27319
rect 7849 27285 7883 27319
rect 10609 27285 10643 27319
rect 11253 27285 11287 27319
rect 19625 27285 19659 27319
rect 20085 27285 20119 27319
rect 27353 27285 27387 27319
rect 29745 27285 29779 27319
rect 32505 27285 32539 27319
rect 33057 27285 33091 27319
rect 4169 27081 4203 27115
rect 20085 27081 20119 27115
rect 22477 27081 22511 27115
rect 24777 27081 24811 27115
rect 26341 27081 26375 27115
rect 29101 27081 29135 27115
rect 36185 27081 36219 27115
rect 37933 27081 37967 27115
rect 3056 27013 3090 27047
rect 5089 27013 5123 27047
rect 22017 27013 22051 27047
rect 26157 27013 26191 27047
rect 32956 27013 32990 27047
rect 37841 27013 37875 27047
rect 2789 26945 2823 26979
rect 5549 26945 5583 26979
rect 7021 26945 7055 26979
rect 8493 26945 8527 26979
rect 8585 26945 8619 26979
rect 9229 26945 9263 26979
rect 9413 26945 9447 26979
rect 10793 26945 10827 26979
rect 13369 26945 13403 26979
rect 13553 26945 13587 26979
rect 13645 26945 13679 26979
rect 14381 26945 14415 26979
rect 17049 26945 17083 26979
rect 17325 26945 17359 26979
rect 17877 26945 17911 26979
rect 18153 26945 18187 26979
rect 18889 26945 18923 26979
rect 19257 26945 19291 26979
rect 19993 26945 20027 26979
rect 20177 26945 20211 26979
rect 20821 26945 20855 26979
rect 22293 26945 22327 26979
rect 22937 26945 22971 26979
rect 23213 26945 23247 26979
rect 24593 26945 24627 26979
rect 24777 26945 24811 26979
rect 27261 26945 27295 26979
rect 28089 26945 28123 26979
rect 29101 26945 29135 26979
rect 29745 26945 29779 26979
rect 31033 26945 31067 26979
rect 31125 26945 31159 26979
rect 31309 26945 31343 26979
rect 31401 26945 31435 26979
rect 32689 26945 32723 26979
rect 35173 26945 35207 26979
rect 35357 26945 35391 26979
rect 35449 26945 35483 26979
rect 35541 26945 35575 26979
rect 36369 26945 36403 26979
rect 36645 26945 36679 26979
rect 5365 26877 5399 26911
rect 6837 26877 6871 26911
rect 10885 26877 10919 26911
rect 10977 26877 11011 26911
rect 14657 26877 14691 26911
rect 17233 26877 17267 26911
rect 19073 26877 19107 26911
rect 20913 26877 20947 26911
rect 22109 26877 22143 26911
rect 23029 26877 23063 26911
rect 38025 26877 38059 26911
rect 5733 26809 5767 26843
rect 7205 26809 7239 26843
rect 8677 26809 8711 26843
rect 17141 26809 17175 26843
rect 18153 26809 18187 26843
rect 19165 26809 19199 26843
rect 21189 26809 21223 26843
rect 26525 26809 26559 26843
rect 34069 26809 34103 26843
rect 5549 26741 5583 26775
rect 9229 26741 9263 26775
rect 10425 26741 10459 26775
rect 13185 26741 13219 26775
rect 16865 26741 16899 26775
rect 19073 26741 19107 26775
rect 21005 26741 21039 26775
rect 22293 26741 22327 26775
rect 23121 26741 23155 26775
rect 23397 26741 23431 26775
rect 26341 26741 26375 26775
rect 28273 26741 28307 26775
rect 30849 26741 30883 26775
rect 35725 26741 35759 26775
rect 36553 26741 36587 26775
rect 37473 26741 37507 26775
rect 4905 26537 4939 26571
rect 6009 26537 6043 26571
rect 9137 26537 9171 26571
rect 11989 26537 12023 26571
rect 13277 26537 13311 26571
rect 22293 26537 22327 26571
rect 22753 26537 22787 26571
rect 27537 26537 27571 26571
rect 35265 26537 35299 26571
rect 38117 26537 38151 26571
rect 34253 26469 34287 26503
rect 4353 26401 4387 26435
rect 5089 26401 5123 26435
rect 10609 26401 10643 26435
rect 15669 26401 15703 26435
rect 24869 26401 24903 26435
rect 27997 26401 28031 26435
rect 28549 26401 28583 26435
rect 31217 26401 31251 26435
rect 32229 26401 32263 26435
rect 4261 26333 4295 26367
rect 4445 26333 4479 26367
rect 5181 26333 5215 26367
rect 5273 26333 5307 26367
rect 5365 26333 5399 26367
rect 6285 26333 6319 26367
rect 6745 26333 6779 26367
rect 6929 26333 6963 26367
rect 9321 26333 9355 26367
rect 9505 26333 9539 26367
rect 9781 26333 9815 26367
rect 10876 26333 10910 26367
rect 13461 26333 13495 26367
rect 13737 26333 13771 26367
rect 15577 26333 15611 26367
rect 15945 26333 15979 26367
rect 16037 26333 16071 26367
rect 16865 26333 16899 26367
rect 17141 26333 17175 26367
rect 17417 26333 17451 26367
rect 17785 26333 17819 26367
rect 20637 26333 20671 26367
rect 20821 26333 20855 26367
rect 21281 26333 21315 26367
rect 21465 26333 21499 26367
rect 21741 26333 21775 26367
rect 22293 26333 22327 26367
rect 22477 26333 22511 26367
rect 22569 26333 22603 26367
rect 23213 26333 23247 26367
rect 23397 26333 23431 26367
rect 24593 26333 24627 26367
rect 24781 26335 24815 26369
rect 24961 26333 24995 26367
rect 25145 26333 25179 26367
rect 27169 26333 27203 26367
rect 28181 26333 28215 26367
rect 31861 26333 31895 26367
rect 33149 26333 33183 26367
rect 33241 26333 33275 26367
rect 33425 26333 33459 26367
rect 33517 26333 33551 26367
rect 33977 26333 34011 26367
rect 34161 26333 34195 26367
rect 35449 26333 35483 26367
rect 35541 26333 35575 26367
rect 35725 26333 35759 26367
rect 35817 26333 35851 26367
rect 36737 26333 36771 26367
rect 37004 26333 37038 26367
rect 6009 26265 6043 26299
rect 6193 26265 6227 26299
rect 6837 26265 6871 26299
rect 9413 26265 9447 26299
rect 9623 26265 9657 26299
rect 13645 26265 13679 26299
rect 14933 26265 14967 26299
rect 25789 26265 25823 26299
rect 25973 26265 26007 26299
rect 27353 26265 27387 26299
rect 31033 26265 31067 26299
rect 32965 26265 32999 26299
rect 17785 26197 17819 26231
rect 20729 26197 20763 26231
rect 21649 26197 21683 26231
rect 23489 26197 23523 26231
rect 25329 26197 25363 26231
rect 26157 26197 26191 26231
rect 28457 26197 28491 26231
rect 30573 26197 30607 26231
rect 30941 26197 30975 26231
rect 5457 25993 5491 26027
rect 8049 25993 8083 26027
rect 8217 25993 8251 26027
rect 14565 25993 14599 26027
rect 18153 25993 18187 26027
rect 22569 25993 22603 26027
rect 24501 25993 24535 26027
rect 33333 25993 33367 26027
rect 6561 25925 6595 25959
rect 7849 25925 7883 25959
rect 13430 25925 13464 25959
rect 17141 25925 17175 25959
rect 30757 25925 30791 25959
rect 5273 25857 5307 25891
rect 5549 25857 5583 25891
rect 6745 25857 6779 25891
rect 6837 25857 6871 25891
rect 10149 25857 10183 25891
rect 10333 25857 10367 25891
rect 16957 25857 16991 25891
rect 18337 25857 18371 25891
rect 18613 25857 18647 25891
rect 19441 25857 19475 25891
rect 20637 25857 20671 25891
rect 20821 25857 20855 25891
rect 21189 25857 21223 25891
rect 23121 25857 23155 25891
rect 23673 25857 23707 25891
rect 24685 25857 24719 25891
rect 24961 25857 24995 25891
rect 25145 25857 25179 25891
rect 27537 25857 27571 25891
rect 27721 25857 27755 25891
rect 27813 25857 27847 25891
rect 27905 25857 27939 25891
rect 28549 25857 28583 25891
rect 33149 25857 33183 25891
rect 37841 25857 37875 25891
rect 13185 25789 13219 25823
rect 19625 25789 19659 25823
rect 19901 25789 19935 25823
rect 19993 25789 20027 25823
rect 29009 25789 29043 25823
rect 31585 25789 31619 25823
rect 32965 25789 32999 25823
rect 38117 25789 38151 25823
rect 5089 25721 5123 25755
rect 24777 25721 24811 25755
rect 24869 25721 24903 25755
rect 4813 25653 4847 25687
rect 5181 25653 5215 25687
rect 6561 25653 6595 25687
rect 8033 25653 8067 25687
rect 10149 25653 10183 25687
rect 17233 25653 17267 25687
rect 28089 25653 28123 25687
rect 6285 25449 6319 25483
rect 9321 25449 9355 25483
rect 12909 25449 12943 25483
rect 21925 25449 21959 25483
rect 27629 25449 27663 25483
rect 7941 25381 7975 25415
rect 16589 25381 16623 25415
rect 26065 25381 26099 25415
rect 28641 25381 28675 25415
rect 32873 25381 32907 25415
rect 4353 25313 4387 25347
rect 4905 25313 4939 25347
rect 5273 25313 5307 25347
rect 6469 25313 6503 25347
rect 6561 25313 6595 25347
rect 18337 25313 18371 25347
rect 25513 25313 25547 25347
rect 30021 25313 30055 25347
rect 34069 25313 34103 25347
rect 34345 25313 34379 25347
rect 4169 25245 4203 25279
rect 4445 25245 4479 25279
rect 5365 25245 5399 25279
rect 6653 25245 6687 25279
rect 6745 25245 6779 25279
rect 8125 25245 8159 25279
rect 8401 25245 8435 25279
rect 10517 25245 10551 25279
rect 10701 25245 10735 25279
rect 10793 25245 10827 25279
rect 10885 25245 10919 25279
rect 11529 25245 11563 25279
rect 14289 25245 14323 25279
rect 14657 25245 14691 25279
rect 16773 25245 16807 25279
rect 18521 25245 18555 25279
rect 18889 25245 18923 25279
rect 19533 25245 19567 25279
rect 19625 25245 19659 25279
rect 20637 25245 20671 25279
rect 21005 25245 21039 25279
rect 21649 25245 21683 25279
rect 21833 25245 21867 25279
rect 22753 25245 22787 25279
rect 22937 25245 22971 25279
rect 24961 25245 24995 25279
rect 25145 25245 25179 25279
rect 25973 25245 26007 25279
rect 26525 25245 26559 25279
rect 26801 25245 26835 25279
rect 27537 25245 27571 25279
rect 28457 25245 28491 25279
rect 28549 25245 28583 25279
rect 28733 25245 28767 25279
rect 32413 25245 32447 25279
rect 32597 25245 32631 25279
rect 32965 25245 32999 25279
rect 33977 25245 34011 25279
rect 34897 25245 34931 25279
rect 36829 25245 36863 25279
rect 9137 25177 9171 25211
rect 11774 25177 11808 25211
rect 14473 25177 14507 25211
rect 14565 25177 14599 25211
rect 16865 25177 16899 25211
rect 30288 25177 30322 25211
rect 35142 25177 35176 25211
rect 37096 25177 37130 25211
rect 3985 25109 4019 25143
rect 5549 25109 5583 25143
rect 9321 25109 9355 25143
rect 9505 25109 9539 25143
rect 11069 25109 11103 25143
rect 14841 25109 14875 25143
rect 16957 25109 16991 25143
rect 17141 25109 17175 25143
rect 18797 25109 18831 25143
rect 19533 25109 19567 25143
rect 20545 25109 20579 25143
rect 23029 25109 23063 25143
rect 28273 25109 28307 25143
rect 31401 25109 31435 25143
rect 36277 25109 36311 25143
rect 38209 25109 38243 25143
rect 4721 24905 4755 24939
rect 5917 24905 5951 24939
rect 23765 24905 23799 24939
rect 23857 24905 23891 24939
rect 32965 24905 32999 24939
rect 33885 24905 33919 24939
rect 37473 24905 37507 24939
rect 37841 24905 37875 24939
rect 2964 24837 2998 24871
rect 33517 24837 33551 24871
rect 36093 24837 36127 24871
rect 2697 24769 2731 24803
rect 4905 24769 4939 24803
rect 4997 24769 5031 24803
rect 5181 24769 5215 24803
rect 5825 24769 5859 24803
rect 6009 24769 6043 24803
rect 6561 24769 6595 24803
rect 6745 24769 6779 24803
rect 6929 24769 6963 24803
rect 7665 24769 7699 24803
rect 7849 24769 7883 24803
rect 9597 24769 9631 24803
rect 9873 24769 9907 24803
rect 10517 24769 10551 24803
rect 10701 24769 10735 24803
rect 10793 24769 10827 24803
rect 10885 24769 10919 24803
rect 14381 24769 14415 24803
rect 16865 24769 16899 24803
rect 17693 24769 17727 24803
rect 17877 24769 17911 24803
rect 18521 24769 18555 24803
rect 19165 24769 19199 24803
rect 19441 24769 19475 24803
rect 19625 24769 19659 24803
rect 20269 24769 20303 24803
rect 22753 24769 22787 24803
rect 23029 24769 23063 24803
rect 23933 24769 23967 24803
rect 25237 24769 25271 24803
rect 25513 24769 25547 24803
rect 27629 24769 27663 24803
rect 29009 24769 29043 24803
rect 29193 24769 29227 24803
rect 29285 24769 29319 24803
rect 29745 24769 29779 24803
rect 30021 24769 30055 24803
rect 32321 24769 32355 24803
rect 32414 24769 32448 24803
rect 32597 24769 32631 24803
rect 32686 24769 32720 24803
rect 32786 24769 32820 24803
rect 33701 24769 33735 24803
rect 34345 24769 34379 24803
rect 34529 24769 34563 24803
rect 34621 24769 34655 24803
rect 35265 24769 35299 24803
rect 5089 24701 5123 24735
rect 9689 24701 9723 24735
rect 14105 24701 14139 24735
rect 19349 24701 19383 24735
rect 20545 24701 20579 24735
rect 23581 24701 23615 24735
rect 24317 24701 24351 24735
rect 25697 24701 25731 24735
rect 28457 24701 28491 24735
rect 30481 24701 30515 24735
rect 37933 24701 37967 24735
rect 38025 24701 38059 24735
rect 18429 24633 18463 24667
rect 19257 24633 19291 24667
rect 29009 24633 29043 24667
rect 29837 24633 29871 24667
rect 34345 24633 34379 24667
rect 4077 24565 4111 24599
rect 7665 24565 7699 24599
rect 9873 24565 9907 24599
rect 10057 24565 10091 24599
rect 11069 24565 11103 24599
rect 15669 24565 15703 24599
rect 18981 24565 19015 24599
rect 22569 24565 22603 24599
rect 22937 24565 22971 24599
rect 6837 24361 6871 24395
rect 9505 24361 9539 24395
rect 12081 24361 12115 24395
rect 23857 24361 23891 24395
rect 27905 24361 27939 24395
rect 33609 24361 33643 24395
rect 7941 24293 7975 24327
rect 20085 24293 20119 24327
rect 20177 24293 20211 24327
rect 24869 24293 24903 24327
rect 8493 24225 8527 24259
rect 10701 24225 10735 24259
rect 16773 24225 16807 24259
rect 30021 24225 30055 24259
rect 30665 24225 30699 24259
rect 6653 24157 6687 24191
rect 10968 24157 11002 24191
rect 14289 24157 14323 24191
rect 14545 24157 14579 24191
rect 17141 24157 17175 24191
rect 17325 24157 17359 24191
rect 17509 24157 17543 24191
rect 17693 24157 17727 24191
rect 18705 24157 18739 24191
rect 19993 24157 20027 24191
rect 20269 24157 20303 24191
rect 21005 24157 21039 24191
rect 22661 24157 22695 24191
rect 22845 24157 22879 24191
rect 23029 24157 23063 24191
rect 23305 24157 23339 24191
rect 23857 24157 23891 24191
rect 24041 24157 24075 24191
rect 24685 24157 24719 24191
rect 24777 24157 24811 24191
rect 25973 24157 26007 24191
rect 26157 24157 26191 24191
rect 26341 24157 26375 24191
rect 27261 24157 27295 24191
rect 27409 24157 27443 24191
rect 27767 24157 27801 24191
rect 29929 24157 29963 24191
rect 30205 24157 30239 24191
rect 31861 24157 31895 24191
rect 31954 24157 31988 24191
rect 32137 24157 32171 24191
rect 32365 24157 32399 24191
rect 32965 24157 32999 24191
rect 33113 24157 33147 24191
rect 33430 24157 33464 24191
rect 37841 24157 37875 24191
rect 8217 24089 8251 24123
rect 9321 24089 9355 24123
rect 9505 24089 9539 24123
rect 20821 24089 20855 24123
rect 26249 24089 26283 24123
rect 27537 24089 27571 24123
rect 27629 24089 27663 24123
rect 32229 24089 32263 24123
rect 33241 24089 33275 24123
rect 33333 24089 33367 24123
rect 38117 24089 38151 24123
rect 8125 24021 8159 24055
rect 8309 24021 8343 24055
rect 9689 24021 9723 24055
rect 15669 24021 15703 24055
rect 18153 24021 18187 24055
rect 18797 24021 18831 24055
rect 19809 24021 19843 24055
rect 21097 24021 21131 24055
rect 22661 24021 22695 24055
rect 26525 24021 26559 24055
rect 32505 24021 32539 24055
rect 4077 23817 4111 23851
rect 21097 23817 21131 23851
rect 7297 23749 7331 23783
rect 19717 23749 19751 23783
rect 24869 23749 24903 23783
rect 25237 23749 25271 23783
rect 27169 23749 27203 23783
rect 28641 23749 28675 23783
rect 30665 23749 30699 23783
rect 35081 23749 35115 23783
rect 35173 23749 35207 23783
rect 35909 23749 35943 23783
rect 37933 23749 37967 23783
rect 2697 23681 2731 23715
rect 2964 23681 2998 23715
rect 4721 23681 4755 23715
rect 4813 23681 4847 23715
rect 4997 23681 5031 23715
rect 5089 23681 5123 23715
rect 5549 23681 5583 23715
rect 5733 23681 5767 23715
rect 6009 23681 6043 23715
rect 7113 23681 7147 23715
rect 7389 23681 7423 23715
rect 8401 23681 8435 23715
rect 9321 23681 9355 23715
rect 10425 23681 10459 23715
rect 19901 23681 19935 23715
rect 21005 23681 21039 23715
rect 23213 23681 23247 23715
rect 23397 23681 23431 23715
rect 23765 23681 23799 23715
rect 25053 23681 25087 23715
rect 25697 23681 25731 23715
rect 26249 23681 26283 23715
rect 27353 23681 27387 23715
rect 27629 23681 27663 23715
rect 28365 23681 28399 23715
rect 28503 23681 28537 23715
rect 28757 23681 28791 23715
rect 29929 23681 29963 23715
rect 30205 23681 30239 23715
rect 32597 23681 32631 23715
rect 32689 23681 32723 23715
rect 32965 23681 32999 23715
rect 34805 23681 34839 23715
rect 34898 23681 34932 23715
rect 35270 23681 35304 23715
rect 36093 23681 36127 23715
rect 36185 23681 36219 23715
rect 36461 23681 36495 23715
rect 37841 23681 37875 23715
rect 9505 23613 9539 23647
rect 10241 23613 10275 23647
rect 21281 23613 21315 23647
rect 26065 23613 26099 23647
rect 26157 23613 26191 23647
rect 36369 23613 36403 23647
rect 38025 23613 38059 23647
rect 23673 23545 23707 23579
rect 30021 23545 30055 23579
rect 32413 23545 32447 23579
rect 35449 23545 35483 23579
rect 4537 23477 4571 23511
rect 5917 23477 5951 23511
rect 6929 23477 6963 23511
rect 8493 23477 8527 23511
rect 10609 23477 10643 23511
rect 20085 23477 20119 23511
rect 20637 23477 20671 23511
rect 27537 23477 27571 23511
rect 28917 23477 28951 23511
rect 32873 23477 32907 23511
rect 37473 23477 37507 23511
rect 3985 23273 4019 23307
rect 10517 23273 10551 23307
rect 21281 23273 21315 23307
rect 22569 23273 22603 23307
rect 34989 23273 35023 23307
rect 38117 23273 38151 23307
rect 6929 23205 6963 23239
rect 15301 23205 15335 23239
rect 23121 23205 23155 23239
rect 4537 23137 4571 23171
rect 6837 23137 6871 23171
rect 20545 23137 20579 23171
rect 20637 23137 20671 23171
rect 21833 23137 21867 23171
rect 26709 23137 26743 23171
rect 35633 23137 35667 23171
rect 4353 23069 4387 23103
rect 4445 23069 4479 23103
rect 5825 23069 5859 23103
rect 6745 23069 6779 23103
rect 7021 23069 7055 23103
rect 7757 23069 7791 23103
rect 8033 23069 8067 23103
rect 9137 23069 9171 23103
rect 12081 23069 12115 23103
rect 14657 23069 14691 23103
rect 15577 23069 15611 23103
rect 16037 23069 16071 23103
rect 16957 23069 16991 23103
rect 22477 23069 22511 23103
rect 22753 23069 22787 23103
rect 22937 23069 22971 23103
rect 25973 23069 26007 23103
rect 26617 23069 26651 23103
rect 26893 23069 26927 23103
rect 27813 23069 27847 23103
rect 27997 23069 28031 23103
rect 28457 23069 28491 23103
rect 28605 23069 28639 23103
rect 28733 23069 28767 23103
rect 28922 23069 28956 23103
rect 29837 23069 29871 23103
rect 30297 23069 30331 23103
rect 30665 23069 30699 23103
rect 35173 23069 35207 23103
rect 35265 23069 35299 23103
rect 35541 23069 35575 23103
rect 36737 23069 36771 23103
rect 37004 23069 37038 23103
rect 5917 23001 5951 23035
rect 9382 23001 9416 23035
rect 12348 23001 12382 23035
rect 15301 23001 15335 23035
rect 17224 23001 17258 23035
rect 21741 23001 21775 23035
rect 27905 23001 27939 23035
rect 28825 23001 28859 23035
rect 6561 22933 6595 22967
rect 7573 22933 7607 22967
rect 7941 22933 7975 22967
rect 13461 22933 13495 22967
rect 14749 22933 14783 22967
rect 15485 22933 15519 22967
rect 16129 22933 16163 22967
rect 18337 22933 18371 22967
rect 20085 22933 20119 22967
rect 20453 22933 20487 22967
rect 21649 22933 21683 22967
rect 29101 22933 29135 22967
rect 30941 22933 30975 22967
rect 4813 22729 4847 22763
rect 8953 22729 8987 22763
rect 12357 22729 12391 22763
rect 15669 22729 15703 22763
rect 21189 22729 21223 22763
rect 28273 22729 28307 22763
rect 33517 22729 33551 22763
rect 7205 22661 7239 22695
rect 11069 22661 11103 22695
rect 12081 22661 12115 22695
rect 15945 22661 15979 22695
rect 16155 22661 16189 22695
rect 16865 22661 16899 22695
rect 19165 22661 19199 22695
rect 20076 22661 20110 22695
rect 29561 22661 29595 22695
rect 29653 22661 29687 22695
rect 31769 22661 31803 22695
rect 35817 22661 35851 22695
rect 4721 22593 4755 22627
rect 4905 22593 4939 22627
rect 7481 22593 7515 22627
rect 9137 22593 9171 22627
rect 9413 22593 9447 22627
rect 10885 22593 10919 22627
rect 11161 22593 11195 22627
rect 11805 22593 11839 22627
rect 11989 22593 12023 22627
rect 12173 22593 12207 22627
rect 14381 22593 14415 22627
rect 14565 22593 14599 22627
rect 15025 22593 15059 22627
rect 15853 22593 15887 22627
rect 16038 22593 16072 22627
rect 17049 22593 17083 22627
rect 18337 22593 18371 22627
rect 19809 22593 19843 22627
rect 22661 22593 22695 22627
rect 22937 22593 22971 22627
rect 23581 22593 23615 22627
rect 24501 22593 24535 22627
rect 24869 22593 24903 22627
rect 27629 22593 27663 22627
rect 27722 22593 27756 22627
rect 27905 22593 27939 22627
rect 27997 22593 28031 22627
rect 28135 22593 28169 22627
rect 29377 22593 29411 22627
rect 29745 22593 29779 22627
rect 31217 22593 31251 22627
rect 31585 22593 31619 22627
rect 33149 22593 33183 22627
rect 33333 22593 33367 22627
rect 35449 22593 35483 22627
rect 35725 22593 35759 22627
rect 37841 22593 37875 22627
rect 7297 22525 7331 22559
rect 9229 22525 9263 22559
rect 9321 22525 9355 22559
rect 16313 22525 16347 22559
rect 17417 22525 17451 22559
rect 18521 22525 18555 22559
rect 23397 22525 23431 22559
rect 25329 22525 25363 22559
rect 30757 22525 30791 22559
rect 35357 22525 35391 22559
rect 38117 22525 38151 22559
rect 24409 22457 24443 22491
rect 7205 22389 7239 22423
rect 7665 22389 7699 22423
rect 10701 22389 10735 22423
rect 14473 22389 14507 22423
rect 15117 22389 15151 22423
rect 29929 22389 29963 22423
rect 35173 22389 35207 22423
rect 7205 22185 7239 22219
rect 11897 22185 11931 22219
rect 15117 22185 15151 22219
rect 16405 22185 16439 22219
rect 27905 22185 27939 22219
rect 23305 22117 23339 22151
rect 4629 22049 4663 22083
rect 15761 22049 15795 22083
rect 23029 22049 23063 22083
rect 25789 22049 25823 22083
rect 31217 22049 31251 22083
rect 31309 22049 31343 22083
rect 33793 22049 33827 22083
rect 34253 22049 34287 22083
rect 4445 21981 4479 22015
rect 7481 21981 7515 22015
rect 7573 21981 7607 22015
rect 7665 21981 7699 22015
rect 7849 21981 7883 22015
rect 9229 21981 9263 22015
rect 9321 21981 9355 22015
rect 10517 21981 10551 22015
rect 12357 21981 12391 22015
rect 14289 21981 14323 22015
rect 14473 21981 14507 22015
rect 15301 21981 15335 22015
rect 15485 21981 15519 22015
rect 16221 21981 16255 22015
rect 16405 21981 16439 22015
rect 22937 21981 22971 22015
rect 23857 21981 23891 22015
rect 24041 21981 24075 22015
rect 24869 21981 24903 22015
rect 25329 21981 25363 22015
rect 26801 21981 26835 22015
rect 27169 21981 27203 22015
rect 27905 21981 27939 22015
rect 28089 21981 28123 22015
rect 30849 21981 30883 22015
rect 30941 21981 30975 22015
rect 32597 21981 32631 22015
rect 32745 21981 32779 22015
rect 33062 21981 33096 22015
rect 33885 21981 33919 22015
rect 34897 21981 34931 22015
rect 36921 21981 36955 22015
rect 9505 21913 9539 21947
rect 10762 21913 10796 21947
rect 12602 21913 12636 21947
rect 14657 21913 14691 21947
rect 15393 21913 15427 21947
rect 15623 21913 15657 21947
rect 26985 21913 27019 21947
rect 27077 21913 27111 21947
rect 32873 21913 32907 21947
rect 32965 21913 32999 21947
rect 35142 21913 35176 21947
rect 37188 21913 37222 21947
rect 3985 21845 4019 21879
rect 4353 21845 4387 21879
rect 13737 21845 13771 21879
rect 16589 21845 16623 21879
rect 23949 21845 23983 21879
rect 24869 21845 24903 21879
rect 27353 21845 27387 21879
rect 30665 21845 30699 21879
rect 33241 21845 33275 21879
rect 36277 21845 36311 21879
rect 38301 21845 38335 21879
rect 9255 21641 9289 21675
rect 9873 21641 9907 21675
rect 26525 21641 26559 21675
rect 32873 21641 32907 21675
rect 35633 21641 35667 21675
rect 37473 21641 37507 21675
rect 3056 21573 3090 21607
rect 6837 21573 6871 21607
rect 9045 21573 9079 21607
rect 10149 21573 10183 21607
rect 22293 21573 22327 21607
rect 27445 21573 27479 21607
rect 28641 21573 28675 21607
rect 32689 21573 32723 21607
rect 35357 21573 35391 21607
rect 36093 21573 36127 21607
rect 37933 21573 37967 21607
rect 2789 21505 2823 21539
rect 5733 21505 5767 21539
rect 6561 21505 6595 21539
rect 6745 21505 6779 21539
rect 6929 21505 6963 21539
rect 7849 21505 7883 21539
rect 9873 21505 9907 21539
rect 14749 21505 14783 21539
rect 15025 21505 15059 21539
rect 15853 21505 15887 21539
rect 15945 21505 15979 21539
rect 16865 21505 16899 21539
rect 22017 21505 22051 21539
rect 22201 21505 22235 21539
rect 22390 21505 22424 21539
rect 24777 21505 24811 21539
rect 26341 21505 26375 21539
rect 26617 21505 26651 21539
rect 27169 21505 27203 21539
rect 27353 21505 27387 21539
rect 27537 21505 27571 21539
rect 28365 21505 28399 21539
rect 28513 21505 28547 21539
rect 28733 21505 28767 21539
rect 28830 21505 28864 21539
rect 30481 21505 30515 21539
rect 30757 21505 30791 21539
rect 31217 21505 31251 21539
rect 31585 21505 31619 21539
rect 32965 21505 32999 21539
rect 34989 21505 35023 21539
rect 35082 21505 35116 21539
rect 35265 21505 35299 21539
rect 35495 21505 35529 21539
rect 36277 21505 36311 21539
rect 36369 21505 36403 21539
rect 36645 21505 36679 21539
rect 37841 21505 37875 21539
rect 5549 21437 5583 21471
rect 5917 21437 5951 21471
rect 7941 21437 7975 21471
rect 8033 21437 8067 21471
rect 8125 21437 8159 21471
rect 9965 21437 9999 21471
rect 14933 21437 14967 21471
rect 16221 21437 16255 21471
rect 16313 21437 16347 21471
rect 17601 21437 17635 21471
rect 26157 21437 26191 21471
rect 31033 21437 31067 21471
rect 38025 21437 38059 21471
rect 4169 21369 4203 21403
rect 22569 21369 22603 21403
rect 32689 21369 32723 21403
rect 36553 21369 36587 21403
rect 7113 21301 7147 21335
rect 7665 21301 7699 21335
rect 9229 21301 9263 21335
rect 9413 21301 9447 21335
rect 14749 21301 14783 21335
rect 15209 21301 15243 21335
rect 15669 21301 15703 21335
rect 25053 21301 25087 21335
rect 27721 21301 27755 21335
rect 29009 21301 29043 21335
rect 5917 21097 5951 21131
rect 10977 21097 11011 21131
rect 18521 21097 18555 21131
rect 21833 21097 21867 21131
rect 31585 21097 31619 21131
rect 31953 21097 31987 21131
rect 32597 21029 32631 21063
rect 4537 20961 4571 20995
rect 14933 20961 14967 20995
rect 31677 20961 31711 20995
rect 4804 20893 4838 20927
rect 6837 20893 6871 20927
rect 7113 20893 7147 20927
rect 9597 20893 9631 20927
rect 15485 20893 15519 20927
rect 17601 20893 17635 20927
rect 20545 20893 20579 20927
rect 24593 20893 24627 20927
rect 24869 20893 24903 20927
rect 25053 20893 25087 20927
rect 25329 20893 25363 20927
rect 25522 20893 25556 20927
rect 27261 20893 27295 20927
rect 27353 20893 27387 20927
rect 27537 20893 27571 20927
rect 27629 20893 27663 20927
rect 29745 20893 29779 20927
rect 29929 20893 29963 20927
rect 31309 20893 31343 20927
rect 31456 20893 31490 20927
rect 32873 20893 32907 20927
rect 36737 20893 36771 20927
rect 9864 20825 9898 20859
rect 14657 20825 14691 20859
rect 15761 20825 15795 20859
rect 17233 20825 17267 20859
rect 17509 20825 17543 20859
rect 17969 20825 18003 20859
rect 18337 20825 18371 20859
rect 26157 20825 26191 20859
rect 32597 20825 32631 20859
rect 37004 20825 37038 20859
rect 6653 20757 6687 20791
rect 7021 20757 7055 20791
rect 14289 20757 14323 20791
rect 14749 20757 14783 20791
rect 27077 20757 27111 20791
rect 29837 20757 29871 20791
rect 32781 20757 32815 20791
rect 38117 20757 38151 20791
rect 4353 20553 4387 20587
rect 9965 20553 9999 20587
rect 13553 20553 13587 20587
rect 14105 20553 14139 20587
rect 18153 20553 18187 20587
rect 23397 20553 23431 20587
rect 24869 20553 24903 20587
rect 27813 20553 27847 20587
rect 33149 20553 33183 20587
rect 33977 20553 34011 20587
rect 37473 20553 37507 20587
rect 9597 20485 9631 20519
rect 9689 20485 9723 20519
rect 12440 20485 12474 20519
rect 15301 20485 15335 20519
rect 28457 20485 28491 20519
rect 29285 20485 29319 20519
rect 32873 20485 32907 20519
rect 33609 20485 33643 20519
rect 4261 20417 4295 20451
rect 6828 20417 6862 20451
rect 9413 20417 9447 20451
rect 9781 20417 9815 20451
rect 14473 20417 14507 20451
rect 15485 20417 15519 20451
rect 15577 20417 15611 20451
rect 15853 20417 15887 20451
rect 17969 20417 18003 20451
rect 19441 20417 19475 20451
rect 19697 20417 19731 20451
rect 22017 20417 22051 20451
rect 22284 20417 22318 20451
rect 24041 20417 24075 20451
rect 25053 20417 25087 20451
rect 25237 20417 25271 20451
rect 25329 20417 25363 20451
rect 25881 20417 25915 20451
rect 26028 20417 26062 20451
rect 28089 20417 28123 20451
rect 29469 20417 29503 20451
rect 29653 20417 29687 20451
rect 29745 20417 29779 20451
rect 30758 20417 30792 20451
rect 32505 20417 32539 20451
rect 32653 20417 32687 20451
rect 32781 20417 32815 20451
rect 33011 20417 33045 20451
rect 33793 20417 33827 20451
rect 35541 20417 35575 20451
rect 35633 20417 35667 20451
rect 35909 20417 35943 20451
rect 37841 20417 37875 20451
rect 4537 20349 4571 20383
rect 6561 20349 6595 20383
rect 12173 20349 12207 20383
rect 14565 20349 14599 20383
rect 14749 20349 14783 20383
rect 15761 20349 15795 20383
rect 18429 20349 18463 20383
rect 18521 20349 18555 20383
rect 23949 20349 23983 20383
rect 26249 20349 26283 20383
rect 27997 20349 28031 20383
rect 28365 20349 28399 20383
rect 31125 20349 31159 20383
rect 31217 20349 31251 20383
rect 35357 20349 35391 20383
rect 37933 20349 37967 20383
rect 38025 20349 38059 20383
rect 20821 20281 20855 20315
rect 24409 20281 24443 20315
rect 35817 20281 35851 20315
rect 3893 20213 3927 20247
rect 7941 20213 7975 20247
rect 26157 20213 26191 20247
rect 26525 20213 26559 20247
rect 30665 20213 30699 20247
rect 7113 20009 7147 20043
rect 12633 20009 12667 20043
rect 14933 20009 14967 20043
rect 16589 20009 16623 20043
rect 24777 20009 24811 20043
rect 29745 20009 29779 20043
rect 36277 20009 36311 20043
rect 5365 19941 5399 19975
rect 20545 19941 20579 19975
rect 23673 19941 23707 19975
rect 30941 19941 30975 19975
rect 3985 19873 4019 19907
rect 15577 19873 15611 19907
rect 16681 19873 16715 19907
rect 19441 19873 19475 19907
rect 21097 19873 21131 19907
rect 29837 19873 29871 19907
rect 31309 19873 31343 19907
rect 33241 19873 33275 19907
rect 33517 19873 33551 19907
rect 38117 19873 38151 19907
rect 4241 19805 4275 19839
rect 6561 19805 6595 19839
rect 6837 19805 6871 19839
rect 6929 19805 6963 19839
rect 8309 19805 8343 19839
rect 8493 19805 8527 19839
rect 10241 19805 10275 19839
rect 10517 19805 10551 19839
rect 10609 19805 10643 19839
rect 11253 19805 11287 19839
rect 16865 19805 16899 19839
rect 17509 19805 17543 19839
rect 19625 19805 19659 19839
rect 19901 19805 19935 19839
rect 20085 19805 20119 19839
rect 20913 19805 20947 19839
rect 21005 19805 21039 19839
rect 22017 19805 22051 19839
rect 22390 19805 22424 19839
rect 23121 19805 23155 19839
rect 23305 19805 23339 19839
rect 23541 19805 23575 19839
rect 24777 19805 24811 19839
rect 24961 19805 24995 19839
rect 27261 19805 27295 19839
rect 27629 19805 27663 19839
rect 29745 19805 29779 19839
rect 31493 19805 31527 19839
rect 33149 19805 33183 19839
rect 34897 19805 34931 19839
rect 37841 19805 37875 19839
rect 6745 19737 6779 19771
rect 10425 19737 10459 19771
rect 11498 19737 11532 19771
rect 15393 19737 15427 19771
rect 16589 19737 16623 19771
rect 18705 19737 18739 19771
rect 22201 19737 22235 19771
rect 22293 19737 22327 19771
rect 23397 19737 23431 19771
rect 27077 19737 27111 19771
rect 35142 19737 35176 19771
rect 8401 19669 8435 19703
rect 10793 19669 10827 19703
rect 15301 19669 15335 19703
rect 17049 19669 17083 19703
rect 22577 19669 22611 19703
rect 30113 19669 30147 19703
rect 31401 19669 31435 19703
rect 15301 19465 15335 19499
rect 17417 19465 17451 19499
rect 19349 19465 19383 19499
rect 19809 19465 19843 19499
rect 35541 19465 35575 19499
rect 5457 19397 5491 19431
rect 8217 19397 8251 19431
rect 8309 19397 8343 19431
rect 19717 19397 19751 19431
rect 20729 19397 20763 19431
rect 20913 19397 20947 19431
rect 26249 19397 26283 19431
rect 29009 19397 29043 19431
rect 29101 19397 29135 19431
rect 30205 19397 30239 19431
rect 32873 19397 32907 19431
rect 35173 19397 35207 19431
rect 35265 19397 35299 19431
rect 8033 19329 8067 19363
rect 8401 19329 8435 19363
rect 9413 19329 9447 19363
rect 9680 19329 9714 19363
rect 11713 19329 11747 19363
rect 11989 19329 12023 19363
rect 15669 19329 15703 19363
rect 15761 19329 15795 19363
rect 17601 19329 17635 19363
rect 17785 19329 17819 19363
rect 18521 19329 18555 19363
rect 18613 19329 18647 19363
rect 18889 19329 18923 19363
rect 20545 19329 20579 19363
rect 22109 19329 22143 19363
rect 22569 19329 22603 19363
rect 22661 19329 22695 19363
rect 22937 19329 22971 19363
rect 23213 19329 23247 19363
rect 23397 19329 23431 19363
rect 24409 19329 24443 19363
rect 26065 19329 26099 19363
rect 26341 19329 26375 19363
rect 26433 19329 26467 19363
rect 27169 19329 27203 19363
rect 27629 19329 27663 19363
rect 27905 19329 27939 19363
rect 28733 19329 28767 19363
rect 28826 19329 28860 19363
rect 29239 19329 29273 19363
rect 29844 19329 29878 19363
rect 29930 19329 29964 19363
rect 30113 19329 30147 19363
rect 30302 19329 30336 19363
rect 33057 19329 33091 19363
rect 33149 19329 33183 19363
rect 34897 19329 34931 19363
rect 35045 19329 35079 19363
rect 35403 19329 35437 19363
rect 37841 19329 37875 19363
rect 38117 19329 38151 19363
rect 5549 19261 5583 19295
rect 5733 19261 5767 19295
rect 15945 19261 15979 19295
rect 17877 19261 17911 19295
rect 19901 19261 19935 19295
rect 24685 19261 24719 19295
rect 10793 19193 10827 19227
rect 24961 19193 24995 19227
rect 5089 19125 5123 19159
rect 8585 19125 8619 19159
rect 18337 19125 18371 19159
rect 18797 19125 18831 19159
rect 24501 19125 24535 19159
rect 26617 19125 26651 19159
rect 29377 19125 29411 19159
rect 30481 19125 30515 19159
rect 32873 19125 32907 19159
rect 9965 18921 9999 18955
rect 13277 18921 13311 18955
rect 15393 18921 15427 18955
rect 17969 18921 18003 18955
rect 21557 18921 21591 18955
rect 23489 18921 23523 18955
rect 24593 18921 24627 18955
rect 24961 18921 24995 18955
rect 33425 18921 33459 18955
rect 5641 18853 5675 18887
rect 32229 18853 32263 18887
rect 4261 18785 4295 18819
rect 8125 18785 8159 18819
rect 13093 18785 13127 18819
rect 16957 18785 16991 18819
rect 18337 18785 18371 18819
rect 18429 18785 18463 18819
rect 20361 18785 20395 18819
rect 21649 18785 21683 18819
rect 23949 18785 23983 18819
rect 25881 18785 25915 18819
rect 6469 18717 6503 18751
rect 6561 18717 6595 18751
rect 9413 18717 9447 18751
rect 9781 18717 9815 18751
rect 13277 18717 13311 18751
rect 14289 18717 14323 18751
rect 15301 18717 15335 18751
rect 17141 18717 17175 18751
rect 17233 18717 17267 18751
rect 17417 18717 17451 18751
rect 17509 18717 17543 18751
rect 18153 18717 18187 18751
rect 21833 18717 21867 18751
rect 22477 18717 22511 18751
rect 22661 18717 22695 18751
rect 23673 18717 23707 18751
rect 23857 18717 23891 18751
rect 24593 18717 24627 18751
rect 24685 18717 24719 18751
rect 30849 18717 30883 18751
rect 31309 18717 31343 18751
rect 31769 18717 31803 18751
rect 32045 18717 32079 18751
rect 32781 18717 32815 18751
rect 32929 18717 32963 18751
rect 33246 18717 33280 18751
rect 35070 18717 35104 18751
rect 35174 18717 35208 18751
rect 35357 18717 35391 18751
rect 35449 18717 35483 18751
rect 35546 18717 35580 18751
rect 36737 18717 36771 18751
rect 4528 18649 4562 18683
rect 6837 18649 6871 18683
rect 6929 18649 6963 18683
rect 7389 18649 7423 18683
rect 9597 18649 9631 18683
rect 9689 18649 9723 18683
rect 13001 18649 13035 18683
rect 21557 18649 21591 18683
rect 26148 18649 26182 18683
rect 33057 18649 33091 18683
rect 33149 18649 33183 18683
rect 37004 18649 37038 18683
rect 6285 18581 6319 18615
rect 13461 18581 13495 18615
rect 14381 18581 14415 18615
rect 19809 18581 19843 18615
rect 20177 18581 20211 18615
rect 20269 18581 20303 18615
rect 22017 18581 22051 18615
rect 22569 18581 22603 18615
rect 27261 18581 27295 18615
rect 35725 18581 35759 18615
rect 38117 18581 38151 18615
rect 6929 18377 6963 18411
rect 9321 18377 9355 18411
rect 13093 18377 13127 18411
rect 13185 18377 13219 18411
rect 13921 18377 13955 18411
rect 14289 18377 14323 18411
rect 14381 18377 14415 18411
rect 18521 18377 18555 18411
rect 18613 18377 18647 18411
rect 19349 18377 19383 18411
rect 19809 18377 19843 18411
rect 24317 18377 24351 18411
rect 30757 18377 30791 18411
rect 33701 18377 33735 18411
rect 37473 18377 37507 18411
rect 37841 18377 37875 18411
rect 8208 18309 8242 18343
rect 10333 18309 10367 18343
rect 19717 18309 19751 18343
rect 24777 18309 24811 18343
rect 29377 18309 29411 18343
rect 35541 18309 35575 18343
rect 37933 18309 37967 18343
rect 6837 18241 6871 18275
rect 7021 18241 7055 18275
rect 10057 18241 10091 18275
rect 10241 18241 10275 18275
rect 10425 18241 10459 18275
rect 15301 18241 15335 18275
rect 15485 18241 15519 18275
rect 15577 18241 15611 18275
rect 17141 18241 17175 18275
rect 17417 18241 17451 18275
rect 17601 18241 17635 18275
rect 22017 18241 22051 18275
rect 22293 18241 22327 18275
rect 23029 18241 23063 18275
rect 23213 18241 23247 18275
rect 24041 18241 24075 18275
rect 28365 18241 28399 18275
rect 29193 18241 29227 18275
rect 30573 18241 30607 18275
rect 30757 18241 30791 18275
rect 33333 18241 33367 18275
rect 33517 18241 33551 18275
rect 35725 18241 35759 18275
rect 35817 18241 35851 18275
rect 36093 18241 36127 18275
rect 7941 18173 7975 18207
rect 13277 18173 13311 18207
rect 14565 18173 14599 18207
rect 17233 18173 17267 18207
rect 18705 18173 18739 18207
rect 19901 18173 19935 18207
rect 22109 18173 22143 18207
rect 23673 18173 23707 18207
rect 24133 18173 24167 18207
rect 25605 18173 25639 18207
rect 28273 18173 28307 18207
rect 28733 18173 28767 18207
rect 31125 18173 31159 18207
rect 38025 18173 38059 18207
rect 36001 18105 36035 18139
rect 10609 18037 10643 18071
rect 12725 18037 12759 18071
rect 15117 18037 15151 18071
rect 16865 18037 16899 18071
rect 17325 18037 17359 18071
rect 18153 18037 18187 18071
rect 22293 18037 22327 18071
rect 22477 18037 22511 18071
rect 23121 18037 23155 18071
rect 29561 18037 29595 18071
rect 11437 17833 11471 17867
rect 30297 17833 30331 17867
rect 31401 17833 31435 17867
rect 33517 17833 33551 17867
rect 21833 17765 21867 17799
rect 22937 17765 22971 17799
rect 5825 17697 5859 17731
rect 10057 17697 10091 17731
rect 12817 17697 12851 17731
rect 13001 17697 13035 17731
rect 16773 17697 16807 17731
rect 24685 17697 24719 17731
rect 38117 17697 38151 17731
rect 6092 17629 6126 17663
rect 10324 17629 10358 17663
rect 14657 17629 14691 17663
rect 14750 17629 14784 17663
rect 15025 17629 15059 17663
rect 15122 17629 15156 17663
rect 19533 17629 19567 17663
rect 19625 17629 19659 17663
rect 21281 17629 21315 17663
rect 21557 17629 21591 17663
rect 21701 17629 21735 17663
rect 22937 17629 22971 17663
rect 23213 17629 23247 17663
rect 23673 17629 23707 17663
rect 24777 17629 24811 17663
rect 25237 17629 25271 17663
rect 25329 17629 25363 17663
rect 27077 17629 27111 17663
rect 27170 17629 27204 17663
rect 27542 17629 27576 17663
rect 29870 17629 29904 17663
rect 30389 17629 30423 17663
rect 30849 17629 30883 17663
rect 31217 17629 31251 17663
rect 31861 17629 31895 17663
rect 32045 17629 32079 17663
rect 32229 17629 32263 17663
rect 33149 17629 33183 17663
rect 33517 17629 33551 17663
rect 37841 17629 37875 17663
rect 14933 17561 14967 17595
rect 16589 17561 16623 17595
rect 21465 17561 21499 17595
rect 23857 17561 23891 17595
rect 27353 17561 27387 17595
rect 27445 17561 27479 17595
rect 31033 17561 31067 17595
rect 31125 17561 31159 17595
rect 32137 17561 32171 17595
rect 7205 17493 7239 17527
rect 12357 17493 12391 17527
rect 12725 17493 12759 17527
rect 15301 17493 15335 17527
rect 16129 17493 16163 17527
rect 16497 17493 16531 17527
rect 19809 17493 19843 17527
rect 23121 17493 23155 17527
rect 24041 17493 24075 17527
rect 25789 17493 25823 17527
rect 27721 17493 27755 17527
rect 29745 17493 29779 17527
rect 29929 17493 29963 17527
rect 32413 17493 32447 17527
rect 33333 17493 33367 17527
rect 14841 17289 14875 17323
rect 15485 17289 15519 17323
rect 19625 17289 19659 17323
rect 23673 17289 23707 17323
rect 24317 17289 24351 17323
rect 26617 17289 26651 17323
rect 8309 17221 8343 17255
rect 8401 17221 8435 17255
rect 11980 17221 12014 17255
rect 18490 17221 18524 17255
rect 22569 17221 22603 17255
rect 22785 17221 22819 17255
rect 26249 17221 26283 17255
rect 27353 17221 27387 17255
rect 28457 17221 28491 17255
rect 30113 17221 30147 17255
rect 35449 17221 35483 17255
rect 36185 17221 36219 17255
rect 37933 17221 37967 17255
rect 8125 17153 8159 17187
rect 8493 17153 8527 17187
rect 14749 17153 14783 17187
rect 14933 17153 14967 17187
rect 15669 17153 15703 17187
rect 15853 17153 15887 17187
rect 15945 17153 15979 17187
rect 18245 17153 18279 17187
rect 23397 17153 23431 17187
rect 23581 17153 23615 17187
rect 24501 17153 24535 17187
rect 24593 17153 24627 17187
rect 26065 17153 26099 17187
rect 26341 17153 26375 17187
rect 26433 17153 26467 17187
rect 27169 17153 27203 17187
rect 27445 17153 27479 17187
rect 27537 17153 27571 17187
rect 28181 17153 28215 17187
rect 28365 17153 28399 17187
rect 28549 17153 28583 17187
rect 29837 17153 29871 17187
rect 30021 17153 30055 17187
rect 30205 17153 30239 17187
rect 32965 17153 32999 17187
rect 33425 17153 33459 17187
rect 35081 17153 35115 17187
rect 35174 17153 35208 17187
rect 35357 17153 35391 17187
rect 35546 17153 35580 17187
rect 36369 17153 36403 17187
rect 36461 17153 36495 17187
rect 36737 17153 36771 17187
rect 37841 17153 37875 17187
rect 11713 17085 11747 17119
rect 24685 17085 24719 17119
rect 24777 17085 24811 17119
rect 32873 17085 32907 17119
rect 36645 17085 36679 17119
rect 38025 17085 38059 17119
rect 13093 17017 13127 17051
rect 22937 17017 22971 17051
rect 33793 17017 33827 17051
rect 35725 17017 35759 17051
rect 8677 16949 8711 16983
rect 22713 16949 22747 16983
rect 27721 16949 27755 16983
rect 28733 16949 28767 16983
rect 30389 16949 30423 16983
rect 37473 16949 37507 16983
rect 8033 16745 8067 16779
rect 10517 16745 10551 16779
rect 22845 16745 22879 16779
rect 32505 16745 32539 16779
rect 38209 16745 38243 16779
rect 15669 16677 15703 16711
rect 17601 16677 17635 16711
rect 9137 16609 9171 16643
rect 13369 16609 13403 16643
rect 16221 16609 16255 16643
rect 19993 16609 20027 16643
rect 29101 16609 29135 16643
rect 33609 16609 33643 16643
rect 34069 16609 34103 16643
rect 36829 16609 36863 16643
rect 5641 16541 5675 16575
rect 8033 16541 8067 16575
rect 8217 16541 8251 16575
rect 9393 16541 9427 16575
rect 11529 16541 11563 16575
rect 11897 16541 11931 16575
rect 12541 16541 12575 16575
rect 15393 16541 15427 16575
rect 15485 16541 15519 16575
rect 16477 16541 16511 16575
rect 20249 16541 20283 16575
rect 22477 16541 22511 16575
rect 22937 16541 22971 16575
rect 26525 16541 26559 16575
rect 26709 16541 26743 16575
rect 26893 16541 26927 16575
rect 28825 16541 28859 16575
rect 28917 16541 28951 16575
rect 29193 16541 29227 16575
rect 31033 16541 31067 16575
rect 31125 16541 31159 16575
rect 31309 16541 31343 16575
rect 31401 16541 31435 16575
rect 31861 16541 31895 16575
rect 31954 16541 31988 16575
rect 32229 16541 32263 16575
rect 32367 16541 32401 16575
rect 33701 16541 33735 16575
rect 35081 16541 35115 16575
rect 35174 16541 35208 16575
rect 35357 16541 35391 16575
rect 35546 16541 35580 16575
rect 37096 16541 37130 16575
rect 5908 16473 5942 16507
rect 11713 16473 11747 16507
rect 11805 16473 11839 16507
rect 26801 16473 26835 16507
rect 32137 16473 32171 16507
rect 35449 16473 35483 16507
rect 7021 16405 7055 16439
rect 12081 16405 12115 16439
rect 21373 16405 21407 16439
rect 27077 16405 27111 16439
rect 28641 16405 28675 16439
rect 30849 16405 30883 16439
rect 35725 16405 35759 16439
rect 6561 16201 6595 16235
rect 7941 16201 7975 16235
rect 13553 16201 13587 16235
rect 18889 16201 18923 16235
rect 25329 16201 25363 16235
rect 30481 16201 30515 16235
rect 37841 16201 37875 16235
rect 6929 16133 6963 16167
rect 12418 16133 12452 16167
rect 15853 16133 15887 16167
rect 22753 16133 22787 16167
rect 22969 16133 23003 16167
rect 31033 16133 31067 16167
rect 31125 16133 31159 16167
rect 32597 16133 32631 16167
rect 7938 16065 7972 16099
rect 14197 16065 14231 16099
rect 17601 16065 17635 16099
rect 17785 16065 17819 16099
rect 17877 16065 17911 16099
rect 19073 16065 19107 16099
rect 19257 16065 19291 16099
rect 19625 16065 19659 16099
rect 25145 16065 25179 16099
rect 27445 16065 27479 16099
rect 27629 16065 27663 16099
rect 27757 16065 27791 16099
rect 29193 16065 29227 16099
rect 29285 16065 29319 16099
rect 29469 16065 29503 16099
rect 30665 16065 30699 16099
rect 30758 16066 30792 16100
rect 32321 16065 32355 16099
rect 32505 16065 32539 16099
rect 32689 16065 32723 16099
rect 35725 16065 35759 16099
rect 35817 16065 35851 16099
rect 36093 16065 36127 16099
rect 7021 15997 7055 16031
rect 7205 15997 7239 16031
rect 8401 15997 8435 16031
rect 12173 15997 12207 16031
rect 14473 15997 14507 16031
rect 25421 15997 25455 16031
rect 27541 15997 27575 16031
rect 29377 15997 29411 16031
rect 35541 15997 35575 16031
rect 37933 15997 37967 16031
rect 38025 15997 38059 16031
rect 23121 15929 23155 15963
rect 32873 15929 32907 15963
rect 36001 15929 36035 15963
rect 7757 15861 7791 15895
rect 8309 15861 8343 15895
rect 17417 15861 17451 15895
rect 22937 15861 22971 15895
rect 24869 15861 24903 15895
rect 27261 15861 27295 15895
rect 29009 15861 29043 15895
rect 37473 15861 37507 15895
rect 8125 15657 8159 15691
rect 24961 15657 24995 15691
rect 27077 15657 27111 15691
rect 29837 15657 29871 15691
rect 36369 15657 36403 15691
rect 11161 15589 11195 15623
rect 20177 15589 20211 15623
rect 25881 15589 25915 15623
rect 33333 15589 33367 15623
rect 34161 15589 34195 15623
rect 6745 15521 6779 15555
rect 18429 15521 18463 15555
rect 19809 15521 19843 15555
rect 21097 15521 21131 15555
rect 24869 15521 24903 15555
rect 31585 15521 31619 15555
rect 31677 15521 31711 15555
rect 33885 15521 33919 15555
rect 38117 15521 38151 15555
rect 7012 15453 7046 15487
rect 9781 15453 9815 15487
rect 15393 15453 15427 15487
rect 15761 15453 15795 15487
rect 16037 15453 16071 15487
rect 17601 15453 17635 15487
rect 18153 15453 18187 15487
rect 21281 15453 21315 15487
rect 21557 15453 21591 15487
rect 21925 15453 21959 15487
rect 22201 15453 22235 15487
rect 23121 15453 23155 15487
rect 23305 15453 23339 15487
rect 23489 15453 23523 15487
rect 24777 15453 24811 15487
rect 25881 15453 25915 15487
rect 26065 15453 26099 15487
rect 26157 15453 26191 15487
rect 26985 15453 27019 15487
rect 27169 15453 27203 15487
rect 28089 15453 28123 15487
rect 28273 15453 28307 15487
rect 28549 15453 28583 15487
rect 29745 15453 29779 15487
rect 29929 15453 29963 15487
rect 32965 15453 32999 15487
rect 34989 15453 35023 15487
rect 37841 15453 37875 15487
rect 10048 15385 10082 15419
rect 35234 15385 35268 15419
rect 15301 15317 15335 15351
rect 17693 15317 17727 15351
rect 20269 15317 20303 15351
rect 25145 15317 25179 15351
rect 28457 15317 28491 15351
rect 31125 15317 31159 15351
rect 31493 15317 31527 15351
rect 33425 15317 33459 15351
rect 34345 15317 34379 15351
rect 8861 15113 8895 15147
rect 10057 15113 10091 15147
rect 13737 15113 13771 15147
rect 18981 15113 19015 15147
rect 21097 15045 21131 15079
rect 25605 15045 25639 15079
rect 25697 15045 25731 15079
rect 31493 15045 31527 15079
rect 38117 15045 38151 15079
rect 8769 14977 8803 15011
rect 10241 14977 10275 15011
rect 10517 14977 10551 15011
rect 11805 14977 11839 15011
rect 13369 14977 13403 15011
rect 15025 14977 15059 15011
rect 15209 14977 15243 15011
rect 15945 14977 15979 15011
rect 16313 14977 16347 15011
rect 17095 14977 17129 15011
rect 17233 14977 17267 15011
rect 17346 14980 17380 15014
rect 17509 14977 17543 15011
rect 19211 14977 19245 15011
rect 19349 14977 19383 15011
rect 19441 14977 19475 15011
rect 19625 14977 19659 15011
rect 20821 14977 20855 15011
rect 21005 14977 21039 15011
rect 21241 14977 21275 15011
rect 22017 14977 22051 15011
rect 22201 14977 22235 15011
rect 22293 14977 22327 15011
rect 22437 14977 22471 15011
rect 22586 14977 22620 15011
rect 24225 14977 24259 15011
rect 24501 14977 24535 15011
rect 25421 14977 25455 15011
rect 25794 14977 25828 15011
rect 27813 14977 27847 15011
rect 28181 14977 28215 15011
rect 31217 14977 31251 15011
rect 33517 14977 33551 15011
rect 33701 14977 33735 15011
rect 37841 14977 37875 15011
rect 9045 14909 9079 14943
rect 10425 14909 10459 14943
rect 11713 14909 11747 14943
rect 12265 14909 12299 14943
rect 13461 14909 13495 14943
rect 17969 14909 18003 14943
rect 27629 14909 27663 14943
rect 15393 14841 15427 14875
rect 18337 14841 18371 14875
rect 28089 14841 28123 14875
rect 8401 14773 8435 14807
rect 16865 14773 16899 14807
rect 18429 14773 18463 14807
rect 21373 14773 21407 14807
rect 24041 14773 24075 14807
rect 24409 14773 24443 14807
rect 25973 14773 26007 14807
rect 33517 14773 33551 14807
rect 13461 14569 13495 14603
rect 17141 14569 17175 14603
rect 19533 14569 19567 14603
rect 25421 14569 25455 14603
rect 27813 14569 27847 14603
rect 34897 14569 34931 14603
rect 38301 14569 38335 14603
rect 22017 14501 22051 14535
rect 29193 14501 29227 14535
rect 8401 14433 8435 14467
rect 17785 14433 17819 14467
rect 20177 14433 20211 14467
rect 24041 14433 24075 14467
rect 28733 14433 28767 14467
rect 29837 14433 29871 14467
rect 33333 14433 33367 14467
rect 35081 14433 35115 14467
rect 35449 14433 35483 14467
rect 7665 14365 7699 14399
rect 11897 14365 11931 14399
rect 12081 14365 12115 14399
rect 12265 14365 12299 14399
rect 13369 14365 13403 14399
rect 13553 14365 13587 14399
rect 15209 14365 15243 14399
rect 17509 14365 17543 14399
rect 18705 14365 18739 14399
rect 18889 14365 18923 14399
rect 21465 14365 21499 14399
rect 21649 14365 21683 14399
rect 21885 14365 21919 14399
rect 23561 14365 23595 14399
rect 23673 14365 23707 14399
rect 24593 14365 24627 14399
rect 24777 14365 24811 14399
rect 25421 14365 25455 14399
rect 25605 14365 25639 14399
rect 27721 14365 27755 14399
rect 28825 14365 28859 14399
rect 29929 14365 29963 14399
rect 33241 14365 33275 14399
rect 35174 14365 35208 14399
rect 36921 14365 36955 14399
rect 37188 14365 37222 14399
rect 15485 14297 15519 14331
rect 17601 14297 17635 14331
rect 21741 14297 21775 14331
rect 23949 14297 23983 14331
rect 35541 14297 35575 14331
rect 18797 14229 18831 14263
rect 19901 14229 19935 14263
rect 19993 14229 20027 14263
rect 23397 14229 23431 14263
rect 24961 14229 24995 14263
rect 30297 14229 30331 14263
rect 33609 14229 33643 14263
rect 9321 14025 9355 14059
rect 17509 14025 17543 14059
rect 19901 14025 19935 14059
rect 22753 14025 22787 14059
rect 24409 14025 24443 14059
rect 31769 14025 31803 14059
rect 32781 14025 32815 14059
rect 35265 14025 35299 14059
rect 8208 13957 8242 13991
rect 16865 13957 16899 13991
rect 19257 13957 19291 13991
rect 23765 13957 23799 13991
rect 24961 13957 24995 13991
rect 27169 13957 27203 13991
rect 27353 13957 27387 13991
rect 33425 13957 33459 13991
rect 36461 13957 36495 13991
rect 7941 13889 7975 13923
rect 10609 13889 10643 13923
rect 11713 13889 11747 13923
rect 11897 13889 11931 13923
rect 12909 13889 12943 13923
rect 13001 13889 13035 13923
rect 13369 13889 13403 13923
rect 14381 13889 14415 13923
rect 14841 13889 14875 13923
rect 15393 13889 15427 13923
rect 17233 13889 17267 13923
rect 19625 13889 19659 13923
rect 19717 13889 19751 13923
rect 22937 13889 22971 13923
rect 23213 13889 23247 13923
rect 24225 13889 24259 13923
rect 24869 13889 24903 13923
rect 25053 13889 25087 13923
rect 26065 13889 26099 13923
rect 26341 13889 26375 13923
rect 27445 13889 27479 13923
rect 27997 13889 28031 13923
rect 28825 13889 28859 13923
rect 30656 13889 30690 13923
rect 33057 13889 33091 13923
rect 33885 13889 33919 13923
rect 34141 13889 34175 13923
rect 36093 13889 36127 13923
rect 36369 13889 36403 13923
rect 10701 13821 10735 13855
rect 12081 13821 12115 13855
rect 13093 13821 13127 13855
rect 15209 13821 15243 13855
rect 17325 13821 17359 13855
rect 23029 13821 23063 13855
rect 23121 13821 23155 13855
rect 24133 13821 24167 13855
rect 25513 13821 25547 13855
rect 26525 13821 26559 13855
rect 30389 13821 30423 13855
rect 32965 13821 32999 13855
rect 33333 13821 33367 13855
rect 36001 13821 36035 13855
rect 38301 13821 38335 13855
rect 10977 13753 11011 13787
rect 13829 13753 13863 13787
rect 15025 13753 15059 13787
rect 35817 13753 35851 13787
rect 27169 13685 27203 13719
rect 28181 13685 28215 13719
rect 29285 13685 29319 13719
rect 10701 13481 10735 13515
rect 15853 13481 15887 13515
rect 23581 13481 23615 13515
rect 37105 13481 37139 13515
rect 25881 13413 25915 13447
rect 27169 13413 27203 13447
rect 10517 13345 10551 13379
rect 14289 13345 14323 13379
rect 21833 13345 21867 13379
rect 26985 13345 27019 13379
rect 28457 13345 28491 13379
rect 30849 13345 30883 13379
rect 35725 13345 35759 13379
rect 10425 13277 10459 13311
rect 12173 13277 12207 13311
rect 14473 13277 14507 13311
rect 14841 13277 14875 13311
rect 16221 13277 16255 13311
rect 16497 13277 16531 13311
rect 16589 13277 16623 13311
rect 16865 13277 16899 13311
rect 17141 13277 17175 13311
rect 17693 13277 17727 13311
rect 17877 13277 17911 13311
rect 17969 13277 18003 13311
rect 18153 13277 18187 13311
rect 18245 13277 18279 13311
rect 20913 13277 20947 13311
rect 21097 13277 21131 13311
rect 21557 13277 21591 13311
rect 21649 13277 21683 13311
rect 23581 13277 23615 13311
rect 23857 13277 23891 13311
rect 25881 13277 25915 13311
rect 26157 13277 26191 13311
rect 27261 13277 27295 13311
rect 28365 13277 28399 13311
rect 28733 13277 28767 13311
rect 28825 13277 28859 13311
rect 30941 13277 30975 13311
rect 31125 13277 31159 13311
rect 35981 13277 36015 13311
rect 12909 13209 12943 13243
rect 23765 13209 23799 13243
rect 26065 13209 26099 13243
rect 27721 13209 27755 13243
rect 31585 13209 31619 13243
rect 14473 13141 14507 13175
rect 21097 13141 21131 13175
rect 21833 13141 21867 13175
rect 26801 13141 26835 13175
rect 13737 12937 13771 12971
rect 14381 12937 14415 12971
rect 15945 12937 15979 12971
rect 17785 12937 17819 12971
rect 33057 12937 33091 12971
rect 11161 12869 11195 12903
rect 13277 12869 13311 12903
rect 22017 12869 22051 12903
rect 29285 12869 29319 12903
rect 7665 12801 7699 12835
rect 7932 12801 7966 12835
rect 9505 12801 9539 12835
rect 12541 12801 12575 12835
rect 12725 12801 12759 12835
rect 12817 12801 12851 12835
rect 14378 12801 14412 12835
rect 15669 12801 15703 12835
rect 15761 12801 15795 12835
rect 17417 12801 17451 12835
rect 17601 12801 17635 12835
rect 19533 12801 19567 12835
rect 19717 12801 19751 12835
rect 19809 12801 19843 12835
rect 21097 12801 21131 12835
rect 21189 12801 21223 12835
rect 21465 12801 21499 12835
rect 22201 12801 22235 12835
rect 22385 12801 22419 12835
rect 25421 12801 25455 12835
rect 25605 12801 25639 12835
rect 25789 12801 25823 12835
rect 25881 12801 25915 12835
rect 28273 12801 28307 12835
rect 28733 12801 28767 12835
rect 28917 12801 28951 12835
rect 32965 12801 32999 12835
rect 9781 12733 9815 12767
rect 14841 12733 14875 12767
rect 15945 12733 15979 12767
rect 22477 12733 22511 12767
rect 27997 12733 28031 12767
rect 33149 12733 33183 12767
rect 13645 12665 13679 12699
rect 28181 12665 28215 12699
rect 29193 12665 29227 12699
rect 9045 12597 9079 12631
rect 12541 12597 12575 12631
rect 14197 12597 14231 12631
rect 14749 12597 14783 12631
rect 19349 12597 19383 12631
rect 20913 12597 20947 12631
rect 21373 12597 21407 12631
rect 27813 12597 27847 12631
rect 32597 12597 32631 12631
rect 38301 12597 38335 12631
rect 9689 12393 9723 12427
rect 13185 12393 13219 12427
rect 15025 12393 15059 12427
rect 16957 12393 16991 12427
rect 21005 12393 21039 12427
rect 25421 12393 25455 12427
rect 28273 12393 28307 12427
rect 29009 12393 29043 12427
rect 33885 12393 33919 12427
rect 12357 12325 12391 12359
rect 16313 12325 16347 12359
rect 24593 12325 24627 12359
rect 9229 12257 9263 12291
rect 12449 12257 12483 12291
rect 15577 12257 15611 12291
rect 16497 12257 16531 12291
rect 17141 12257 17175 12291
rect 17233 12257 17267 12291
rect 18685 12257 18719 12291
rect 19901 12257 19935 12291
rect 22017 12257 22051 12291
rect 25789 12257 25823 12291
rect 25973 12257 26007 12291
rect 31677 12257 31711 12291
rect 35541 12257 35575 12291
rect 36829 12257 36863 12291
rect 9321 12189 9355 12223
rect 12173 12189 12207 12223
rect 12265 12189 12299 12223
rect 13185 12189 13219 12223
rect 13369 12189 13403 12223
rect 16221 12189 16255 12223
rect 17325 12189 17359 12223
rect 17417 12189 17451 12223
rect 18797 12189 18831 12223
rect 18889 12189 18923 12223
rect 19625 12189 19659 12223
rect 19717 12189 19751 12223
rect 19993 12189 20027 12223
rect 21189 12189 21223 12223
rect 21373 12189 21407 12223
rect 21465 12189 21499 12223
rect 21925 12189 21959 12223
rect 22109 12189 22143 12223
rect 24869 12189 24903 12223
rect 28273 12189 28307 12223
rect 28549 12189 28583 12223
rect 29009 12189 29043 12223
rect 29193 12189 29227 12223
rect 32505 12189 32539 12223
rect 32761 12189 32795 12223
rect 15301 12121 15335 12155
rect 16497 12121 16531 12155
rect 18613 12121 18647 12155
rect 24593 12121 24627 12155
rect 31585 12121 31619 12155
rect 35357 12121 35391 12155
rect 37096 12121 37130 12155
rect 15485 12053 15519 12087
rect 19441 12053 19475 12087
rect 24777 12053 24811 12087
rect 25881 12053 25915 12087
rect 28457 12053 28491 12087
rect 31125 12053 31159 12087
rect 31493 12053 31527 12087
rect 34989 12053 35023 12087
rect 35449 12053 35483 12087
rect 38209 12053 38243 12087
rect 9321 11849 9355 11883
rect 10425 11849 10459 11883
rect 14749 11849 14783 11883
rect 15117 11849 15151 11883
rect 19073 11849 19107 11883
rect 19625 11849 19659 11883
rect 24777 11849 24811 11883
rect 25237 11849 25271 11883
rect 26341 11849 26375 11883
rect 35173 11849 35207 11883
rect 37473 11849 37507 11883
rect 37841 11849 37875 11883
rect 8208 11781 8242 11815
rect 12357 11781 12391 11815
rect 12541 11781 12575 11815
rect 17509 11781 17543 11815
rect 25973 11781 26007 11815
rect 26173 11781 26207 11815
rect 30656 11781 30690 11815
rect 10609 11713 10643 11747
rect 10793 11713 10827 11747
rect 10885 11713 10919 11747
rect 15209 11713 15243 11747
rect 17693 11713 17727 11747
rect 18981 11713 19015 11747
rect 19165 11713 19199 11747
rect 19809 11713 19843 11747
rect 19993 11713 20027 11747
rect 20085 11713 20119 11747
rect 22937 11713 22971 11747
rect 23204 11713 23238 11747
rect 25145 11713 25179 11747
rect 29285 11713 29319 11747
rect 30389 11713 30423 11747
rect 32321 11713 32355 11747
rect 32873 11713 32907 11747
rect 33149 11713 33183 11747
rect 33793 11713 33827 11747
rect 35081 11713 35115 11747
rect 35909 11713 35943 11747
rect 36553 11713 36587 11747
rect 7941 11645 7975 11679
rect 15393 11645 15427 11679
rect 25421 11645 25455 11679
rect 29377 11645 29411 11679
rect 29469 11645 29503 11679
rect 33057 11645 33091 11679
rect 33517 11645 33551 11679
rect 35817 11645 35851 11679
rect 36277 11645 36311 11679
rect 37933 11645 37967 11679
rect 38117 11645 38151 11679
rect 17877 11577 17911 11611
rect 24317 11577 24351 11611
rect 31769 11577 31803 11611
rect 12725 11509 12759 11543
rect 26157 11509 26191 11543
rect 28917 11509 28951 11543
rect 10977 11305 11011 11339
rect 12265 11305 12299 11339
rect 15025 11305 15059 11339
rect 19717 11305 19751 11339
rect 21649 11305 21683 11339
rect 36277 11305 36311 11339
rect 18061 11237 18095 11271
rect 29837 11237 29871 11271
rect 10149 11169 10183 11203
rect 25421 11169 25455 11203
rect 25605 11169 25639 11203
rect 30481 11169 30515 11203
rect 33885 11169 33919 11203
rect 34897 11169 34931 11203
rect 10057 11101 10091 11135
rect 10333 11101 10367 11135
rect 10425 11101 10459 11135
rect 11161 11101 11195 11135
rect 11253 11101 11287 11135
rect 11437 11101 11471 11135
rect 11529 11101 11563 11135
rect 12265 11101 12299 11135
rect 12541 11101 12575 11135
rect 15025 11101 15059 11135
rect 15301 11101 15335 11135
rect 16497 11101 16531 11135
rect 16681 11101 16715 11135
rect 17141 11101 17175 11135
rect 19625 11101 19659 11135
rect 19809 11101 19843 11135
rect 21557 11101 21591 11135
rect 21833 11101 21867 11135
rect 26709 11101 26743 11135
rect 29745 11101 29779 11135
rect 30573 11101 30607 11135
rect 31033 11101 31067 11135
rect 31401 11101 31435 11135
rect 36737 11101 36771 11135
rect 15209 11033 15243 11067
rect 16589 11033 16623 11067
rect 17785 11033 17819 11067
rect 25329 11033 25363 11067
rect 26976 11033 27010 11067
rect 33149 11033 33183 11067
rect 35142 11033 35176 11067
rect 37004 11033 37038 11067
rect 10517 10965 10551 10999
rect 12449 10965 12483 10999
rect 17233 10965 17267 10999
rect 18245 10965 18279 10999
rect 22109 10965 22143 10999
rect 24961 10965 24995 10999
rect 28089 10965 28123 10999
rect 38117 10965 38151 10999
rect 17785 10761 17819 10795
rect 18521 10761 18555 10795
rect 21097 10761 21131 10795
rect 25973 10761 26007 10795
rect 27169 10761 27203 10795
rect 27537 10761 27571 10795
rect 30113 10761 30147 10795
rect 37473 10761 37507 10795
rect 17693 10693 17727 10727
rect 22293 10693 22327 10727
rect 29000 10693 29034 10727
rect 37933 10693 37967 10727
rect 11805 10625 11839 10659
rect 11989 10625 12023 10659
rect 13185 10625 13219 10659
rect 13369 10625 13403 10659
rect 15393 10625 15427 10659
rect 15577 10625 15611 10659
rect 18889 10625 18923 10659
rect 22017 10625 22051 10659
rect 22201 10625 22235 10659
rect 22385 10625 22419 10659
rect 24860 10625 24894 10659
rect 27629 10625 27663 10659
rect 28733 10625 28767 10659
rect 34253 10625 34287 10659
rect 37841 10625 37875 10659
rect 17877 10557 17911 10591
rect 18981 10557 19015 10591
rect 21189 10557 21223 10591
rect 21281 10557 21315 10591
rect 24593 10557 24627 10591
rect 27721 10557 27755 10591
rect 34345 10557 34379 10591
rect 34437 10557 34471 10591
rect 38117 10557 38151 10591
rect 22569 10489 22603 10523
rect 11897 10421 11931 10455
rect 13553 10421 13587 10455
rect 15393 10421 15427 10455
rect 17325 10421 17359 10455
rect 19165 10421 19199 10455
rect 20729 10421 20763 10455
rect 33885 10421 33919 10455
rect 10701 10217 10735 10251
rect 13185 10217 13219 10251
rect 21925 10217 21959 10251
rect 24869 10217 24903 10251
rect 24961 10217 24995 10251
rect 31861 10217 31895 10251
rect 17233 10149 17267 10183
rect 21833 10149 21867 10183
rect 22569 10149 22603 10183
rect 34345 10149 34379 10183
rect 35081 10149 35115 10183
rect 9137 10081 9171 10115
rect 13277 10081 13311 10115
rect 15669 10081 15703 10115
rect 22017 10081 22051 10115
rect 25053 10081 25087 10115
rect 26893 10081 26927 10115
rect 32965 10081 32999 10115
rect 35725 10081 35759 10115
rect 36185 10081 36219 10115
rect 38117 10081 38151 10115
rect 9413 10013 9447 10047
rect 11253 10013 11287 10047
rect 11529 10013 11563 10047
rect 13185 10013 13219 10047
rect 15393 10013 15427 10047
rect 16405 10013 16439 10047
rect 16773 10013 16807 10047
rect 17417 10013 17451 10047
rect 18705 10013 18739 10047
rect 18889 10013 18923 10047
rect 21741 10013 21775 10047
rect 22477 10013 22511 10047
rect 22661 10013 22695 10047
rect 24777 10013 24811 10047
rect 32137 10013 32171 10047
rect 32229 10013 32263 10047
rect 32321 10013 32355 10047
rect 32505 10013 32539 10047
rect 33232 10013 33266 10047
rect 34989 10013 35023 10047
rect 35909 10013 35943 10047
rect 36461 10013 36495 10047
rect 37841 10013 37875 10047
rect 11437 9945 11471 9979
rect 16221 9945 16255 9979
rect 17785 9945 17819 9979
rect 18797 9945 18831 9979
rect 26157 9945 26191 9979
rect 11345 9877 11379 9911
rect 13553 9877 13587 9911
rect 15025 9877 15059 9911
rect 15485 9877 15519 9911
rect 17509 9877 17543 9911
rect 17601 9877 17635 9911
rect 15485 9673 15519 9707
rect 24133 9673 24167 9707
rect 33609 9673 33643 9707
rect 11069 9605 11103 9639
rect 14657 9605 14691 9639
rect 24961 9605 24995 9639
rect 25053 9605 25087 9639
rect 26341 9605 26375 9639
rect 29193 9605 29227 9639
rect 30849 9605 30883 9639
rect 32689 9605 32723 9639
rect 38117 9605 38151 9639
rect 10885 9537 10919 9571
rect 11161 9537 11195 9571
rect 11989 9537 12023 9571
rect 12081 9537 12115 9571
rect 12173 9537 12207 9571
rect 13277 9537 13311 9571
rect 15577 9537 15611 9571
rect 18337 9537 18371 9571
rect 19165 9537 19199 9571
rect 19533 9537 19567 9571
rect 21097 9537 21131 9571
rect 21189 9537 21223 9571
rect 22753 9537 22787 9571
rect 23020 9537 23054 9571
rect 25881 9537 25915 9571
rect 27353 9537 27387 9571
rect 27620 9537 27654 9571
rect 29469 9537 29503 9571
rect 29561 9537 29595 9571
rect 29653 9537 29687 9571
rect 29837 9537 29871 9571
rect 30297 9537 30331 9571
rect 30389 9537 30423 9571
rect 34161 9537 34195 9571
rect 34713 9537 34747 9571
rect 37841 9537 37875 9571
rect 12449 9469 12483 9503
rect 13001 9469 13035 9503
rect 15761 9469 15795 9503
rect 21373 9469 21407 9503
rect 25237 9469 25271 9503
rect 32781 9469 32815 9503
rect 32873 9469 32907 9503
rect 10701 9401 10735 9435
rect 11713 9401 11747 9435
rect 24593 9401 24627 9435
rect 28733 9401 28767 9435
rect 12357 9333 12391 9367
rect 15117 9333 15151 9367
rect 20729 9333 20763 9367
rect 32321 9333 32355 9367
rect 10885 9129 10919 9163
rect 26249 9129 26283 9163
rect 27997 9129 28031 9163
rect 32597 9129 32631 9163
rect 33425 9129 33459 9163
rect 18521 9061 18555 9095
rect 19441 9061 19475 9095
rect 20821 9061 20855 9095
rect 35449 9061 35483 9095
rect 10517 8993 10551 9027
rect 12633 8993 12667 9027
rect 13001 8993 13035 9027
rect 13093 8993 13127 9027
rect 16957 8993 16991 9027
rect 18705 8993 18739 9027
rect 20085 8993 20119 9027
rect 21373 8993 21407 9027
rect 25513 8993 25547 9027
rect 25697 8993 25731 9027
rect 28457 8993 28491 9027
rect 28549 8993 28583 9027
rect 36093 8993 36127 9027
rect 36553 8993 36587 9027
rect 10701 8925 10735 8959
rect 14473 8925 14507 8959
rect 14657 8925 14691 8959
rect 15669 8925 15703 8959
rect 15761 8925 15795 8959
rect 16773 8925 16807 8959
rect 17509 8925 17543 8959
rect 18521 8925 18555 8959
rect 25421 8925 25455 8959
rect 26433 8925 26467 8959
rect 26709 8925 26743 8959
rect 28365 8925 28399 8959
rect 30021 8925 30055 8959
rect 30113 8925 30147 8959
rect 31217 8925 31251 8959
rect 31484 8925 31518 8959
rect 33241 8925 33275 8959
rect 35449 8925 35483 8959
rect 36185 8925 36219 8959
rect 36829 8925 36863 8959
rect 37841 8925 37875 8959
rect 14841 8857 14875 8891
rect 16681 8857 16715 8891
rect 17601 8857 17635 8891
rect 18889 8857 18923 8891
rect 21097 8857 21131 8891
rect 21281 8857 21315 8891
rect 26617 8857 26651 8891
rect 30573 8857 30607 8891
rect 33057 8857 33091 8891
rect 38117 8857 38151 8891
rect 13277 8789 13311 8823
rect 16313 8789 16347 8823
rect 19809 8789 19843 8823
rect 19901 8789 19935 8823
rect 25053 8789 25087 8823
rect 12081 8585 12115 8619
rect 16957 8585 16991 8619
rect 21373 8585 21407 8619
rect 25881 8585 25915 8619
rect 27629 8585 27663 8619
rect 31401 8585 31435 8619
rect 32965 8585 32999 8619
rect 36185 8585 36219 8619
rect 37841 8585 37875 8619
rect 18521 8517 18555 8551
rect 20177 8517 20211 8551
rect 22017 8517 22051 8551
rect 22201 8517 22235 8551
rect 24768 8517 24802 8551
rect 29837 8517 29871 8551
rect 33793 8517 33827 8551
rect 11805 8449 11839 8483
rect 11897 8449 11931 8483
rect 13921 8449 13955 8483
rect 14841 8449 14875 8483
rect 16129 8449 16163 8483
rect 16865 8449 16899 8483
rect 17049 8449 17083 8483
rect 18705 8449 18739 8483
rect 20361 8449 20395 8483
rect 21097 8449 21131 8483
rect 21281 8449 21315 8483
rect 24501 8449 24535 8483
rect 27537 8449 27571 8483
rect 29285 8449 29319 8483
rect 29377 8449 29411 8483
rect 30941 8449 30975 8483
rect 31033 8449 31067 8483
rect 32873 8449 32907 8483
rect 33977 8449 34011 8483
rect 35072 8449 35106 8483
rect 16221 8381 16255 8415
rect 20545 8381 20579 8415
rect 20637 8381 20671 8415
rect 27721 8381 27755 8415
rect 29101 8381 29135 8415
rect 33057 8381 33091 8415
rect 34805 8381 34839 8415
rect 37933 8381 37967 8415
rect 38117 8381 38151 8415
rect 22385 8313 22419 8347
rect 34161 8313 34195 8347
rect 37473 8313 37507 8347
rect 14197 8245 14231 8279
rect 18797 8245 18831 8279
rect 27169 8245 27203 8279
rect 32505 8245 32539 8279
rect 11805 8041 11839 8075
rect 12817 8041 12851 8075
rect 15577 8041 15611 8075
rect 17601 8041 17635 8075
rect 23029 8041 23063 8075
rect 27905 8041 27939 8075
rect 28733 8041 28767 8075
rect 32045 8041 32079 8075
rect 35081 8041 35115 8075
rect 38301 8041 38335 8075
rect 18521 7905 18555 7939
rect 35633 7905 35667 7939
rect 11989 7837 12023 7871
rect 12265 7837 12299 7871
rect 12725 7837 12759 7871
rect 13001 7837 13035 7871
rect 14289 7837 14323 7871
rect 14933 7837 14967 7871
rect 16405 7837 16439 7871
rect 16497 7837 16531 7871
rect 16681 7837 16715 7871
rect 16773 7837 16807 7871
rect 17417 7837 17451 7871
rect 17693 7837 17727 7871
rect 18429 7837 18463 7871
rect 18705 7837 18739 7871
rect 19533 7837 19567 7871
rect 19625 7837 19659 7871
rect 20453 7837 20487 7871
rect 20545 7837 20579 7871
rect 20729 7837 20763 7871
rect 21649 7837 21683 7871
rect 26525 7837 26559 7871
rect 26792 7837 26826 7871
rect 28549 7837 28583 7871
rect 30665 7837 30699 7871
rect 33241 7837 33275 7871
rect 36921 7837 36955 7871
rect 37188 7837 37222 7871
rect 12909 7769 12943 7803
rect 14749 7769 14783 7803
rect 21189 7769 21223 7803
rect 21894 7769 21928 7803
rect 28365 7769 28399 7803
rect 30932 7769 30966 7803
rect 33977 7769 34011 7803
rect 35449 7769 35483 7803
rect 12173 7701 12207 7735
rect 16221 7701 16255 7735
rect 17233 7701 17267 7735
rect 35541 7701 35575 7735
rect 21465 7497 21499 7531
rect 24241 7497 24275 7531
rect 33793 7497 33827 7531
rect 34529 7497 34563 7531
rect 37841 7497 37875 7531
rect 37933 7497 37967 7531
rect 13369 7429 13403 7463
rect 21097 7429 21131 7463
rect 24041 7429 24075 7463
rect 29561 7429 29595 7463
rect 11713 7361 11747 7395
rect 14381 7361 14415 7395
rect 14473 7361 14507 7395
rect 14749 7361 14783 7395
rect 14933 7361 14967 7395
rect 17233 7361 17267 7395
rect 17417 7361 17451 7395
rect 18521 7361 18555 7395
rect 19073 7361 19107 7395
rect 20269 7361 20303 7395
rect 20361 7361 20395 7395
rect 20637 7361 20671 7395
rect 21281 7361 21315 7395
rect 29653 7361 29687 7395
rect 32413 7361 32447 7395
rect 32680 7361 32714 7395
rect 34805 7361 34839 7395
rect 34897 7361 34931 7395
rect 34989 7361 35023 7395
rect 35173 7361 35207 7395
rect 11989 7293 12023 7327
rect 17509 7293 17543 7327
rect 18153 7293 18187 7327
rect 18797 7293 18831 7327
rect 20545 7293 20579 7327
rect 38025 7293 38059 7327
rect 14565 7225 14599 7259
rect 18705 7225 18739 7259
rect 17049 7157 17083 7191
rect 20085 7157 20119 7191
rect 24225 7157 24259 7191
rect 24409 7157 24443 7191
rect 29377 7157 29411 7191
rect 29837 7157 29871 7191
rect 37473 7157 37507 7191
rect 21649 6953 21683 6987
rect 23857 6953 23891 6987
rect 25145 6953 25179 6987
rect 32965 6953 32999 6987
rect 34897 6953 34931 6987
rect 38117 6953 38151 6987
rect 14289 6885 14323 6919
rect 12541 6817 12575 6851
rect 16313 6817 16347 6851
rect 17969 6817 18003 6851
rect 18521 6817 18555 6851
rect 20821 6817 20855 6851
rect 25697 6817 25731 6851
rect 27629 6817 27663 6851
rect 28181 6817 28215 6851
rect 30757 6817 30791 6851
rect 33517 6817 33551 6851
rect 36737 6817 36771 6851
rect 12265 6749 12299 6783
rect 12357 6749 12391 6783
rect 14473 6749 14507 6783
rect 14565 6749 14599 6783
rect 14749 6749 14783 6783
rect 14841 6749 14875 6783
rect 15669 6749 15703 6783
rect 16037 6749 16071 6783
rect 17417 6749 17451 6783
rect 17693 6749 17727 6783
rect 18245 6749 18279 6783
rect 19993 6749 20027 6783
rect 20545 6749 20579 6783
rect 21557 6749 21591 6783
rect 21741 6749 21775 6783
rect 22477 6749 22511 6783
rect 26249 6749 26283 6783
rect 27721 6749 27755 6783
rect 30021 6749 30055 6783
rect 30113 6749 30147 6783
rect 30297 6749 30331 6783
rect 33333 6749 33367 6783
rect 35127 6749 35161 6783
rect 35265 6749 35299 6783
rect 35357 6749 35391 6783
rect 35541 6749 35575 6783
rect 37004 6749 37038 6783
rect 22744 6681 22778 6715
rect 25421 6681 25455 6715
rect 27077 6681 27111 6715
rect 15577 6613 15611 6647
rect 20085 6613 20119 6647
rect 25605 6613 25639 6647
rect 33425 6613 33459 6647
rect 20561 6409 20595 6443
rect 20729 6409 20763 6443
rect 23305 6409 23339 6443
rect 23673 6409 23707 6443
rect 24599 6409 24633 6443
rect 26249 6409 26283 6443
rect 28825 6409 28859 6443
rect 29285 6409 29319 6443
rect 30481 6409 30515 6443
rect 33977 6409 34011 6443
rect 20361 6341 20395 6375
rect 23765 6341 23799 6375
rect 24501 6341 24535 6375
rect 29653 6341 29687 6375
rect 33609 6341 33643 6375
rect 34805 6341 34839 6375
rect 38117 6341 38151 6375
rect 15577 6273 15611 6307
rect 16037 6273 16071 6307
rect 18153 6273 18187 6307
rect 18613 6273 18647 6307
rect 21189 6273 21223 6307
rect 21373 6273 21407 6307
rect 24685 6273 24719 6307
rect 24777 6273 24811 6307
rect 26065 6273 26099 6307
rect 26341 6273 26375 6307
rect 27712 6273 27746 6307
rect 30849 6273 30883 6307
rect 33793 6273 33827 6307
rect 35081 6273 35115 6307
rect 35173 6273 35207 6307
rect 35265 6273 35299 6307
rect 35449 6273 35483 6307
rect 37841 6273 37875 6307
rect 23949 6205 23983 6239
rect 27445 6205 27479 6239
rect 29745 6205 29779 6239
rect 29929 6205 29963 6239
rect 30941 6205 30975 6239
rect 31033 6205 31067 6239
rect 15669 6069 15703 6103
rect 20545 6069 20579 6103
rect 21189 6069 21223 6103
rect 25881 6069 25915 6103
rect 17141 5865 17175 5899
rect 25973 5865 26007 5899
rect 28089 5865 28123 5899
rect 35265 5865 35299 5899
rect 38301 5865 38335 5899
rect 22477 5797 22511 5831
rect 25881 5797 25915 5831
rect 20913 5729 20947 5763
rect 25053 5729 25087 5763
rect 25237 5729 25271 5763
rect 26065 5729 26099 5763
rect 28549 5729 28583 5763
rect 28641 5729 28675 5763
rect 34161 5729 34195 5763
rect 36921 5729 36955 5763
rect 15485 5661 15519 5695
rect 16037 5661 16071 5695
rect 18245 5661 18279 5695
rect 18429 5661 18463 5695
rect 21189 5661 21223 5695
rect 25789 5661 25823 5695
rect 28457 5661 28491 5695
rect 30481 5661 30515 5695
rect 33977 5661 34011 5695
rect 30726 5593 30760 5627
rect 34897 5593 34931 5627
rect 35081 5593 35115 5627
rect 37188 5593 37222 5627
rect 18337 5525 18371 5559
rect 24593 5525 24627 5559
rect 24961 5525 24995 5559
rect 31861 5525 31895 5559
rect 33609 5525 33643 5559
rect 34069 5525 34103 5559
rect 21281 5321 21315 5355
rect 23581 5321 23615 5355
rect 25421 5321 25455 5355
rect 30481 5321 30515 5355
rect 30849 5321 30883 5355
rect 33701 5321 33735 5355
rect 36645 5321 36679 5355
rect 37473 5321 37507 5355
rect 37841 5321 37875 5355
rect 18061 5253 18095 5287
rect 24308 5253 24342 5287
rect 26341 5253 26375 5287
rect 30941 5253 30975 5287
rect 37933 5253 37967 5287
rect 19717 5185 19751 5219
rect 22201 5185 22235 5219
rect 22468 5185 22502 5219
rect 26249 5185 26283 5219
rect 32321 5185 32355 5219
rect 32588 5185 32622 5219
rect 35532 5185 35566 5219
rect 19993 5117 20027 5151
rect 24041 5117 24075 5151
rect 26525 5117 26559 5151
rect 31033 5117 31067 5151
rect 35265 5117 35299 5151
rect 38025 5117 38059 5151
rect 18337 5049 18371 5083
rect 18521 4981 18555 5015
rect 25881 4981 25915 5015
rect 23029 4777 23063 4811
rect 26985 4777 27019 4811
rect 28825 4777 28859 4811
rect 31125 4777 31159 4811
rect 32597 4777 32631 4811
rect 35633 4777 35667 4811
rect 17509 4709 17543 4743
rect 16221 4641 16255 4675
rect 23581 4641 23615 4675
rect 33149 4641 33183 4675
rect 36093 4641 36127 4675
rect 36185 4641 36219 4675
rect 38117 4641 38151 4675
rect 15945 4573 15979 4607
rect 23397 4573 23431 4607
rect 25605 4573 25639 4607
rect 27445 4573 27479 4607
rect 29745 4573 29779 4607
rect 32965 4573 32999 4607
rect 36001 4573 36035 4607
rect 37841 4573 37875 4607
rect 25872 4505 25906 4539
rect 27712 4505 27746 4539
rect 30012 4505 30046 4539
rect 23489 4437 23523 4471
rect 33057 4437 33091 4471
rect 27905 4233 27939 4267
rect 28273 4233 28307 4267
rect 29929 4233 29963 4267
rect 30297 4233 30331 4267
rect 30389 4165 30423 4199
rect 18153 4097 18187 4131
rect 18429 4097 18463 4131
rect 28365 4097 28399 4131
rect 33609 4097 33643 4131
rect 33865 4097 33899 4131
rect 37841 4097 37875 4131
rect 38117 4097 38151 4131
rect 19533 4029 19567 4063
rect 28457 4029 28491 4063
rect 30481 4029 30515 4063
rect 34989 3893 35023 3927
rect 37841 3009 37875 3043
rect 38117 2941 38151 2975
rect 37841 2397 37875 2431
rect 38117 2329 38151 2363
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 9398 37272 9404 37324
rect 9456 37312 9462 37324
rect 9677 37315 9735 37321
rect 9677 37312 9689 37315
rect 9456 37284 9689 37312
rect 9456 37272 9462 37284
rect 9677 37281 9689 37284
rect 9723 37281 9735 37315
rect 12158 37312 12164 37324
rect 12119 37284 12164 37312
rect 9677 37275 9735 37281
rect 12158 37272 12164 37284
rect 12216 37272 12222 37324
rect 26510 37312 26516 37324
rect 26471 37284 26516 37312
rect 26510 37272 26516 37284
rect 26568 37272 26574 37324
rect 28074 37272 28080 37324
rect 28132 37312 28138 37324
rect 28629 37315 28687 37321
rect 28629 37312 28641 37315
rect 28132 37284 28641 37312
rect 28132 37272 28138 37284
rect 28629 37281 28641 37284
rect 28675 37281 28687 37315
rect 28629 37275 28687 37281
rect 30466 37272 30472 37324
rect 30524 37312 30530 37324
rect 32585 37315 32643 37321
rect 32585 37312 32597 37315
rect 30524 37284 32597 37312
rect 30524 37272 30530 37284
rect 32585 37281 32597 37284
rect 32631 37281 32643 37315
rect 32585 37275 32643 37281
rect 32674 37272 32680 37324
rect 32732 37312 32738 37324
rect 33597 37315 33655 37321
rect 33597 37312 33609 37315
rect 32732 37284 33609 37312
rect 32732 37272 32738 37284
rect 33597 37281 33609 37284
rect 33643 37281 33655 37315
rect 33597 37275 33655 37281
rect 1762 37204 1768 37256
rect 1820 37244 1826 37256
rect 1857 37247 1915 37253
rect 1857 37244 1869 37247
rect 1820 37216 1869 37244
rect 1820 37204 1826 37216
rect 1857 37213 1869 37216
rect 1903 37213 1915 37247
rect 5074 37244 5080 37256
rect 5035 37216 5080 37244
rect 1857 37207 1915 37213
rect 5074 37204 5080 37216
rect 5132 37204 5138 37256
rect 7929 37247 7987 37253
rect 7929 37213 7941 37247
rect 7975 37244 7987 37247
rect 8386 37244 8392 37256
rect 7975 37216 8392 37244
rect 7975 37213 7987 37216
rect 7929 37207 7987 37213
rect 8386 37204 8392 37216
rect 8444 37204 8450 37256
rect 11698 37204 11704 37256
rect 11756 37244 11762 37256
rect 11793 37247 11851 37253
rect 11793 37244 11805 37247
rect 11756 37216 11805 37244
rect 11756 37204 11762 37216
rect 11793 37213 11805 37216
rect 11839 37213 11851 37247
rect 15194 37244 15200 37256
rect 15155 37216 15200 37244
rect 11793 37207 11851 37213
rect 15194 37204 15200 37216
rect 15252 37204 15258 37256
rect 18233 37247 18291 37253
rect 15672 37216 17816 37244
rect 2685 37179 2743 37185
rect 2685 37145 2697 37179
rect 2731 37176 2743 37179
rect 5534 37176 5540 37188
rect 2731 37148 5540 37176
rect 2731 37145 2743 37148
rect 2685 37139 2743 37145
rect 5534 37136 5540 37148
rect 5592 37136 5598 37188
rect 5718 37136 5724 37188
rect 5776 37176 5782 37188
rect 5813 37179 5871 37185
rect 5813 37176 5825 37179
rect 5776 37148 5825 37176
rect 5776 37136 5782 37148
rect 5813 37145 5825 37148
rect 5859 37145 5871 37179
rect 5813 37139 5871 37145
rect 8481 37179 8539 37185
rect 8481 37145 8493 37179
rect 8527 37176 8539 37179
rect 9306 37176 9312 37188
rect 8527 37148 9312 37176
rect 8527 37145 8539 37148
rect 8481 37139 8539 37145
rect 9306 37136 9312 37148
rect 9364 37136 9370 37188
rect 9490 37176 9496 37188
rect 9403 37148 9496 37176
rect 9490 37136 9496 37148
rect 9548 37176 9554 37188
rect 15672 37176 15700 37216
rect 9548 37148 15700 37176
rect 15749 37179 15807 37185
rect 9548 37136 9554 37148
rect 15749 37145 15761 37179
rect 15795 37176 15807 37179
rect 16022 37176 16028 37188
rect 15795 37148 16028 37176
rect 15795 37145 15807 37148
rect 15749 37139 15807 37145
rect 16022 37136 16028 37148
rect 16080 37136 16086 37188
rect 17788 37176 17816 37216
rect 18233 37213 18245 37247
rect 18279 37244 18291 37247
rect 18322 37244 18328 37256
rect 18279 37216 18328 37244
rect 18279 37213 18291 37216
rect 18233 37207 18291 37213
rect 18322 37204 18328 37216
rect 18380 37204 18386 37256
rect 22094 37204 22100 37256
rect 22152 37244 22158 37256
rect 22152 37216 22197 37244
rect 22152 37204 22158 37216
rect 24946 37204 24952 37256
rect 25004 37244 25010 37256
rect 25133 37247 25191 37253
rect 25133 37244 25145 37247
rect 25004 37216 25145 37244
rect 25004 37204 25010 37216
rect 25133 37213 25145 37216
rect 25179 37213 25191 37247
rect 25133 37207 25191 37213
rect 26234 37204 26240 37256
rect 26292 37244 26298 37256
rect 26421 37247 26479 37253
rect 26421 37244 26433 37247
rect 26292 37216 26433 37244
rect 26292 37204 26298 37216
rect 26421 37213 26433 37216
rect 26467 37213 26479 37247
rect 26421 37207 26479 37213
rect 26605 37247 26663 37253
rect 26605 37213 26617 37247
rect 26651 37244 26663 37247
rect 27430 37244 27436 37256
rect 26651 37216 27436 37244
rect 26651 37213 26663 37216
rect 26605 37207 26663 37213
rect 27430 37204 27436 37216
rect 27488 37204 27494 37256
rect 28258 37204 28264 37256
rect 28316 37244 28322 37256
rect 28445 37247 28503 37253
rect 28445 37244 28457 37247
rect 28316 37216 28457 37244
rect 28316 37204 28322 37216
rect 28445 37213 28457 37216
rect 28491 37213 28503 37247
rect 28445 37207 28503 37213
rect 31754 37204 31760 37256
rect 31812 37244 31818 37256
rect 32401 37247 32459 37253
rect 32401 37244 32413 37247
rect 31812 37216 32413 37244
rect 31812 37204 31818 37216
rect 32401 37213 32413 37216
rect 32447 37213 32459 37247
rect 33778 37244 33784 37256
rect 33739 37216 33784 37244
rect 32401 37207 32459 37213
rect 33778 37204 33784 37216
rect 33836 37204 33842 37256
rect 36446 37244 36452 37256
rect 36407 37216 36452 37244
rect 36446 37204 36452 37216
rect 36504 37204 36510 37256
rect 37645 37247 37703 37253
rect 37645 37213 37657 37247
rect 37691 37244 37703 37247
rect 38102 37244 38108 37256
rect 37691 37216 38108 37244
rect 37691 37213 37703 37216
rect 37645 37207 37703 37213
rect 38102 37204 38108 37216
rect 38160 37204 38166 37256
rect 18598 37176 18604 37188
rect 17788 37148 18604 37176
rect 18598 37136 18604 37148
rect 18656 37136 18662 37188
rect 22833 37179 22891 37185
rect 22833 37176 22845 37179
rect 22066 37148 22845 37176
rect 9122 37108 9128 37120
rect 9083 37080 9128 37108
rect 9122 37068 9128 37080
rect 9180 37068 9186 37120
rect 9582 37068 9588 37120
rect 9640 37108 9646 37120
rect 9640 37080 9685 37108
rect 9640 37068 9646 37080
rect 12986 37068 12992 37120
rect 13044 37108 13050 37120
rect 22066 37108 22094 37148
rect 22833 37145 22845 37148
rect 22879 37176 22891 37179
rect 24302 37176 24308 37188
rect 22879 37148 24308 37176
rect 22879 37145 22891 37148
rect 22833 37139 22891 37145
rect 24302 37136 24308 37148
rect 24360 37136 24366 37188
rect 25501 37179 25559 37185
rect 25501 37145 25513 37179
rect 25547 37145 25559 37179
rect 36722 37176 36728 37188
rect 36683 37148 36728 37176
rect 25501 37139 25559 37145
rect 13044 37080 22094 37108
rect 13044 37068 13050 37080
rect 22462 37068 22468 37120
rect 22520 37108 22526 37120
rect 25516 37108 25544 37139
rect 36722 37136 36728 37148
rect 36780 37136 36786 37188
rect 38010 37176 38016 37188
rect 37971 37148 38016 37176
rect 38010 37136 38016 37148
rect 38068 37136 38074 37188
rect 28442 37108 28448 37120
rect 22520 37080 28448 37108
rect 22520 37068 22526 37080
rect 28442 37068 28448 37080
rect 28500 37108 28506 37120
rect 31018 37108 31024 37120
rect 28500 37080 31024 37108
rect 28500 37068 28506 37080
rect 31018 37068 31024 37080
rect 31076 37068 31082 37120
rect 33962 37108 33968 37120
rect 33923 37080 33968 37108
rect 33962 37068 33968 37080
rect 34020 37068 34026 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 6549 36907 6607 36913
rect 6549 36873 6561 36907
rect 6595 36873 6607 36907
rect 6549 36867 6607 36873
rect 9309 36907 9367 36913
rect 9309 36873 9321 36907
rect 9355 36904 9367 36907
rect 9582 36904 9588 36916
rect 9355 36876 9588 36904
rect 9355 36873 9367 36876
rect 9309 36867 9367 36873
rect 4700 36839 4758 36845
rect 4700 36805 4712 36839
rect 4746 36836 4758 36839
rect 6564 36836 6592 36867
rect 9582 36864 9588 36876
rect 9640 36864 9646 36916
rect 14292 36876 15884 36904
rect 4746 36808 6592 36836
rect 8196 36839 8254 36845
rect 4746 36805 4758 36808
rect 4700 36799 4758 36805
rect 8196 36805 8208 36839
rect 8242 36836 8254 36839
rect 9122 36836 9128 36848
rect 8242 36808 9128 36836
rect 8242 36805 8254 36808
rect 8196 36799 8254 36805
rect 9122 36796 9128 36808
rect 9180 36796 9186 36848
rect 12084 36808 13400 36836
rect 4433 36771 4491 36777
rect 4433 36737 4445 36771
rect 4479 36768 4491 36771
rect 4522 36768 4528 36780
rect 4479 36740 4528 36768
rect 4479 36737 4491 36740
rect 4433 36731 4491 36737
rect 4522 36728 4528 36740
rect 4580 36728 4586 36780
rect 5534 36728 5540 36780
rect 5592 36768 5598 36780
rect 6917 36771 6975 36777
rect 6917 36768 6929 36771
rect 5592 36740 6929 36768
rect 5592 36728 5598 36740
rect 6917 36737 6929 36740
rect 6963 36768 6975 36771
rect 11514 36768 11520 36780
rect 6963 36740 11520 36768
rect 6963 36737 6975 36740
rect 6917 36731 6975 36737
rect 11514 36728 11520 36740
rect 11572 36728 11578 36780
rect 12084 36777 12112 36808
rect 13372 36780 13400 36808
rect 12069 36771 12127 36777
rect 12069 36737 12081 36771
rect 12115 36737 12127 36771
rect 12069 36731 12127 36737
rect 12336 36771 12394 36777
rect 12336 36737 12348 36771
rect 12382 36768 12394 36771
rect 12618 36768 12624 36780
rect 12382 36740 12624 36768
rect 12382 36737 12394 36740
rect 12336 36731 12394 36737
rect 12618 36728 12624 36740
rect 12676 36728 12682 36780
rect 13354 36728 13360 36780
rect 13412 36768 13418 36780
rect 14292 36777 14320 36876
rect 15856 36848 15884 36876
rect 17788 36876 22048 36904
rect 15286 36796 15292 36848
rect 15344 36796 15350 36848
rect 15838 36796 15844 36848
rect 15896 36836 15902 36848
rect 17788 36836 17816 36876
rect 15896 36808 17816 36836
rect 15896 36796 15902 36808
rect 14277 36771 14335 36777
rect 14277 36768 14289 36771
rect 13412 36740 14289 36768
rect 13412 36728 13418 36740
rect 14277 36737 14289 36740
rect 14323 36737 14335 36771
rect 14277 36731 14335 36737
rect 16482 36728 16488 36780
rect 16540 36768 16546 36780
rect 17788 36777 17816 36808
rect 20180 36808 21956 36836
rect 16853 36771 16911 36777
rect 16853 36768 16865 36771
rect 16540 36740 16865 36768
rect 16540 36728 16546 36740
rect 16853 36737 16865 36740
rect 16899 36737 16911 36771
rect 16853 36731 16911 36737
rect 17773 36771 17831 36777
rect 17773 36737 17785 36771
rect 17819 36737 17831 36771
rect 19518 36768 19524 36780
rect 19182 36740 19524 36768
rect 17773 36731 17831 36737
rect 19518 36728 19524 36740
rect 19576 36728 19582 36780
rect 19978 36728 19984 36780
rect 20036 36768 20042 36780
rect 20180 36768 20208 36808
rect 20036 36754 20208 36768
rect 20036 36740 20194 36754
rect 20036 36728 20042 36740
rect 7009 36703 7067 36709
rect 7009 36700 7021 36703
rect 5828 36672 7021 36700
rect 5626 36592 5632 36644
rect 5684 36632 5690 36644
rect 5828 36641 5856 36672
rect 7009 36669 7021 36672
rect 7055 36669 7067 36703
rect 7009 36663 7067 36669
rect 7193 36703 7251 36709
rect 7193 36669 7205 36703
rect 7239 36700 7251 36703
rect 7650 36700 7656 36712
rect 7239 36672 7656 36700
rect 7239 36669 7251 36672
rect 7193 36663 7251 36669
rect 7650 36660 7656 36672
rect 7708 36660 7714 36712
rect 7926 36700 7932 36712
rect 7887 36672 7932 36700
rect 7926 36660 7932 36672
rect 7984 36660 7990 36712
rect 14550 36700 14556 36712
rect 14511 36672 14556 36700
rect 14550 36660 14556 36672
rect 14608 36660 14614 36712
rect 18046 36700 18052 36712
rect 18007 36672 18052 36700
rect 18046 36660 18052 36672
rect 18104 36660 18110 36712
rect 20257 36703 20315 36709
rect 20257 36669 20269 36703
rect 20303 36700 20315 36703
rect 20806 36700 20812 36712
rect 20303 36672 20812 36700
rect 20303 36669 20315 36672
rect 20257 36663 20315 36669
rect 20806 36660 20812 36672
rect 20864 36660 20870 36712
rect 20993 36703 21051 36709
rect 20993 36669 21005 36703
rect 21039 36669 21051 36703
rect 20993 36663 21051 36669
rect 5813 36635 5871 36641
rect 5813 36632 5825 36635
rect 5684 36604 5825 36632
rect 5684 36592 5690 36604
rect 5813 36601 5825 36604
rect 5859 36601 5871 36635
rect 5813 36595 5871 36601
rect 16025 36635 16083 36641
rect 16025 36601 16037 36635
rect 16071 36632 16083 36635
rect 17678 36632 17684 36644
rect 16071 36604 17684 36632
rect 16071 36601 16083 36604
rect 16025 36595 16083 36601
rect 17678 36592 17684 36604
rect 17736 36592 17742 36644
rect 20070 36592 20076 36644
rect 20128 36632 20134 36644
rect 21008 36632 21036 36663
rect 20128 36604 21036 36632
rect 20128 36592 20134 36604
rect 13078 36524 13084 36576
rect 13136 36564 13142 36576
rect 13449 36567 13507 36573
rect 13449 36564 13461 36567
rect 13136 36536 13461 36564
rect 13136 36524 13142 36536
rect 13449 36533 13461 36536
rect 13495 36533 13507 36567
rect 16942 36564 16948 36576
rect 16903 36536 16948 36564
rect 13449 36527 13507 36533
rect 16942 36524 16948 36536
rect 17000 36524 17006 36576
rect 19521 36567 19579 36573
rect 19521 36533 19533 36567
rect 19567 36564 19579 36567
rect 19886 36564 19892 36576
rect 19567 36536 19892 36564
rect 19567 36533 19579 36536
rect 19521 36527 19579 36533
rect 19886 36524 19892 36536
rect 19944 36524 19950 36576
rect 21928 36564 21956 36808
rect 22020 36777 22048 36876
rect 23952 36876 27568 36904
rect 22005 36771 22063 36777
rect 22005 36737 22017 36771
rect 22051 36737 22063 36771
rect 22005 36731 22063 36737
rect 22094 36728 22100 36780
rect 22152 36768 22158 36780
rect 23952 36777 23980 36876
rect 26329 36839 26387 36845
rect 26329 36836 26341 36839
rect 25438 36808 26341 36836
rect 26329 36805 26341 36808
rect 26375 36805 26387 36839
rect 27540 36836 27568 36876
rect 28350 36864 28356 36916
rect 28408 36904 28414 36916
rect 38010 36904 38016 36916
rect 28408 36876 38016 36904
rect 28408 36864 28414 36876
rect 38010 36864 38016 36876
rect 38068 36864 38074 36916
rect 27614 36836 27620 36848
rect 27527 36808 27620 36836
rect 26329 36799 26387 36805
rect 22261 36771 22319 36777
rect 22261 36768 22273 36771
rect 22152 36740 22273 36768
rect 22152 36728 22158 36740
rect 22261 36737 22273 36740
rect 22307 36737 22319 36771
rect 22261 36731 22319 36737
rect 23937 36771 23995 36777
rect 23937 36737 23949 36771
rect 23983 36737 23995 36771
rect 23937 36731 23995 36737
rect 26237 36771 26295 36777
rect 26237 36737 26249 36771
rect 26283 36768 26295 36771
rect 26418 36768 26424 36780
rect 26283 36740 26424 36768
rect 26283 36737 26295 36740
rect 26237 36731 26295 36737
rect 26418 36728 26424 36740
rect 26476 36768 26482 36780
rect 27540 36777 27568 36808
rect 27614 36796 27620 36808
rect 27672 36836 27678 36848
rect 32766 36836 32772 36848
rect 27672 36808 28672 36836
rect 27672 36796 27678 36808
rect 28644 36780 28672 36808
rect 29472 36808 32772 36836
rect 27525 36771 27583 36777
rect 26476 36740 27200 36768
rect 26476 36728 26482 36740
rect 23014 36660 23020 36712
rect 23072 36700 23078 36712
rect 24213 36703 24271 36709
rect 24213 36700 24225 36703
rect 23072 36672 24225 36700
rect 23072 36660 23078 36672
rect 24213 36669 24225 36672
rect 24259 36669 24271 36703
rect 24213 36663 24271 36669
rect 24302 36660 24308 36712
rect 24360 36700 24366 36712
rect 27062 36700 27068 36712
rect 24360 36672 27068 36700
rect 24360 36660 24366 36672
rect 27062 36660 27068 36672
rect 27120 36660 27126 36712
rect 23216 36604 24072 36632
rect 23216 36564 23244 36604
rect 23382 36564 23388 36576
rect 21928 36536 23244 36564
rect 23343 36536 23388 36564
rect 23382 36524 23388 36536
rect 23440 36524 23446 36576
rect 24044 36564 24072 36604
rect 25682 36564 25688 36576
rect 24044 36536 25688 36564
rect 25682 36524 25688 36536
rect 25740 36524 25746 36576
rect 27172 36564 27200 36740
rect 27525 36737 27537 36771
rect 27571 36737 27583 36771
rect 27525 36731 27583 36737
rect 27792 36771 27850 36777
rect 27792 36737 27804 36771
rect 27838 36768 27850 36771
rect 28166 36768 28172 36780
rect 27838 36740 28172 36768
rect 27838 36737 27850 36740
rect 27792 36731 27850 36737
rect 28166 36728 28172 36740
rect 28224 36728 28230 36780
rect 28626 36728 28632 36780
rect 28684 36768 28690 36780
rect 29472 36777 29500 36808
rect 29457 36771 29515 36777
rect 29457 36768 29469 36771
rect 28684 36740 29469 36768
rect 28684 36728 28690 36740
rect 29457 36737 29469 36740
rect 29503 36737 29515 36771
rect 29457 36731 29515 36737
rect 29724 36771 29782 36777
rect 29724 36737 29736 36771
rect 29770 36768 29782 36771
rect 30466 36768 30472 36780
rect 29770 36740 30472 36768
rect 29770 36737 29782 36740
rect 29724 36731 29782 36737
rect 30466 36728 30472 36740
rect 30524 36728 30530 36780
rect 32324 36777 32352 36808
rect 32766 36796 32772 36808
rect 32824 36796 32830 36848
rect 33962 36796 33968 36848
rect 34020 36836 34026 36848
rect 34486 36839 34544 36845
rect 34486 36836 34498 36839
rect 34020 36808 34498 36836
rect 34020 36796 34026 36808
rect 34486 36805 34498 36808
rect 34532 36805 34544 36839
rect 34486 36799 34544 36805
rect 36725 36839 36783 36845
rect 36725 36805 36737 36839
rect 36771 36836 36783 36839
rect 36814 36836 36820 36848
rect 36771 36808 36820 36836
rect 36771 36805 36783 36808
rect 36725 36799 36783 36805
rect 36814 36796 36820 36808
rect 36872 36796 36878 36848
rect 32309 36771 32367 36777
rect 32309 36737 32321 36771
rect 32355 36737 32367 36771
rect 32309 36731 32367 36737
rect 32398 36728 32404 36780
rect 32456 36768 32462 36780
rect 32565 36771 32623 36777
rect 32565 36768 32577 36771
rect 32456 36740 32577 36768
rect 32456 36728 32462 36740
rect 32565 36737 32577 36740
rect 32611 36737 32623 36771
rect 32565 36731 32623 36737
rect 35986 36728 35992 36780
rect 36044 36768 36050 36780
rect 36449 36771 36507 36777
rect 36449 36768 36461 36771
rect 36044 36740 36461 36768
rect 36044 36728 36050 36740
rect 36449 36737 36461 36740
rect 36495 36737 36507 36771
rect 36449 36731 36507 36737
rect 37734 36728 37740 36780
rect 37792 36768 37798 36780
rect 37829 36771 37887 36777
rect 37829 36768 37841 36771
rect 37792 36740 37841 36768
rect 37792 36728 37798 36740
rect 37829 36737 37841 36740
rect 37875 36737 37887 36771
rect 37829 36731 37887 36737
rect 34238 36700 34244 36712
rect 34199 36672 34244 36700
rect 34238 36660 34244 36672
rect 34296 36660 34302 36712
rect 38102 36700 38108 36712
rect 38063 36672 38108 36700
rect 38102 36660 38108 36672
rect 38160 36660 38166 36712
rect 28258 36564 28264 36576
rect 27172 36536 28264 36564
rect 28258 36524 28264 36536
rect 28316 36524 28322 36576
rect 28905 36567 28963 36573
rect 28905 36533 28917 36567
rect 28951 36564 28963 36567
rect 29270 36564 29276 36576
rect 28951 36536 29276 36564
rect 28951 36533 28963 36536
rect 28905 36527 28963 36533
rect 29270 36524 29276 36536
rect 29328 36524 29334 36576
rect 30098 36524 30104 36576
rect 30156 36564 30162 36576
rect 30837 36567 30895 36573
rect 30837 36564 30849 36567
rect 30156 36536 30849 36564
rect 30156 36524 30162 36536
rect 30837 36533 30849 36536
rect 30883 36533 30895 36567
rect 33686 36564 33692 36576
rect 33647 36536 33692 36564
rect 30837 36527 30895 36533
rect 33686 36524 33692 36536
rect 33744 36524 33750 36576
rect 35618 36564 35624 36576
rect 35579 36536 35624 36564
rect 35618 36524 35624 36536
rect 35676 36524 35682 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 12618 36360 12624 36372
rect 12579 36332 12624 36360
rect 12618 36320 12624 36332
rect 12676 36320 12682 36372
rect 15286 36360 15292 36372
rect 15247 36332 15292 36360
rect 15286 36320 15292 36332
rect 15344 36320 15350 36372
rect 19518 36360 19524 36372
rect 15396 36332 16988 36360
rect 19479 36332 19524 36360
rect 8570 36252 8576 36304
rect 8628 36292 8634 36304
rect 9217 36295 9275 36301
rect 9217 36292 9229 36295
rect 8628 36264 9229 36292
rect 8628 36252 8634 36264
rect 9217 36261 9229 36264
rect 9263 36261 9275 36295
rect 9217 36255 9275 36261
rect 9306 36252 9312 36304
rect 9364 36292 9370 36304
rect 9364 36264 9720 36292
rect 9364 36252 9370 36264
rect 5626 36224 5632 36236
rect 5587 36196 5632 36224
rect 5626 36184 5632 36196
rect 5684 36184 5690 36236
rect 5813 36227 5871 36233
rect 5813 36193 5825 36227
rect 5859 36224 5871 36227
rect 5902 36224 5908 36236
rect 5859 36196 5908 36224
rect 5859 36193 5871 36196
rect 5813 36187 5871 36193
rect 5902 36184 5908 36196
rect 5960 36184 5966 36236
rect 9490 36184 9496 36236
rect 9548 36224 9554 36236
rect 9585 36227 9643 36233
rect 9585 36224 9597 36227
rect 9548 36196 9597 36224
rect 9548 36184 9554 36196
rect 9585 36193 9597 36196
rect 9631 36193 9643 36227
rect 9692 36224 9720 36264
rect 11514 36252 11520 36304
rect 11572 36292 11578 36304
rect 13998 36292 14004 36304
rect 11572 36264 14004 36292
rect 11572 36252 11578 36264
rect 13998 36252 14004 36264
rect 14056 36252 14062 36304
rect 13078 36224 13084 36236
rect 9692 36196 10640 36224
rect 13039 36196 13084 36224
rect 9585 36187 9643 36193
rect 4614 36116 4620 36168
rect 4672 36156 4678 36168
rect 6365 36159 6423 36165
rect 6365 36156 6377 36159
rect 4672 36128 6377 36156
rect 4672 36116 4678 36128
rect 6365 36125 6377 36128
rect 6411 36156 6423 36159
rect 7926 36156 7932 36168
rect 6411 36128 7932 36156
rect 6411 36125 6423 36128
rect 6365 36119 6423 36125
rect 7926 36116 7932 36128
rect 7984 36156 7990 36168
rect 9674 36156 9680 36168
rect 7984 36128 9680 36156
rect 7984 36116 7990 36128
rect 9674 36116 9680 36128
rect 9732 36156 9738 36168
rect 10505 36159 10563 36165
rect 10505 36156 10517 36159
rect 9732 36128 10517 36156
rect 9732 36116 9738 36128
rect 10505 36125 10517 36128
rect 10551 36125 10563 36159
rect 10612 36156 10640 36196
rect 13078 36184 13084 36196
rect 13136 36184 13142 36236
rect 13262 36224 13268 36236
rect 13223 36196 13268 36224
rect 13262 36184 13268 36196
rect 13320 36184 13326 36236
rect 13538 36184 13544 36236
rect 13596 36224 13602 36236
rect 15396 36224 15424 36332
rect 16960 36292 16988 36332
rect 19518 36320 19524 36332
rect 19576 36320 19582 36372
rect 27430 36360 27436 36372
rect 23216 36332 27436 36360
rect 23216 36292 23244 36332
rect 27430 36320 27436 36332
rect 27488 36320 27494 36372
rect 28166 36360 28172 36372
rect 28127 36332 28172 36360
rect 28166 36320 28172 36332
rect 28224 36320 28230 36372
rect 30098 36360 30104 36372
rect 30059 36332 30104 36360
rect 30098 36320 30104 36332
rect 30156 36320 30162 36372
rect 31573 36363 31631 36369
rect 31573 36329 31585 36363
rect 31619 36360 31631 36363
rect 32398 36360 32404 36372
rect 31619 36332 32404 36360
rect 31619 36329 31631 36332
rect 31573 36323 31631 36329
rect 32398 36320 32404 36332
rect 32456 36320 32462 36372
rect 32674 36360 32680 36372
rect 32635 36332 32680 36360
rect 32674 36320 32680 36332
rect 32732 36320 32738 36372
rect 33597 36363 33655 36369
rect 33597 36329 33609 36363
rect 33643 36360 33655 36363
rect 33778 36360 33784 36372
rect 33643 36332 33784 36360
rect 33643 36329 33655 36332
rect 33597 36323 33655 36329
rect 33778 36320 33784 36332
rect 33836 36320 33842 36372
rect 16960 36264 20760 36292
rect 15838 36224 15844 36236
rect 13596 36196 15424 36224
rect 15799 36196 15844 36224
rect 13596 36184 13602 36196
rect 15838 36184 15844 36196
rect 15896 36184 15902 36236
rect 16482 36224 16488 36236
rect 16040 36196 16488 36224
rect 10612 36128 12434 36156
rect 10505 36119 10563 36125
rect 5534 36088 5540 36100
rect 5495 36060 5540 36088
rect 5534 36048 5540 36060
rect 5592 36048 5598 36100
rect 6632 36091 6690 36097
rect 6632 36057 6644 36091
rect 6678 36088 6690 36091
rect 7098 36088 7104 36100
rect 6678 36060 7104 36088
rect 6678 36057 6690 36060
rect 6632 36051 6690 36057
rect 7098 36048 7104 36060
rect 7156 36048 7162 36100
rect 7834 36048 7840 36100
rect 7892 36088 7898 36100
rect 9769 36091 9827 36097
rect 9769 36088 9781 36091
rect 7892 36060 9781 36088
rect 7892 36048 7898 36060
rect 9769 36057 9781 36060
rect 9815 36057 9827 36091
rect 9769 36051 9827 36057
rect 10772 36091 10830 36097
rect 10772 36057 10784 36091
rect 10818 36088 10830 36091
rect 11698 36088 11704 36100
rect 10818 36060 11704 36088
rect 10818 36057 10830 36060
rect 10772 36051 10830 36057
rect 11698 36048 11704 36060
rect 11756 36048 11762 36100
rect 5169 36023 5227 36029
rect 5169 35989 5181 36023
rect 5215 36020 5227 36023
rect 5258 36020 5264 36032
rect 5215 35992 5264 36020
rect 5215 35989 5227 35992
rect 5169 35983 5227 35989
rect 5258 35980 5264 35992
rect 5316 35980 5322 36032
rect 7742 36020 7748 36032
rect 7703 35992 7748 36020
rect 7742 35980 7748 35992
rect 7800 35980 7806 36032
rect 9582 35980 9588 36032
rect 9640 36020 9646 36032
rect 9677 36023 9735 36029
rect 9677 36020 9689 36023
rect 9640 35992 9689 36020
rect 9640 35980 9646 35992
rect 9677 35989 9689 35992
rect 9723 35989 9735 36023
rect 11882 36020 11888 36032
rect 11843 35992 11888 36020
rect 9677 35983 9735 35989
rect 11882 35980 11888 35992
rect 11940 35980 11946 36032
rect 12406 36020 12434 36128
rect 12710 36116 12716 36168
rect 12768 36156 12774 36168
rect 12986 36156 12992 36168
rect 12768 36128 12992 36156
rect 12768 36116 12774 36128
rect 12986 36116 12992 36128
rect 13044 36116 13050 36168
rect 15194 36156 15200 36168
rect 15107 36128 15200 36156
rect 15194 36116 15200 36128
rect 15252 36156 15258 36168
rect 16040 36156 16068 36196
rect 16482 36184 16488 36196
rect 16540 36224 16546 36236
rect 20622 36224 20628 36236
rect 16540 36196 20628 36224
rect 16540 36184 16546 36196
rect 16206 36156 16212 36168
rect 15252 36128 16068 36156
rect 16167 36128 16212 36156
rect 15252 36116 15258 36128
rect 16206 36116 16212 36128
rect 16264 36116 16270 36168
rect 18414 36156 18420 36168
rect 18375 36128 18420 36156
rect 18414 36116 18420 36128
rect 18472 36116 18478 36168
rect 19444 36165 19472 36196
rect 20622 36184 20628 36196
rect 20680 36184 20686 36236
rect 20732 36224 20760 36264
rect 22066 36264 23244 36292
rect 22066 36224 22094 36264
rect 20732 36196 22094 36224
rect 23216 36210 23244 36264
rect 24854 36252 24860 36304
rect 24912 36292 24918 36304
rect 25133 36295 25191 36301
rect 25133 36292 25145 36295
rect 24912 36264 25145 36292
rect 24912 36252 24918 36264
rect 25133 36261 25145 36264
rect 25179 36261 25191 36295
rect 25133 36255 25191 36261
rect 27062 36252 27068 36304
rect 27120 36292 27126 36304
rect 32306 36292 32312 36304
rect 27120 36264 32312 36292
rect 27120 36252 27126 36264
rect 32306 36252 32312 36264
rect 32364 36252 32370 36304
rect 23937 36227 23995 36233
rect 23937 36193 23949 36227
rect 23983 36224 23995 36227
rect 24946 36224 24952 36236
rect 23983 36196 24952 36224
rect 23983 36193 23995 36196
rect 23937 36187 23995 36193
rect 24946 36184 24952 36196
rect 25004 36224 25010 36236
rect 25225 36227 25283 36233
rect 25225 36224 25237 36227
rect 25004 36196 25237 36224
rect 25004 36184 25010 36196
rect 25225 36193 25237 36196
rect 25271 36193 25283 36227
rect 25225 36187 25283 36193
rect 26053 36227 26111 36233
rect 26053 36193 26065 36227
rect 26099 36224 26111 36227
rect 27614 36224 27620 36236
rect 26099 36196 27620 36224
rect 26099 36193 26111 36196
rect 26053 36187 26111 36193
rect 27614 36184 27620 36196
rect 27672 36184 27678 36236
rect 30466 36224 30472 36236
rect 29748 36196 30472 36224
rect 19429 36159 19487 36165
rect 19429 36125 19441 36159
rect 19475 36125 19487 36159
rect 19429 36119 19487 36125
rect 19886 36116 19892 36168
rect 19944 36156 19950 36168
rect 20257 36159 20315 36165
rect 20257 36156 20269 36159
rect 19944 36128 20269 36156
rect 19944 36116 19950 36128
rect 20257 36125 20269 36128
rect 20303 36156 20315 36159
rect 20438 36156 20444 36168
rect 20303 36128 20444 36156
rect 20303 36125 20315 36128
rect 20257 36119 20315 36125
rect 20438 36116 20444 36128
rect 20496 36116 20502 36168
rect 22922 36116 22928 36168
rect 22980 36156 22986 36168
rect 23382 36156 23388 36168
rect 22980 36128 23388 36156
rect 22980 36116 22986 36128
rect 23382 36116 23388 36128
rect 23440 36116 23446 36168
rect 24670 36156 24676 36168
rect 24631 36128 24676 36156
rect 24670 36116 24676 36128
rect 24728 36116 24734 36168
rect 24765 36159 24823 36165
rect 24765 36125 24777 36159
rect 24811 36125 24823 36159
rect 26326 36156 26332 36168
rect 26287 36128 26332 36156
rect 24765 36119 24823 36125
rect 16942 36048 16948 36100
rect 17000 36048 17006 36100
rect 18230 36048 18236 36100
rect 18288 36088 18294 36100
rect 18693 36091 18751 36097
rect 18693 36088 18705 36091
rect 18288 36060 18705 36088
rect 18288 36048 18294 36060
rect 18693 36057 18705 36060
rect 18739 36057 18751 36091
rect 18693 36051 18751 36057
rect 20533 36091 20591 36097
rect 20533 36057 20545 36091
rect 20579 36088 20591 36091
rect 20806 36088 20812 36100
rect 20579 36060 20812 36088
rect 20579 36057 20591 36060
rect 20533 36051 20591 36057
rect 20806 36048 20812 36060
rect 20864 36048 20870 36100
rect 20990 36048 20996 36100
rect 21048 36088 21054 36100
rect 21453 36091 21511 36097
rect 21453 36088 21465 36091
rect 21048 36060 21465 36088
rect 21048 36048 21054 36060
rect 21453 36057 21465 36060
rect 21499 36057 21511 36091
rect 23750 36088 23756 36100
rect 23711 36060 23756 36088
rect 21453 36051 21511 36057
rect 23750 36048 23756 36060
rect 23808 36048 23814 36100
rect 23842 36048 23848 36100
rect 23900 36088 23906 36100
rect 24780 36088 24808 36119
rect 26326 36116 26332 36128
rect 26384 36116 26390 36168
rect 28350 36156 28356 36168
rect 28311 36128 28356 36156
rect 28350 36116 28356 36128
rect 28408 36116 28414 36168
rect 29748 36165 29776 36196
rect 30466 36184 30472 36196
rect 30524 36184 30530 36236
rect 31202 36224 31208 36236
rect 31163 36196 31208 36224
rect 31202 36184 31208 36196
rect 31260 36184 31266 36236
rect 32692 36224 32720 36320
rect 31726 36196 32720 36224
rect 28629 36159 28687 36165
rect 28629 36156 28641 36159
rect 28460 36128 28641 36156
rect 23900 36060 24808 36088
rect 23900 36048 23906 36060
rect 27522 36048 27528 36100
rect 27580 36088 27586 36100
rect 28460 36088 28488 36128
rect 28629 36125 28641 36128
rect 28675 36125 28687 36159
rect 28629 36119 28687 36125
rect 29733 36159 29791 36165
rect 29733 36125 29745 36159
rect 29779 36125 29791 36159
rect 30006 36156 30012 36168
rect 29967 36128 30012 36156
rect 29733 36119 29791 36125
rect 30006 36116 30012 36128
rect 30064 36116 30070 36168
rect 31297 36159 31355 36165
rect 31297 36125 31309 36159
rect 31343 36156 31355 36159
rect 31726 36156 31754 36196
rect 34238 36184 34244 36236
rect 34296 36224 34302 36236
rect 34885 36227 34943 36233
rect 34885 36224 34897 36227
rect 34296 36196 34897 36224
rect 34296 36184 34302 36196
rect 34885 36193 34897 36196
rect 34931 36193 34943 36227
rect 34885 36187 34943 36193
rect 32582 36156 32588 36168
rect 31343 36128 31754 36156
rect 32543 36128 32588 36156
rect 31343 36125 31355 36128
rect 31297 36119 31355 36125
rect 32582 36116 32588 36128
rect 32640 36116 32646 36168
rect 32769 36159 32827 36165
rect 32769 36125 32781 36159
rect 32815 36156 32827 36159
rect 33413 36159 33471 36165
rect 33413 36156 33425 36159
rect 32815 36128 33425 36156
rect 32815 36125 32827 36128
rect 32769 36119 32827 36125
rect 33413 36125 33425 36128
rect 33459 36156 33471 36159
rect 33778 36156 33784 36168
rect 33459 36128 33784 36156
rect 33459 36125 33471 36128
rect 33413 36119 33471 36125
rect 33778 36116 33784 36128
rect 33836 36116 33842 36168
rect 34900 36156 34928 36187
rect 36262 36156 36268 36168
rect 34900 36128 36268 36156
rect 36262 36116 36268 36128
rect 36320 36156 36326 36168
rect 36817 36159 36875 36165
rect 36817 36156 36829 36159
rect 36320 36128 36829 36156
rect 36320 36116 36326 36128
rect 36817 36125 36829 36128
rect 36863 36125 36875 36159
rect 36817 36119 36875 36125
rect 27580 36060 28488 36088
rect 28537 36091 28595 36097
rect 27580 36048 27586 36060
rect 28537 36057 28549 36091
rect 28583 36088 28595 36091
rect 29270 36088 29276 36100
rect 28583 36060 29276 36088
rect 28583 36057 28595 36060
rect 28537 36051 28595 36057
rect 29270 36048 29276 36060
rect 29328 36048 29334 36100
rect 32600 36088 32628 36116
rect 33229 36091 33287 36097
rect 33229 36088 33241 36091
rect 32600 36060 33241 36088
rect 33229 36057 33241 36060
rect 33275 36057 33287 36091
rect 33229 36051 33287 36057
rect 34514 36048 34520 36100
rect 34572 36088 34578 36100
rect 35130 36091 35188 36097
rect 35130 36088 35142 36091
rect 34572 36060 35142 36088
rect 34572 36048 34578 36060
rect 35130 36057 35142 36060
rect 35176 36057 35188 36091
rect 35130 36051 35188 36057
rect 37084 36091 37142 36097
rect 37084 36057 37096 36091
rect 37130 36088 37142 36091
rect 37458 36088 37464 36100
rect 37130 36060 37464 36088
rect 37130 36057 37142 36060
rect 37084 36051 37142 36057
rect 37458 36048 37464 36060
rect 37516 36048 37522 36100
rect 16114 36020 16120 36032
rect 12406 35992 16120 36020
rect 16114 35980 16120 35992
rect 16172 35980 16178 36032
rect 17635 36023 17693 36029
rect 17635 35989 17647 36023
rect 17681 36020 17693 36023
rect 18782 36020 18788 36032
rect 17681 35992 18788 36020
rect 17681 35989 17693 35992
rect 17635 35983 17693 35989
rect 18782 35980 18788 35992
rect 18840 35980 18846 36032
rect 22462 35980 22468 36032
rect 22520 36020 22526 36032
rect 25501 36023 25559 36029
rect 22520 35992 22565 36020
rect 22520 35980 22526 35992
rect 25501 35989 25513 36023
rect 25547 36020 25559 36023
rect 26786 36020 26792 36032
rect 25547 35992 26792 36020
rect 25547 35989 25559 35992
rect 25501 35983 25559 35989
rect 26786 35980 26792 35992
rect 26844 35980 26850 36032
rect 29086 35980 29092 36032
rect 29144 36020 29150 36032
rect 30285 36023 30343 36029
rect 30285 36020 30297 36023
rect 29144 35992 30297 36020
rect 29144 35980 29150 35992
rect 30285 35989 30297 35992
rect 30331 35989 30343 36023
rect 30285 35983 30343 35989
rect 36078 35980 36084 36032
rect 36136 36020 36142 36032
rect 36265 36023 36323 36029
rect 36265 36020 36277 36023
rect 36136 35992 36277 36020
rect 36136 35980 36142 35992
rect 36265 35989 36277 35992
rect 36311 35989 36323 36023
rect 36265 35983 36323 35989
rect 37826 35980 37832 36032
rect 37884 36020 37890 36032
rect 38197 36023 38255 36029
rect 38197 36020 38209 36023
rect 37884 35992 38209 36020
rect 37884 35980 37890 35992
rect 38197 35989 38209 35992
rect 38243 35989 38255 36023
rect 38197 35983 38255 35989
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 7098 35816 7104 35828
rect 7059 35788 7104 35816
rect 7098 35776 7104 35788
rect 7156 35776 7162 35828
rect 7561 35819 7619 35825
rect 7561 35785 7573 35819
rect 7607 35816 7619 35819
rect 7742 35816 7748 35828
rect 7607 35788 7748 35816
rect 7607 35785 7619 35788
rect 7561 35779 7619 35785
rect 7742 35776 7748 35788
rect 7800 35776 7806 35828
rect 11698 35816 11704 35828
rect 11659 35788 11704 35816
rect 11698 35776 11704 35788
rect 11756 35776 11762 35828
rect 11882 35776 11888 35828
rect 11940 35816 11946 35828
rect 12161 35819 12219 35825
rect 12161 35816 12173 35819
rect 11940 35788 12173 35816
rect 11940 35776 11946 35788
rect 12161 35785 12173 35788
rect 12207 35785 12219 35819
rect 12161 35779 12219 35785
rect 13262 35776 13268 35828
rect 13320 35816 13326 35828
rect 22005 35819 22063 35825
rect 13320 35788 20576 35816
rect 13320 35776 13326 35788
rect 7469 35751 7527 35757
rect 7469 35717 7481 35751
rect 7515 35748 7527 35751
rect 8294 35748 8300 35760
rect 7515 35720 8300 35748
rect 7515 35717 7527 35720
rect 7469 35711 7527 35717
rect 8294 35708 8300 35720
rect 8352 35748 8358 35760
rect 9306 35748 9312 35760
rect 8352 35720 9312 35748
rect 8352 35708 8358 35720
rect 9306 35708 9312 35720
rect 9364 35708 9370 35760
rect 19996 35720 20300 35748
rect 9950 35680 9956 35692
rect 9911 35652 9956 35680
rect 9950 35640 9956 35652
rect 10008 35640 10014 35692
rect 11606 35640 11612 35692
rect 11664 35680 11670 35692
rect 12069 35683 12127 35689
rect 12069 35680 12081 35683
rect 11664 35652 12081 35680
rect 11664 35640 11670 35652
rect 12069 35649 12081 35652
rect 12115 35680 12127 35683
rect 12158 35680 12164 35692
rect 12115 35652 12164 35680
rect 12115 35649 12127 35652
rect 12069 35643 12127 35649
rect 12158 35640 12164 35652
rect 12216 35640 12222 35692
rect 13354 35680 13360 35692
rect 13315 35652 13360 35680
rect 13354 35640 13360 35652
rect 13412 35640 13418 35692
rect 14734 35640 14740 35692
rect 14792 35640 14798 35692
rect 16482 35640 16488 35692
rect 16540 35680 16546 35692
rect 16853 35683 16911 35689
rect 16853 35680 16865 35683
rect 16540 35652 16865 35680
rect 16540 35640 16546 35652
rect 16853 35649 16865 35652
rect 16899 35649 16911 35683
rect 17678 35680 17684 35692
rect 17639 35652 17684 35680
rect 16853 35643 16911 35649
rect 17678 35640 17684 35652
rect 17736 35640 17742 35692
rect 18782 35680 18788 35692
rect 18743 35652 18788 35680
rect 18782 35640 18788 35652
rect 18840 35640 18846 35692
rect 19797 35683 19855 35689
rect 19797 35649 19809 35683
rect 19843 35680 19855 35683
rect 19886 35680 19892 35692
rect 19843 35652 19892 35680
rect 19843 35649 19855 35652
rect 19797 35643 19855 35649
rect 19886 35640 19892 35652
rect 19944 35640 19950 35692
rect 19996 35689 20024 35720
rect 19981 35683 20039 35689
rect 19981 35649 19993 35683
rect 20027 35649 20039 35683
rect 19981 35643 20039 35649
rect 7650 35612 7656 35624
rect 7611 35584 7656 35612
rect 7650 35572 7656 35584
rect 7708 35572 7714 35624
rect 10042 35612 10048 35624
rect 10003 35584 10048 35612
rect 10042 35572 10048 35584
rect 10100 35572 10106 35624
rect 10137 35615 10195 35621
rect 10137 35581 10149 35615
rect 10183 35612 10195 35615
rect 12253 35615 12311 35621
rect 12253 35612 12265 35615
rect 10183 35584 12265 35612
rect 10183 35581 10195 35584
rect 10137 35575 10195 35581
rect 12253 35581 12265 35584
rect 12299 35612 12311 35615
rect 13630 35612 13636 35624
rect 12299 35584 12434 35612
rect 13591 35584 13636 35612
rect 12299 35581 12311 35584
rect 12253 35575 12311 35581
rect 7668 35544 7696 35572
rect 9398 35544 9404 35556
rect 7668 35516 9404 35544
rect 9398 35504 9404 35516
rect 9456 35544 9462 35556
rect 10152 35544 10180 35575
rect 9456 35516 10180 35544
rect 12406 35544 12434 35584
rect 13630 35572 13636 35584
rect 13688 35572 13694 35624
rect 17954 35612 17960 35624
rect 17915 35584 17960 35612
rect 17954 35572 17960 35584
rect 18012 35572 18018 35624
rect 19061 35615 19119 35621
rect 19061 35581 19073 35615
rect 19107 35612 19119 35615
rect 19150 35612 19156 35624
rect 19107 35584 19156 35612
rect 19107 35581 19119 35584
rect 19061 35575 19119 35581
rect 19150 35572 19156 35584
rect 19208 35572 19214 35624
rect 13262 35544 13268 35556
rect 12406 35516 13268 35544
rect 9456 35504 9462 35516
rect 13262 35504 13268 35516
rect 13320 35504 13326 35556
rect 18414 35504 18420 35556
rect 18472 35544 18478 35556
rect 19702 35544 19708 35556
rect 18472 35516 19708 35544
rect 18472 35504 18478 35516
rect 19702 35504 19708 35516
rect 19760 35504 19766 35556
rect 19904 35544 19932 35640
rect 20272 35612 20300 35720
rect 20438 35680 20444 35692
rect 20399 35652 20444 35680
rect 20438 35640 20444 35652
rect 20496 35640 20502 35692
rect 20548 35680 20576 35788
rect 22005 35785 22017 35819
rect 22051 35816 22063 35819
rect 22094 35816 22100 35828
rect 22051 35788 22100 35816
rect 22051 35785 22063 35788
rect 22005 35779 22063 35785
rect 22094 35776 22100 35788
rect 22152 35776 22158 35828
rect 22465 35819 22523 35825
rect 22465 35785 22477 35819
rect 22511 35816 22523 35819
rect 22922 35816 22928 35828
rect 22511 35788 22928 35816
rect 22511 35785 22523 35788
rect 22465 35779 22523 35785
rect 22922 35776 22928 35788
rect 22980 35776 22986 35828
rect 23198 35776 23204 35828
rect 23256 35816 23262 35828
rect 26513 35819 26571 35825
rect 26513 35816 26525 35819
rect 23256 35788 26525 35816
rect 23256 35776 23262 35788
rect 26513 35785 26525 35788
rect 26559 35785 26571 35819
rect 26513 35779 26571 35785
rect 33689 35819 33747 35825
rect 33689 35785 33701 35819
rect 33735 35816 33747 35819
rect 34514 35816 34520 35828
rect 33735 35788 34520 35816
rect 33735 35785 33747 35788
rect 33689 35779 33747 35785
rect 34514 35776 34520 35788
rect 34572 35776 34578 35828
rect 36446 35776 36452 35828
rect 36504 35816 36510 35828
rect 36817 35819 36875 35825
rect 36817 35816 36829 35819
rect 36504 35788 36829 35816
rect 36504 35776 36510 35788
rect 36817 35785 36829 35788
rect 36863 35785 36875 35819
rect 37458 35816 37464 35828
rect 37419 35788 37464 35816
rect 36817 35779 36875 35785
rect 37458 35776 37464 35788
rect 37516 35776 37522 35828
rect 20622 35708 20628 35760
rect 20680 35748 20686 35760
rect 26329 35751 26387 35757
rect 26329 35748 26341 35751
rect 20680 35720 26341 35748
rect 20680 35708 20686 35720
rect 22373 35683 22431 35689
rect 20548 35652 22094 35680
rect 20717 35615 20775 35621
rect 20717 35612 20729 35615
rect 20272 35584 20729 35612
rect 20717 35581 20729 35584
rect 20763 35612 20775 35615
rect 21358 35612 21364 35624
rect 20763 35584 21364 35612
rect 20763 35581 20775 35584
rect 20717 35575 20775 35581
rect 21358 35572 21364 35584
rect 21416 35572 21422 35624
rect 22066 35544 22094 35652
rect 22373 35649 22385 35683
rect 22419 35680 22431 35683
rect 22462 35680 22468 35692
rect 22419 35652 22468 35680
rect 22419 35649 22431 35652
rect 22373 35643 22431 35649
rect 22462 35640 22468 35652
rect 22520 35640 22526 35692
rect 22922 35640 22928 35692
rect 22980 35680 22986 35692
rect 23198 35680 23204 35692
rect 22980 35652 23204 35680
rect 22980 35640 22986 35652
rect 23198 35640 23204 35652
rect 23256 35640 23262 35692
rect 23400 35689 23428 35720
rect 26329 35717 26341 35720
rect 26375 35748 26387 35751
rect 26418 35748 26424 35760
rect 26375 35720 26424 35748
rect 26375 35717 26387 35720
rect 26329 35711 26387 35717
rect 26418 35708 26424 35720
rect 26476 35708 26482 35760
rect 32030 35708 32036 35760
rect 32088 35748 32094 35760
rect 35618 35748 35624 35760
rect 32088 35720 35624 35748
rect 32088 35708 32094 35720
rect 35618 35708 35624 35720
rect 35676 35708 35682 35760
rect 23385 35683 23443 35689
rect 23385 35649 23397 35683
rect 23431 35649 23443 35683
rect 24946 35680 24952 35692
rect 24907 35652 24952 35680
rect 23385 35643 23443 35649
rect 24946 35640 24952 35652
rect 25004 35640 25010 35692
rect 26510 35640 26516 35692
rect 26568 35680 26574 35692
rect 26605 35683 26663 35689
rect 26605 35680 26617 35683
rect 26568 35652 26617 35680
rect 26568 35640 26574 35652
rect 26605 35649 26617 35652
rect 26651 35649 26663 35683
rect 27246 35680 27252 35692
rect 27207 35652 27252 35680
rect 26605 35643 26663 35649
rect 27246 35640 27252 35652
rect 27304 35640 27310 35692
rect 28626 35680 28632 35692
rect 28587 35652 28632 35680
rect 28626 35640 28632 35652
rect 28684 35640 28690 35692
rect 28902 35689 28908 35692
rect 28896 35643 28908 35689
rect 28960 35680 28966 35692
rect 28960 35652 28996 35680
rect 28902 35640 28908 35643
rect 28960 35640 28966 35652
rect 32674 35640 32680 35692
rect 32732 35680 32738 35692
rect 32769 35683 32827 35689
rect 32769 35680 32781 35683
rect 32732 35652 32781 35680
rect 32732 35640 32738 35652
rect 32769 35649 32781 35652
rect 32815 35649 32827 35683
rect 32950 35680 32956 35692
rect 32911 35652 32956 35680
rect 32769 35643 32827 35649
rect 32950 35640 32956 35652
rect 33008 35640 33014 35692
rect 33042 35640 33048 35692
rect 33100 35680 33106 35692
rect 33597 35683 33655 35689
rect 33100 35652 33145 35680
rect 33100 35640 33106 35652
rect 33597 35649 33609 35683
rect 33643 35649 33655 35683
rect 33778 35680 33784 35692
rect 33739 35652 33784 35680
rect 33597 35643 33655 35649
rect 22649 35615 22707 35621
rect 22649 35581 22661 35615
rect 22695 35612 22707 35615
rect 23661 35615 23719 35621
rect 23661 35612 23673 35615
rect 22695 35584 23673 35612
rect 22695 35581 22707 35584
rect 22649 35575 22707 35581
rect 23661 35581 23673 35584
rect 23707 35581 23719 35615
rect 24854 35612 24860 35624
rect 24815 35584 24860 35612
rect 23661 35575 23719 35581
rect 22664 35544 22692 35575
rect 24854 35572 24860 35584
rect 24912 35572 24918 35624
rect 25406 35612 25412 35624
rect 25367 35584 25412 35612
rect 25406 35572 25412 35584
rect 25464 35572 25470 35624
rect 26234 35612 26240 35624
rect 25992 35584 26240 35612
rect 25992 35544 26020 35584
rect 26234 35572 26240 35584
rect 26292 35612 26298 35624
rect 27522 35612 27528 35624
rect 26292 35584 27528 35612
rect 26292 35572 26298 35584
rect 27522 35572 27528 35584
rect 27580 35612 27586 35624
rect 27798 35612 27804 35624
rect 27580 35584 27804 35612
rect 27580 35572 27586 35584
rect 27798 35572 27804 35584
rect 27856 35572 27862 35624
rect 33612 35612 33640 35643
rect 33778 35640 33784 35652
rect 33836 35640 33842 35692
rect 35986 35640 35992 35692
rect 36044 35680 36050 35692
rect 36725 35683 36783 35689
rect 36725 35680 36737 35683
rect 36044 35652 36737 35680
rect 36044 35640 36050 35652
rect 36725 35649 36737 35652
rect 36771 35649 36783 35683
rect 37826 35680 37832 35692
rect 37787 35652 37832 35680
rect 36725 35643 36783 35649
rect 37826 35640 37832 35652
rect 37884 35640 37890 35692
rect 32784 35584 33640 35612
rect 26326 35544 26332 35556
rect 19904 35516 20208 35544
rect 22066 35516 22692 35544
rect 23584 35516 26020 35544
rect 26287 35516 26332 35544
rect 20180 35488 20208 35516
rect 9582 35476 9588 35488
rect 9543 35448 9588 35476
rect 9582 35436 9588 35448
rect 9640 35436 9646 35488
rect 14826 35436 14832 35488
rect 14884 35476 14890 35488
rect 15105 35479 15163 35485
rect 15105 35476 15117 35479
rect 14884 35448 15117 35476
rect 14884 35436 14890 35448
rect 15105 35445 15117 35448
rect 15151 35476 15163 35479
rect 16574 35476 16580 35488
rect 15151 35448 16580 35476
rect 15151 35445 15163 35448
rect 15105 35439 15163 35445
rect 16574 35436 16580 35448
rect 16632 35436 16638 35488
rect 16942 35476 16948 35488
rect 16903 35448 16948 35476
rect 16942 35436 16948 35448
rect 17000 35436 17006 35488
rect 19797 35479 19855 35485
rect 19797 35445 19809 35479
rect 19843 35476 19855 35479
rect 19886 35476 19892 35488
rect 19843 35448 19892 35476
rect 19843 35445 19855 35448
rect 19797 35439 19855 35445
rect 19886 35436 19892 35448
rect 19944 35436 19950 35488
rect 20162 35436 20168 35488
rect 20220 35436 20226 35488
rect 20530 35436 20536 35488
rect 20588 35476 20594 35488
rect 23584 35476 23612 35516
rect 26326 35504 26332 35516
rect 26384 35504 26390 35556
rect 32784 35553 32812 35584
rect 37734 35572 37740 35624
rect 37792 35612 37798 35624
rect 37921 35615 37979 35621
rect 37921 35612 37933 35615
rect 37792 35584 37933 35612
rect 37792 35572 37798 35584
rect 37921 35581 37933 35584
rect 37967 35581 37979 35615
rect 37921 35575 37979 35581
rect 38010 35572 38016 35624
rect 38068 35612 38074 35624
rect 38068 35584 38113 35612
rect 38068 35572 38074 35584
rect 32769 35547 32827 35553
rect 32769 35513 32781 35547
rect 32815 35513 32827 35547
rect 32769 35507 32827 35513
rect 20588 35448 23612 35476
rect 20588 35436 20594 35448
rect 23658 35436 23664 35488
rect 23716 35476 23722 35488
rect 24670 35476 24676 35488
rect 23716 35448 24676 35476
rect 23716 35436 23722 35448
rect 24670 35436 24676 35448
rect 24728 35476 24734 35488
rect 25317 35479 25375 35485
rect 25317 35476 25329 35479
rect 24728 35448 25329 35476
rect 24728 35436 24734 35448
rect 25317 35445 25329 35448
rect 25363 35445 25375 35479
rect 25317 35439 25375 35445
rect 25685 35479 25743 35485
rect 25685 35445 25697 35479
rect 25731 35476 25743 35479
rect 26418 35476 26424 35488
rect 25731 35448 26424 35476
rect 25731 35445 25743 35448
rect 25685 35439 25743 35445
rect 26418 35436 26424 35448
rect 26476 35436 26482 35488
rect 28534 35436 28540 35488
rect 28592 35476 28598 35488
rect 30006 35476 30012 35488
rect 28592 35448 30012 35476
rect 28592 35436 28598 35448
rect 30006 35436 30012 35448
rect 30064 35436 30070 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 10042 35232 10048 35284
rect 10100 35272 10106 35284
rect 10505 35275 10563 35281
rect 10505 35272 10517 35275
rect 10100 35244 10517 35272
rect 10100 35232 10106 35244
rect 10505 35241 10517 35244
rect 10551 35241 10563 35275
rect 10505 35235 10563 35241
rect 14734 35232 14740 35284
rect 14792 35272 14798 35284
rect 14829 35275 14887 35281
rect 14829 35272 14841 35275
rect 14792 35244 14841 35272
rect 14792 35232 14798 35244
rect 14829 35241 14841 35244
rect 14875 35241 14887 35275
rect 14829 35235 14887 35241
rect 17129 35275 17187 35281
rect 17129 35241 17141 35275
rect 17175 35272 17187 35275
rect 18414 35272 18420 35284
rect 17175 35244 18420 35272
rect 17175 35241 17187 35244
rect 17129 35235 17187 35241
rect 18414 35232 18420 35244
rect 18472 35232 18478 35284
rect 19978 35232 19984 35284
rect 20036 35272 20042 35284
rect 20901 35275 20959 35281
rect 20901 35272 20913 35275
rect 20036 35244 20913 35272
rect 20036 35232 20042 35244
rect 20901 35241 20913 35244
rect 20947 35241 20959 35275
rect 23566 35272 23572 35284
rect 23479 35244 23572 35272
rect 20901 35235 20959 35241
rect 23566 35232 23572 35244
rect 23624 35272 23630 35284
rect 24854 35272 24860 35284
rect 23624 35244 24860 35272
rect 23624 35232 23630 35244
rect 24854 35232 24860 35244
rect 24912 35232 24918 35284
rect 28902 35232 28908 35284
rect 28960 35272 28966 35284
rect 28997 35275 29055 35281
rect 28997 35272 29009 35275
rect 28960 35244 29009 35272
rect 28960 35232 28966 35244
rect 28997 35241 29009 35244
rect 29043 35241 29055 35275
rect 28997 35235 29055 35241
rect 31202 35232 31208 35284
rect 31260 35272 31266 35284
rect 31297 35275 31355 35281
rect 31297 35272 31309 35275
rect 31260 35244 31309 35272
rect 31260 35232 31266 35244
rect 31297 35241 31309 35244
rect 31343 35241 31355 35275
rect 31297 35235 31355 35241
rect 32401 35275 32459 35281
rect 32401 35241 32413 35275
rect 32447 35272 32459 35275
rect 32582 35272 32588 35284
rect 32447 35244 32588 35272
rect 32447 35241 32459 35244
rect 32401 35235 32459 35241
rect 32582 35232 32588 35244
rect 32640 35232 32646 35284
rect 32858 35232 32864 35284
rect 32916 35272 32922 35284
rect 33042 35272 33048 35284
rect 32916 35244 33048 35272
rect 32916 35232 32922 35244
rect 33042 35232 33048 35244
rect 33100 35232 33106 35284
rect 33229 35275 33287 35281
rect 33229 35241 33241 35275
rect 33275 35272 33287 35275
rect 33778 35272 33784 35284
rect 33275 35244 33784 35272
rect 33275 35241 33287 35244
rect 33229 35235 33287 35241
rect 33778 35232 33784 35244
rect 33836 35232 33842 35284
rect 11330 35204 11336 35216
rect 11291 35176 11336 35204
rect 11330 35164 11336 35176
rect 11388 35164 11394 35216
rect 11882 35164 11888 35216
rect 11940 35204 11946 35216
rect 18877 35207 18935 35213
rect 11940 35176 13216 35204
rect 11940 35164 11946 35176
rect 5721 35139 5779 35145
rect 5721 35105 5733 35139
rect 5767 35136 5779 35139
rect 7650 35136 7656 35148
rect 5767 35108 7656 35136
rect 5767 35105 5779 35108
rect 5721 35099 5779 35105
rect 7650 35096 7656 35108
rect 7708 35096 7714 35148
rect 12710 35136 12716 35148
rect 12671 35108 12716 35136
rect 12710 35096 12716 35108
rect 12768 35096 12774 35148
rect 13078 35136 13084 35148
rect 12820 35108 13084 35136
rect 9125 35071 9183 35077
rect 9125 35037 9137 35071
rect 9171 35068 9183 35071
rect 9674 35068 9680 35080
rect 9171 35040 9680 35068
rect 9171 35037 9183 35040
rect 9125 35031 9183 35037
rect 9674 35028 9680 35040
rect 9732 35028 9738 35080
rect 12820 35077 12848 35108
rect 13078 35096 13084 35108
rect 13136 35096 13142 35148
rect 12805 35071 12863 35077
rect 12805 35037 12817 35071
rect 12851 35037 12863 35071
rect 12805 35031 12863 35037
rect 12989 35071 13047 35077
rect 12989 35037 13001 35071
rect 13035 35068 13047 35071
rect 13188 35068 13216 35176
rect 18877 35173 18889 35207
rect 18923 35204 18935 35207
rect 19334 35204 19340 35216
rect 18923 35176 19340 35204
rect 18923 35173 18935 35176
rect 18877 35167 18935 35173
rect 19334 35164 19340 35176
rect 19392 35204 19398 35216
rect 19392 35176 20300 35204
rect 19392 35164 19398 35176
rect 15381 35139 15439 35145
rect 15381 35105 15393 35139
rect 15427 35136 15439 35139
rect 15746 35136 15752 35148
rect 15427 35108 15752 35136
rect 15427 35105 15439 35108
rect 15381 35099 15439 35105
rect 15746 35096 15752 35108
rect 15804 35096 15810 35148
rect 19886 35096 19892 35148
rect 19944 35096 19950 35148
rect 20272 35145 20300 35176
rect 31662 35164 31668 35216
rect 31720 35204 31726 35216
rect 31720 35176 32260 35204
rect 31720 35164 31726 35176
rect 20257 35139 20315 35145
rect 20257 35105 20269 35139
rect 20303 35105 20315 35139
rect 20257 35099 20315 35105
rect 22373 35139 22431 35145
rect 22373 35105 22385 35139
rect 22419 35136 22431 35139
rect 23566 35136 23572 35148
rect 22419 35108 23572 35136
rect 22419 35105 22431 35108
rect 22373 35099 22431 35105
rect 23566 35096 23572 35108
rect 23624 35096 23630 35148
rect 23661 35139 23719 35145
rect 23661 35105 23673 35139
rect 23707 35136 23719 35139
rect 23842 35136 23848 35148
rect 23707 35108 23848 35136
rect 23707 35105 23719 35108
rect 23661 35099 23719 35105
rect 23842 35096 23848 35108
rect 23900 35096 23906 35148
rect 29086 35136 29092 35148
rect 29047 35108 29092 35136
rect 29086 35096 29092 35108
rect 29144 35096 29150 35148
rect 32122 35136 32128 35148
rect 31036 35108 32128 35136
rect 13538 35068 13544 35080
rect 13035 35040 13544 35068
rect 13035 35037 13047 35040
rect 12989 35031 13047 35037
rect 13538 35028 13544 35040
rect 13596 35028 13602 35080
rect 14737 35071 14795 35077
rect 14737 35037 14749 35071
rect 14783 35068 14795 35071
rect 15194 35068 15200 35080
rect 14783 35040 15200 35068
rect 14783 35037 14795 35040
rect 14737 35031 14795 35037
rect 15194 35028 15200 35040
rect 15252 35028 15258 35080
rect 18230 35068 18236 35080
rect 18191 35040 18236 35068
rect 18230 35028 18236 35040
rect 18288 35028 18294 35080
rect 19794 35068 19800 35080
rect 19755 35040 19800 35068
rect 19794 35028 19800 35040
rect 19852 35028 19858 35080
rect 19904 35068 19932 35096
rect 31036 35080 31064 35108
rect 32122 35096 32128 35108
rect 32180 35096 32186 35148
rect 20099 35071 20157 35077
rect 20099 35068 20111 35071
rect 19904 35040 20111 35068
rect 20099 35037 20111 35040
rect 20145 35068 20157 35071
rect 20145 35040 20300 35068
rect 20145 35037 20157 35040
rect 20099 35031 20157 35037
rect 5445 35003 5503 35009
rect 5445 34969 5457 35003
rect 5491 35000 5503 35003
rect 5718 35000 5724 35012
rect 5491 34972 5724 35000
rect 5491 34969 5503 34972
rect 5445 34963 5503 34969
rect 5718 34960 5724 34972
rect 5776 34960 5782 35012
rect 9392 35003 9450 35009
rect 9392 34969 9404 35003
rect 9438 35000 9450 35003
rect 9582 35000 9588 35012
rect 9438 34972 9588 35000
rect 9438 34969 9450 34972
rect 9392 34963 9450 34969
rect 9582 34960 9588 34972
rect 9640 34960 9646 35012
rect 11606 35000 11612 35012
rect 11567 34972 11612 35000
rect 11606 34960 11612 34972
rect 11664 34960 11670 35012
rect 11790 35000 11796 35012
rect 11751 34972 11796 35000
rect 11790 34960 11796 34972
rect 11848 34960 11854 35012
rect 11882 34960 11888 35012
rect 11940 35000 11946 35012
rect 13449 35003 13507 35009
rect 13449 35000 13461 35003
rect 11940 34972 11985 35000
rect 12728 34972 13461 35000
rect 11940 34960 11946 34972
rect 12728 34944 12756 34972
rect 13449 34969 13461 34972
rect 13495 34969 13507 35003
rect 13449 34963 13507 34969
rect 15657 35003 15715 35009
rect 15657 34969 15669 35003
rect 15703 35000 15715 35003
rect 15930 35000 15936 35012
rect 15703 34972 15936 35000
rect 15703 34969 15715 34972
rect 15657 34963 15715 34969
rect 15930 34960 15936 34972
rect 15988 34960 15994 35012
rect 16942 35000 16948 35012
rect 16882 34972 16948 35000
rect 16942 34960 16948 34972
rect 17000 34960 17006 35012
rect 18414 34960 18420 35012
rect 18472 35000 18478 35012
rect 18601 35003 18659 35009
rect 18601 35000 18613 35003
rect 18472 34972 18613 35000
rect 18472 34960 18478 34972
rect 18601 34969 18613 34972
rect 18647 34969 18659 35003
rect 18601 34963 18659 34969
rect 18718 35003 18776 35009
rect 18718 34969 18730 35003
rect 18764 35000 18776 35003
rect 19058 35000 19064 35012
rect 18764 34972 19064 35000
rect 18764 34969 18776 34972
rect 18718 34963 18776 34969
rect 19058 34960 19064 34972
rect 19116 34960 19122 35012
rect 19889 35003 19947 35009
rect 19889 34969 19901 35003
rect 19935 34969 19947 35003
rect 19889 34963 19947 34969
rect 5074 34932 5080 34944
rect 5035 34904 5080 34932
rect 5074 34892 5080 34904
rect 5132 34892 5138 34944
rect 5534 34892 5540 34944
rect 5592 34932 5598 34944
rect 5592 34904 5637 34932
rect 5592 34892 5598 34904
rect 12710 34892 12716 34944
rect 12768 34892 12774 34944
rect 18509 34935 18567 34941
rect 18509 34901 18521 34935
rect 18555 34932 18567 34935
rect 19150 34932 19156 34944
rect 18555 34904 19156 34932
rect 18555 34901 18567 34904
rect 18509 34895 18567 34901
rect 19150 34892 19156 34904
rect 19208 34892 19214 34944
rect 19426 34892 19432 34944
rect 19484 34932 19490 34944
rect 19613 34935 19671 34941
rect 19613 34932 19625 34935
rect 19484 34904 19625 34932
rect 19484 34892 19490 34904
rect 19613 34901 19625 34904
rect 19659 34901 19671 34935
rect 19904 34932 19932 34963
rect 19978 34960 19984 35012
rect 20036 35000 20042 35012
rect 20272 35000 20300 35040
rect 20898 35028 20904 35080
rect 20956 35068 20962 35080
rect 22002 35068 22008 35080
rect 20956 35040 22008 35068
rect 20956 35028 20962 35040
rect 22002 35028 22008 35040
rect 22060 35068 22066 35080
rect 22097 35071 22155 35077
rect 22097 35068 22109 35071
rect 22060 35040 22109 35068
rect 22060 35028 22066 35040
rect 22097 35037 22109 35040
rect 22143 35037 22155 35071
rect 22097 35031 22155 35037
rect 23109 35071 23167 35077
rect 23109 35037 23121 35071
rect 23155 35037 23167 35071
rect 23109 35031 23167 35037
rect 20717 35003 20775 35009
rect 20717 35000 20729 35003
rect 20036 34972 20081 35000
rect 20272 34972 20729 35000
rect 20036 34960 20042 34972
rect 20717 34969 20729 34972
rect 20763 34969 20775 35003
rect 23124 35000 23152 35031
rect 23198 35028 23204 35080
rect 23256 35068 23262 35080
rect 24946 35068 24952 35080
rect 23256 35040 24952 35068
rect 23256 35028 23262 35040
rect 24946 35028 24952 35040
rect 25004 35028 25010 35080
rect 27154 35028 27160 35080
rect 27212 35068 27218 35080
rect 27341 35071 27399 35077
rect 27341 35068 27353 35071
rect 27212 35040 27353 35068
rect 27212 35028 27218 35040
rect 27341 35037 27353 35040
rect 27387 35037 27399 35071
rect 27341 35031 27399 35037
rect 27430 35028 27436 35080
rect 27488 35068 27494 35080
rect 28813 35071 28871 35077
rect 27488 35040 27533 35068
rect 27488 35028 27494 35040
rect 28813 35037 28825 35071
rect 28859 35037 28871 35071
rect 28813 35031 28871 35037
rect 23658 35000 23664 35012
rect 23124 34972 23664 35000
rect 20717 34963 20775 34969
rect 23658 34960 23664 34972
rect 23716 34960 23722 35012
rect 25130 35000 25136 35012
rect 25091 34972 25136 35000
rect 25130 34960 25136 34972
rect 25188 34960 25194 35012
rect 28828 35000 28856 35031
rect 28902 35028 28908 35080
rect 28960 35068 28966 35080
rect 30650 35068 30656 35080
rect 28960 35040 29005 35068
rect 30611 35040 30656 35068
rect 28960 35028 28966 35040
rect 30650 35028 30656 35040
rect 30708 35028 30714 35080
rect 30742 35028 30748 35080
rect 30800 35068 30806 35080
rect 31018 35068 31024 35080
rect 30800 35040 30845 35068
rect 30979 35040 31024 35068
rect 30800 35028 30806 35040
rect 31018 35028 31024 35040
rect 31076 35028 31082 35080
rect 31159 35071 31217 35077
rect 31159 35037 31171 35071
rect 31205 35068 31217 35071
rect 31662 35068 31668 35080
rect 31205 35040 31668 35068
rect 31205 35037 31217 35040
rect 31159 35031 31217 35037
rect 31662 35028 31668 35040
rect 31720 35028 31726 35080
rect 31754 35028 31760 35080
rect 31812 35068 31818 35080
rect 31938 35077 31944 35080
rect 31905 35071 31944 35077
rect 31812 35040 31857 35068
rect 31812 35028 31818 35040
rect 31905 35037 31917 35071
rect 31905 35031 31944 35037
rect 31938 35028 31944 35031
rect 31996 35028 32002 35080
rect 32232 35077 32260 35176
rect 36262 35136 36268 35148
rect 36223 35108 36268 35136
rect 36262 35096 36268 35108
rect 36320 35096 36326 35148
rect 32222 35071 32280 35077
rect 32222 35037 32234 35071
rect 32268 35037 32280 35071
rect 34698 35068 34704 35080
rect 32222 35031 32280 35037
rect 32600 35040 34704 35068
rect 29178 35000 29184 35012
rect 28828 34972 29184 35000
rect 29178 34960 29184 34972
rect 29236 34960 29242 35012
rect 30929 35003 30987 35009
rect 30929 34969 30941 35003
rect 30975 35000 30987 35003
rect 32033 35003 32091 35009
rect 32033 35000 32045 35003
rect 30975 34972 32045 35000
rect 30975 34969 30987 34972
rect 30929 34963 30987 34969
rect 31128 34944 31156 34972
rect 32033 34969 32045 34972
rect 32079 34969 32091 35003
rect 32033 34963 32091 34969
rect 32125 35003 32183 35009
rect 32125 34969 32137 35003
rect 32171 35000 32183 35003
rect 32306 35000 32312 35012
rect 32171 34972 32312 35000
rect 32171 34969 32183 34972
rect 32125 34963 32183 34969
rect 32306 34960 32312 34972
rect 32364 35000 32370 35012
rect 32600 35000 32628 35040
rect 34698 35028 34704 35040
rect 34756 35028 34762 35080
rect 32364 34972 32628 35000
rect 32861 35003 32919 35009
rect 32364 34960 32370 34972
rect 32861 34969 32873 35003
rect 32907 35000 32919 35003
rect 32950 35000 32956 35012
rect 32907 34972 32956 35000
rect 32907 34969 32919 34972
rect 32861 34963 32919 34969
rect 32950 34960 32956 34972
rect 33008 34960 33014 35012
rect 36170 34960 36176 35012
rect 36228 35000 36234 35012
rect 36510 35003 36568 35009
rect 36510 35000 36522 35003
rect 36228 34972 36522 35000
rect 36228 34960 36234 34972
rect 36510 34969 36522 34972
rect 36556 34969 36568 35003
rect 36510 34963 36568 34969
rect 20438 34932 20444 34944
rect 19904 34904 20444 34932
rect 19613 34895 19671 34901
rect 20438 34892 20444 34904
rect 20496 34932 20502 34944
rect 20901 34935 20959 34941
rect 20901 34932 20913 34935
rect 20496 34904 20913 34932
rect 20496 34892 20502 34904
rect 20901 34901 20913 34904
rect 20947 34901 20959 34935
rect 21082 34932 21088 34944
rect 21043 34904 21088 34932
rect 20901 34895 20959 34901
rect 21082 34892 21088 34904
rect 21140 34892 21146 34944
rect 22738 34892 22744 34944
rect 22796 34932 22802 34944
rect 23937 34935 23995 34941
rect 23937 34932 23949 34935
rect 22796 34904 23949 34932
rect 22796 34892 22802 34904
rect 23937 34901 23949 34904
rect 23983 34901 23995 34935
rect 23937 34895 23995 34901
rect 24670 34892 24676 34944
rect 24728 34932 24734 34944
rect 26421 34935 26479 34941
rect 26421 34932 26433 34935
rect 24728 34904 26433 34932
rect 24728 34892 24734 34904
rect 26421 34901 26433 34904
rect 26467 34901 26479 34935
rect 27706 34932 27712 34944
rect 27667 34904 27712 34932
rect 26421 34895 26479 34901
rect 27706 34892 27712 34904
rect 27764 34892 27770 34944
rect 31110 34892 31116 34944
rect 31168 34892 31174 34944
rect 31846 34892 31852 34944
rect 31904 34932 31910 34944
rect 32674 34932 32680 34944
rect 31904 34904 32680 34932
rect 31904 34892 31910 34904
rect 32674 34892 32680 34904
rect 32732 34932 32738 34944
rect 33061 34935 33119 34941
rect 33061 34932 33073 34935
rect 32732 34904 33073 34932
rect 32732 34892 32738 34904
rect 33061 34901 33073 34904
rect 33107 34901 33119 34935
rect 33061 34895 33119 34901
rect 35434 34892 35440 34944
rect 35492 34932 35498 34944
rect 37645 34935 37703 34941
rect 37645 34932 37657 34935
rect 35492 34904 37657 34932
rect 35492 34892 35498 34904
rect 37645 34901 37657 34904
rect 37691 34901 37703 34935
rect 37645 34895 37703 34901
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 4614 34728 4620 34740
rect 4356 34700 4620 34728
rect 4356 34601 4384 34700
rect 4614 34688 4620 34700
rect 4672 34688 4678 34740
rect 5534 34688 5540 34740
rect 5592 34728 5598 34740
rect 5721 34731 5779 34737
rect 5721 34728 5733 34731
rect 5592 34700 5733 34728
rect 5592 34688 5598 34700
rect 5721 34697 5733 34700
rect 5767 34697 5779 34731
rect 5721 34691 5779 34697
rect 7006 34688 7012 34740
rect 7064 34728 7070 34740
rect 9585 34731 9643 34737
rect 9585 34728 9597 34731
rect 7064 34700 9597 34728
rect 7064 34688 7070 34700
rect 9585 34697 9597 34700
rect 9631 34697 9643 34731
rect 10042 34728 10048 34740
rect 10003 34700 10048 34728
rect 9585 34691 9643 34697
rect 10042 34688 10048 34700
rect 10100 34688 10106 34740
rect 19150 34688 19156 34740
rect 19208 34728 19214 34740
rect 20438 34728 20444 34740
rect 19208 34700 20300 34728
rect 20399 34700 20444 34728
rect 19208 34688 19214 34700
rect 8294 34660 8300 34672
rect 7576 34632 8300 34660
rect 4341 34595 4399 34601
rect 4341 34561 4353 34595
rect 4387 34561 4399 34595
rect 4341 34555 4399 34561
rect 4608 34595 4666 34601
rect 4608 34561 4620 34595
rect 4654 34592 4666 34595
rect 5074 34592 5080 34604
rect 4654 34564 5080 34592
rect 4654 34561 4666 34564
rect 4608 34555 4666 34561
rect 5074 34552 5080 34564
rect 5132 34552 5138 34604
rect 7576 34601 7604 34632
rect 8294 34620 8300 34632
rect 8352 34620 8358 34672
rect 9950 34660 9956 34672
rect 9863 34632 9956 34660
rect 9950 34620 9956 34632
rect 10008 34660 10014 34672
rect 16022 34660 16028 34672
rect 10008 34632 16028 34660
rect 10008 34620 10014 34632
rect 16022 34620 16028 34632
rect 16080 34620 16086 34672
rect 19168 34660 19196 34688
rect 18892 34632 19196 34660
rect 7561 34595 7619 34601
rect 7561 34561 7573 34595
rect 7607 34561 7619 34595
rect 7561 34555 7619 34561
rect 7653 34595 7711 34601
rect 7653 34561 7665 34595
rect 7699 34592 7711 34595
rect 7742 34592 7748 34604
rect 7699 34564 7748 34592
rect 7699 34561 7711 34564
rect 7653 34555 7711 34561
rect 7742 34552 7748 34564
rect 7800 34552 7806 34604
rect 7834 34552 7840 34604
rect 7892 34592 7898 34604
rect 17681 34595 17739 34601
rect 7892 34564 7985 34592
rect 7892 34552 7898 34564
rect 17681 34561 17693 34595
rect 17727 34561 17739 34595
rect 18230 34592 18236 34604
rect 18191 34564 18236 34592
rect 17681 34555 17739 34561
rect 7852 34524 7880 34552
rect 8297 34527 8355 34533
rect 8297 34524 8309 34527
rect 7668 34496 7880 34524
rect 8220 34496 8309 34524
rect 5902 34416 5908 34468
rect 5960 34456 5966 34468
rect 7668 34456 7696 34496
rect 5960 34428 7696 34456
rect 5960 34416 5966 34428
rect 7668 34388 7696 34428
rect 7742 34416 7748 34468
rect 7800 34456 7806 34468
rect 8220 34456 8248 34496
rect 8297 34493 8309 34496
rect 8343 34493 8355 34527
rect 8297 34487 8355 34493
rect 10137 34527 10195 34533
rect 10137 34493 10149 34527
rect 10183 34493 10195 34527
rect 11882 34524 11888 34536
rect 10137 34487 10195 34493
rect 10980 34496 11888 34524
rect 10152 34456 10180 34487
rect 10980 34456 11008 34496
rect 11882 34484 11888 34496
rect 11940 34484 11946 34536
rect 17402 34484 17408 34536
rect 17460 34524 17466 34536
rect 17696 34524 17724 34555
rect 18230 34552 18236 34564
rect 18288 34552 18294 34604
rect 18892 34601 18920 34632
rect 19426 34620 19432 34672
rect 19484 34660 19490 34672
rect 20070 34660 20076 34672
rect 19484 34632 20076 34660
rect 19484 34620 19490 34632
rect 20070 34620 20076 34632
rect 20128 34620 20134 34672
rect 20272 34660 20300 34700
rect 20438 34688 20444 34700
rect 20496 34688 20502 34740
rect 23842 34728 23848 34740
rect 21192 34700 23848 34728
rect 20898 34660 20904 34672
rect 20272 34632 20904 34660
rect 20272 34601 20300 34632
rect 20898 34620 20904 34632
rect 20956 34620 20962 34672
rect 21192 34601 21220 34700
rect 23842 34688 23848 34700
rect 23900 34688 23906 34740
rect 30742 34688 30748 34740
rect 30800 34728 30806 34740
rect 33686 34728 33692 34740
rect 30800 34700 33692 34728
rect 30800 34688 30806 34700
rect 33686 34688 33692 34700
rect 33744 34688 33750 34740
rect 36170 34728 36176 34740
rect 36131 34700 36176 34728
rect 36170 34688 36176 34700
rect 36228 34688 36234 34740
rect 21358 34620 21364 34672
rect 21416 34660 21422 34672
rect 27430 34660 27436 34672
rect 21416 34632 27436 34660
rect 21416 34620 21422 34632
rect 18877 34595 18935 34601
rect 18877 34561 18889 34595
rect 18923 34561 18935 34595
rect 18877 34555 18935 34561
rect 19245 34595 19303 34601
rect 19245 34561 19257 34595
rect 19291 34561 19303 34595
rect 19245 34555 19303 34561
rect 20257 34595 20315 34601
rect 20257 34561 20269 34595
rect 20303 34561 20315 34595
rect 20257 34555 20315 34561
rect 21177 34595 21235 34601
rect 21177 34561 21189 34595
rect 21223 34561 21235 34595
rect 21177 34555 21235 34561
rect 21269 34595 21327 34601
rect 21269 34561 21281 34595
rect 21315 34561 21327 34595
rect 21269 34555 21327 34561
rect 21453 34595 21511 34601
rect 21453 34561 21465 34595
rect 21499 34592 21511 34595
rect 21818 34592 21824 34604
rect 21499 34564 21824 34592
rect 21499 34561 21511 34564
rect 21453 34555 21511 34561
rect 17954 34524 17960 34536
rect 17460 34496 17960 34524
rect 17460 34484 17466 34496
rect 17954 34484 17960 34496
rect 18012 34524 18018 34536
rect 19058 34524 19064 34536
rect 18012 34496 19064 34524
rect 18012 34484 18018 34496
rect 19058 34484 19064 34496
rect 19116 34484 19122 34536
rect 18414 34456 18420 34468
rect 7800 34428 8248 34456
rect 10060 34428 11008 34456
rect 17972 34428 18420 34456
rect 7800 34416 7806 34428
rect 10060 34388 10088 34428
rect 17972 34400 18000 34428
rect 18414 34416 18420 34428
rect 18472 34456 18478 34468
rect 19260 34456 19288 34555
rect 19886 34484 19892 34536
rect 19944 34524 19950 34536
rect 20073 34527 20131 34533
rect 20073 34524 20085 34527
rect 19944 34496 20085 34524
rect 19944 34484 19950 34496
rect 20073 34493 20085 34496
rect 20119 34493 20131 34527
rect 21284 34524 21312 34555
rect 21818 34552 21824 34564
rect 21876 34552 21882 34604
rect 22002 34592 22008 34604
rect 21963 34564 22008 34592
rect 22002 34552 22008 34564
rect 22060 34552 22066 34604
rect 22370 34552 22376 34604
rect 22428 34592 22434 34604
rect 23477 34595 23535 34601
rect 23477 34592 23489 34595
rect 22428 34564 23489 34592
rect 22428 34552 22434 34564
rect 23477 34561 23489 34564
rect 23523 34561 23535 34595
rect 23477 34555 23535 34561
rect 24670 34552 24676 34604
rect 24728 34592 24734 34604
rect 25041 34595 25099 34601
rect 25041 34592 25053 34595
rect 24728 34564 25053 34592
rect 24728 34552 24734 34564
rect 25041 34561 25053 34564
rect 25087 34561 25099 34595
rect 25041 34555 25099 34561
rect 25682 34552 25688 34604
rect 25740 34592 25746 34604
rect 27154 34592 27160 34604
rect 25740 34564 27160 34592
rect 25740 34552 25746 34564
rect 27154 34552 27160 34564
rect 27212 34552 27218 34604
rect 27356 34601 27384 34632
rect 27430 34620 27436 34632
rect 27488 34620 27494 34672
rect 34394 34663 34452 34669
rect 34394 34660 34406 34663
rect 33428 34632 34406 34660
rect 27341 34595 27399 34601
rect 27341 34561 27353 34595
rect 27387 34561 27399 34595
rect 27341 34555 27399 34561
rect 28353 34595 28411 34601
rect 28353 34561 28365 34595
rect 28399 34592 28411 34595
rect 28534 34592 28540 34604
rect 28399 34564 28540 34592
rect 28399 34561 28411 34564
rect 28353 34555 28411 34561
rect 28534 34552 28540 34564
rect 28592 34552 28598 34604
rect 29086 34592 29092 34604
rect 29047 34564 29092 34592
rect 29086 34552 29092 34564
rect 29144 34552 29150 34604
rect 32950 34552 32956 34604
rect 33008 34592 33014 34604
rect 33045 34595 33103 34601
rect 33045 34592 33057 34595
rect 33008 34564 33057 34592
rect 33008 34552 33014 34564
rect 33045 34561 33057 34564
rect 33091 34561 33103 34595
rect 33045 34555 33103 34561
rect 22278 34524 22284 34536
rect 20073 34487 20131 34493
rect 20272 34496 22284 34524
rect 20272 34468 20300 34496
rect 22278 34484 22284 34496
rect 22336 34484 22342 34536
rect 22557 34527 22615 34533
rect 22557 34493 22569 34527
rect 22603 34524 22615 34527
rect 23198 34524 23204 34536
rect 22603 34496 23204 34524
rect 22603 34493 22615 34496
rect 22557 34487 22615 34493
rect 23198 34484 23204 34496
rect 23256 34484 23262 34536
rect 23658 34524 23664 34536
rect 23619 34496 23664 34524
rect 23658 34484 23664 34496
rect 23716 34484 23722 34536
rect 25866 34524 25872 34536
rect 25827 34496 25872 34524
rect 25866 34484 25872 34496
rect 25924 34484 25930 34536
rect 28445 34527 28503 34533
rect 28445 34493 28457 34527
rect 28491 34524 28503 34527
rect 29178 34524 29184 34536
rect 28491 34496 29184 34524
rect 28491 34493 28503 34496
rect 28445 34487 28503 34493
rect 29178 34484 29184 34496
rect 29236 34484 29242 34536
rect 32858 34484 32864 34536
rect 32916 34524 32922 34536
rect 33428 34533 33456 34632
rect 34394 34629 34406 34632
rect 34440 34629 34452 34663
rect 34394 34623 34452 34629
rect 34149 34595 34207 34601
rect 34149 34561 34161 34595
rect 34195 34592 34207 34595
rect 34238 34592 34244 34604
rect 34195 34564 34244 34592
rect 34195 34561 34207 34564
rect 34149 34555 34207 34561
rect 34238 34552 34244 34564
rect 34296 34552 34302 34604
rect 35434 34552 35440 34604
rect 35492 34592 35498 34604
rect 36541 34595 36599 34601
rect 36541 34592 36553 34595
rect 35492 34564 36553 34592
rect 35492 34552 35498 34564
rect 36541 34561 36553 34564
rect 36587 34561 36599 34595
rect 37829 34595 37887 34601
rect 37829 34592 37841 34595
rect 36541 34555 36599 34561
rect 36648 34564 37841 34592
rect 36648 34536 36676 34564
rect 37829 34561 37841 34564
rect 37875 34561 37887 34595
rect 37829 34555 37887 34561
rect 33137 34527 33195 34533
rect 33137 34524 33149 34527
rect 32916 34496 33149 34524
rect 32916 34484 32922 34496
rect 33137 34493 33149 34496
rect 33183 34493 33195 34527
rect 33137 34487 33195 34493
rect 33413 34527 33471 34533
rect 33413 34493 33425 34527
rect 33459 34493 33471 34527
rect 36630 34524 36636 34536
rect 36591 34496 36636 34524
rect 33413 34487 33471 34493
rect 36630 34484 36636 34496
rect 36688 34484 36694 34536
rect 36817 34527 36875 34533
rect 36817 34493 36829 34527
rect 36863 34493 36875 34527
rect 38102 34524 38108 34536
rect 38063 34496 38108 34524
rect 36817 34487 36875 34493
rect 20254 34456 20260 34468
rect 18472 34428 20260 34456
rect 18472 34416 18478 34428
rect 20254 34416 20260 34428
rect 20312 34416 20318 34468
rect 22465 34459 22523 34465
rect 22465 34425 22477 34459
rect 22511 34456 22523 34459
rect 23566 34456 23572 34468
rect 22511 34428 23572 34456
rect 22511 34425 22523 34428
rect 22465 34419 22523 34425
rect 23566 34416 23572 34428
rect 23624 34416 23630 34468
rect 36832 34456 36860 34487
rect 38102 34484 38108 34496
rect 38160 34484 38166 34536
rect 38010 34456 38016 34468
rect 36832 34428 38016 34456
rect 38010 34416 38016 34428
rect 38068 34416 38074 34468
rect 7668 34360 10088 34388
rect 17954 34348 17960 34400
rect 18012 34348 18018 34400
rect 18138 34388 18144 34400
rect 18099 34360 18144 34388
rect 18138 34348 18144 34360
rect 18196 34348 18202 34400
rect 18230 34348 18236 34400
rect 18288 34388 18294 34400
rect 19886 34388 19892 34400
rect 18288 34360 19892 34388
rect 18288 34348 18294 34360
rect 19886 34348 19892 34360
rect 19944 34388 19950 34400
rect 22370 34388 22376 34400
rect 19944 34360 22376 34388
rect 19944 34348 19950 34360
rect 22370 34348 22376 34360
rect 22428 34348 22434 34400
rect 22646 34388 22652 34400
rect 22607 34360 22652 34388
rect 22646 34348 22652 34360
rect 22704 34348 22710 34400
rect 25130 34348 25136 34400
rect 25188 34388 25194 34400
rect 27433 34391 27491 34397
rect 27433 34388 27445 34391
rect 25188 34360 27445 34388
rect 25188 34348 25194 34360
rect 27433 34357 27445 34360
rect 27479 34357 27491 34391
rect 27433 34351 27491 34357
rect 28994 34348 29000 34400
rect 29052 34388 29058 34400
rect 29181 34391 29239 34397
rect 29181 34388 29193 34391
rect 29052 34360 29193 34388
rect 29052 34348 29058 34360
rect 29181 34357 29193 34360
rect 29227 34357 29239 34391
rect 29181 34351 29239 34357
rect 30742 34348 30748 34400
rect 30800 34388 30806 34400
rect 35342 34388 35348 34400
rect 30800 34360 35348 34388
rect 30800 34348 30806 34360
rect 35342 34348 35348 34360
rect 35400 34388 35406 34400
rect 35529 34391 35587 34397
rect 35529 34388 35541 34391
rect 35400 34360 35541 34388
rect 35400 34348 35406 34360
rect 35529 34357 35541 34360
rect 35575 34357 35587 34391
rect 35529 34351 35587 34357
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 10226 34144 10232 34196
rect 10284 34184 10290 34196
rect 10689 34187 10747 34193
rect 10689 34184 10701 34187
rect 10284 34156 10701 34184
rect 10284 34144 10290 34156
rect 10689 34153 10701 34156
rect 10735 34153 10747 34187
rect 20898 34184 20904 34196
rect 10689 34147 10747 34153
rect 18524 34156 20904 34184
rect 11149 34119 11207 34125
rect 11149 34085 11161 34119
rect 11195 34116 11207 34119
rect 11195 34088 12434 34116
rect 11195 34085 11207 34088
rect 11149 34079 11207 34085
rect 5534 34008 5540 34060
rect 5592 34048 5598 34060
rect 5813 34051 5871 34057
rect 5813 34048 5825 34051
rect 5592 34020 5825 34048
rect 5592 34008 5598 34020
rect 5813 34017 5825 34020
rect 5859 34017 5871 34051
rect 5813 34011 5871 34017
rect 5902 34008 5908 34060
rect 5960 34048 5966 34060
rect 8202 34048 8208 34060
rect 5960 34020 6005 34048
rect 8163 34020 8208 34048
rect 5960 34008 5966 34020
rect 8202 34008 8208 34020
rect 8260 34008 8266 34060
rect 9674 34008 9680 34060
rect 9732 34048 9738 34060
rect 9861 34051 9919 34057
rect 9861 34048 9873 34051
rect 9732 34020 9873 34048
rect 9732 34008 9738 34020
rect 9861 34017 9873 34020
rect 9907 34017 9919 34051
rect 9861 34011 9919 34017
rect 10873 34051 10931 34057
rect 10873 34017 10885 34051
rect 10919 34048 10931 34051
rect 11330 34048 11336 34060
rect 10919 34020 11336 34048
rect 10919 34017 10931 34020
rect 10873 34011 10931 34017
rect 11330 34008 11336 34020
rect 11388 34008 11394 34060
rect 12406 34048 12434 34088
rect 17678 34048 17684 34060
rect 12406 34020 17684 34048
rect 5718 33980 5724 33992
rect 5679 33952 5724 33980
rect 5718 33940 5724 33952
rect 5776 33940 5782 33992
rect 7742 33980 7748 33992
rect 7703 33952 7748 33980
rect 7742 33940 7748 33952
rect 7800 33940 7806 33992
rect 8113 33983 8171 33989
rect 8113 33949 8125 33983
rect 8159 33949 8171 33983
rect 8220 33980 8248 34008
rect 10594 33980 10600 33992
rect 8220 33952 10600 33980
rect 8113 33943 8171 33949
rect 8128 33912 8156 33943
rect 10594 33940 10600 33952
rect 10652 33980 10658 33992
rect 10689 33983 10747 33989
rect 10689 33980 10701 33983
rect 10652 33952 10701 33980
rect 10652 33940 10658 33952
rect 10689 33949 10701 33952
rect 10735 33949 10747 33983
rect 10689 33943 10747 33949
rect 10965 33983 11023 33989
rect 10965 33949 10977 33983
rect 11011 33980 11023 33983
rect 11146 33980 11152 33992
rect 11011 33952 11152 33980
rect 11011 33949 11023 33952
rect 10965 33943 11023 33949
rect 11146 33940 11152 33952
rect 11204 33940 11210 33992
rect 11882 33980 11888 33992
rect 11843 33952 11888 33980
rect 11882 33940 11888 33952
rect 11940 33940 11946 33992
rect 12069 33983 12127 33989
rect 12069 33949 12081 33983
rect 12115 33980 12127 33983
rect 12250 33980 12256 33992
rect 12115 33952 12256 33980
rect 12115 33949 12127 33952
rect 12069 33943 12127 33949
rect 12250 33940 12256 33952
rect 12308 33940 12314 33992
rect 14642 33940 14648 33992
rect 14700 33980 14706 33992
rect 15289 33983 15347 33989
rect 15289 33980 15301 33983
rect 14700 33952 15301 33980
rect 14700 33940 14706 33952
rect 15289 33949 15301 33952
rect 15335 33949 15347 33983
rect 15289 33943 15347 33949
rect 15473 33983 15531 33989
rect 15473 33949 15485 33983
rect 15519 33980 15531 33983
rect 15838 33980 15844 33992
rect 15519 33952 15844 33980
rect 15519 33949 15531 33952
rect 15473 33943 15531 33949
rect 15838 33940 15844 33952
rect 15896 33940 15902 33992
rect 16776 33989 16804 34020
rect 17678 34008 17684 34020
rect 17736 34008 17742 34060
rect 16761 33983 16819 33989
rect 16761 33949 16773 33983
rect 16807 33949 16819 33983
rect 16761 33943 16819 33949
rect 16945 33983 17003 33989
rect 16945 33949 16957 33983
rect 16991 33980 17003 33983
rect 18524 33980 18552 34156
rect 20898 34144 20904 34156
rect 20956 34144 20962 34196
rect 21726 34144 21732 34196
rect 21784 34184 21790 34196
rect 23014 34184 23020 34196
rect 21784 34156 23020 34184
rect 21784 34144 21790 34156
rect 23014 34144 23020 34156
rect 23072 34144 23078 34196
rect 23842 34144 23848 34196
rect 23900 34184 23906 34196
rect 25406 34184 25412 34196
rect 23900 34156 25412 34184
rect 23900 34144 23906 34156
rect 25406 34144 25412 34156
rect 25464 34184 25470 34196
rect 25774 34184 25780 34196
rect 25464 34156 25780 34184
rect 25464 34144 25470 34156
rect 25774 34144 25780 34156
rect 25832 34144 25838 34196
rect 26237 34187 26295 34193
rect 26237 34153 26249 34187
rect 26283 34184 26295 34187
rect 27246 34184 27252 34196
rect 26283 34156 27252 34184
rect 26283 34153 26295 34156
rect 26237 34147 26295 34153
rect 27246 34144 27252 34156
rect 27304 34144 27310 34196
rect 30377 34187 30435 34193
rect 30377 34153 30389 34187
rect 30423 34184 30435 34187
rect 31754 34184 31760 34196
rect 30423 34156 31760 34184
rect 30423 34153 30435 34156
rect 30377 34147 30435 34153
rect 31754 34144 31760 34156
rect 31812 34144 31818 34196
rect 31846 34144 31852 34196
rect 31904 34184 31910 34196
rect 35250 34184 35256 34196
rect 31904 34156 31949 34184
rect 32968 34156 35256 34184
rect 31904 34144 31910 34156
rect 18598 34076 18604 34128
rect 18656 34116 18662 34128
rect 26694 34116 26700 34128
rect 18656 34088 26556 34116
rect 26655 34088 26700 34116
rect 18656 34076 18662 34088
rect 19518 34048 19524 34060
rect 16991 33952 18552 33980
rect 18616 34020 19524 34048
rect 16991 33949 17003 33952
rect 16945 33943 17003 33949
rect 8478 33912 8484 33924
rect 8128 33884 8484 33912
rect 8478 33872 8484 33884
rect 8536 33872 8542 33924
rect 9122 33912 9128 33924
rect 9083 33884 9128 33912
rect 9122 33872 9128 33884
rect 9180 33872 9186 33924
rect 16574 33872 16580 33924
rect 16632 33912 16638 33924
rect 17405 33915 17463 33921
rect 17405 33912 17417 33915
rect 16632 33884 17417 33912
rect 16632 33872 16638 33884
rect 17405 33881 17417 33884
rect 17451 33912 17463 33915
rect 17451 33884 17724 33912
rect 17451 33881 17463 33884
rect 17405 33875 17463 33881
rect 5350 33844 5356 33856
rect 5311 33816 5356 33844
rect 5350 33804 5356 33816
rect 5408 33804 5414 33856
rect 11977 33847 12035 33853
rect 11977 33813 11989 33847
rect 12023 33844 12035 33847
rect 14090 33844 14096 33856
rect 12023 33816 14096 33844
rect 12023 33813 12035 33816
rect 11977 33807 12035 33813
rect 14090 33804 14096 33816
rect 14148 33804 14154 33856
rect 15381 33847 15439 33853
rect 15381 33813 15393 33847
rect 15427 33844 15439 33847
rect 15470 33844 15476 33856
rect 15427 33816 15476 33844
rect 15427 33813 15439 33816
rect 15381 33807 15439 33813
rect 15470 33804 15476 33816
rect 15528 33804 15534 33856
rect 16945 33847 17003 33853
rect 16945 33813 16957 33847
rect 16991 33844 17003 33847
rect 17586 33844 17592 33856
rect 16991 33816 17592 33844
rect 16991 33813 17003 33816
rect 16945 33807 17003 33813
rect 17586 33804 17592 33816
rect 17644 33804 17650 33856
rect 17696 33844 17724 33884
rect 17954 33872 17960 33924
rect 18012 33912 18018 33924
rect 18141 33915 18199 33921
rect 18141 33912 18153 33915
rect 18012 33884 18153 33912
rect 18012 33872 18018 33884
rect 18141 33881 18153 33884
rect 18187 33881 18199 33915
rect 18141 33875 18199 33881
rect 18616 33844 18644 34020
rect 19518 34008 19524 34020
rect 19576 34008 19582 34060
rect 21177 34051 21235 34057
rect 21177 34048 21189 34051
rect 19628 34020 21189 34048
rect 19242 33940 19248 33992
rect 19300 33980 19306 33992
rect 19628 33989 19656 34020
rect 21177 34017 21189 34020
rect 21223 34048 21235 34051
rect 21542 34048 21548 34060
rect 21223 34020 21548 34048
rect 21223 34017 21235 34020
rect 21177 34011 21235 34017
rect 21542 34008 21548 34020
rect 21600 34008 21606 34060
rect 22278 34008 22284 34060
rect 22336 34048 22342 34060
rect 25866 34048 25872 34060
rect 22336 34020 25268 34048
rect 25827 34020 25872 34048
rect 22336 34008 22342 34020
rect 19429 33983 19487 33989
rect 19429 33980 19441 33983
rect 19300 33952 19441 33980
rect 19300 33940 19306 33952
rect 19429 33949 19441 33952
rect 19475 33949 19487 33983
rect 19429 33943 19487 33949
rect 19613 33983 19671 33989
rect 19613 33949 19625 33983
rect 19659 33949 19671 33983
rect 19613 33943 19671 33949
rect 20073 33983 20131 33989
rect 20073 33949 20085 33983
rect 20119 33949 20131 33983
rect 20254 33980 20260 33992
rect 20215 33952 20260 33980
rect 20073 33943 20131 33949
rect 19058 33872 19064 33924
rect 19116 33912 19122 33924
rect 20088 33912 20116 33943
rect 20254 33940 20260 33952
rect 20312 33940 20318 33992
rect 21269 33983 21327 33989
rect 21269 33949 21281 33983
rect 21315 33980 21327 33983
rect 22370 33980 22376 33992
rect 21315 33952 22140 33980
rect 22331 33952 22376 33980
rect 21315 33949 21327 33952
rect 21269 33943 21327 33949
rect 19116 33884 20116 33912
rect 19116 33872 19122 33884
rect 20806 33872 20812 33924
rect 20864 33912 20870 33924
rect 21545 33915 21603 33921
rect 21545 33912 21557 33915
rect 20864 33884 21557 33912
rect 20864 33872 20870 33884
rect 21545 33881 21557 33884
rect 21591 33881 21603 33915
rect 21545 33875 21603 33881
rect 17696 33816 18644 33844
rect 19426 33804 19432 33856
rect 19484 33844 19490 33856
rect 19521 33847 19579 33853
rect 19521 33844 19533 33847
rect 19484 33816 19533 33844
rect 19484 33804 19490 33816
rect 19521 33813 19533 33816
rect 19567 33813 19579 33847
rect 19521 33807 19579 33813
rect 19978 33804 19984 33856
rect 20036 33844 20042 33856
rect 20165 33847 20223 33853
rect 20165 33844 20177 33847
rect 20036 33816 20177 33844
rect 20036 33804 20042 33816
rect 20165 33813 20177 33816
rect 20211 33844 20223 33847
rect 20254 33844 20260 33856
rect 20211 33816 20260 33844
rect 20211 33813 20223 33816
rect 20165 33807 20223 33813
rect 20254 33804 20260 33816
rect 20312 33804 20318 33856
rect 20714 33804 20720 33856
rect 20772 33844 20778 33856
rect 20993 33847 21051 33853
rect 20993 33844 21005 33847
rect 20772 33816 21005 33844
rect 20772 33804 20778 33816
rect 20993 33813 21005 33816
rect 21039 33813 21051 33847
rect 21560 33844 21588 33875
rect 21634 33872 21640 33924
rect 21692 33912 21698 33924
rect 22112 33921 22140 33952
rect 22370 33940 22376 33952
rect 22428 33940 22434 33992
rect 22465 33983 22523 33989
rect 22465 33949 22477 33983
rect 22511 33949 22523 33983
rect 22465 33943 22523 33949
rect 22557 33983 22615 33989
rect 22557 33949 22569 33983
rect 22603 33980 22615 33983
rect 22646 33980 22652 33992
rect 22603 33952 22652 33980
rect 22603 33949 22615 33952
rect 22557 33943 22615 33949
rect 22097 33915 22155 33921
rect 21692 33884 21737 33912
rect 21692 33872 21698 33884
rect 22097 33881 22109 33915
rect 22143 33881 22155 33915
rect 22097 33875 22155 33881
rect 22186 33872 22192 33924
rect 22244 33912 22250 33924
rect 22480 33912 22508 33943
rect 22646 33940 22652 33952
rect 22704 33940 22710 33992
rect 22738 33940 22744 33992
rect 22796 33980 22802 33992
rect 23566 33980 23572 33992
rect 22796 33952 22841 33980
rect 23527 33952 23572 33980
rect 22796 33940 22802 33952
rect 23566 33940 23572 33952
rect 23624 33940 23630 33992
rect 23842 33980 23848 33992
rect 23803 33952 23848 33980
rect 23842 33940 23848 33952
rect 23900 33940 23906 33992
rect 24762 33980 24768 33992
rect 24723 33952 24768 33980
rect 24762 33940 24768 33952
rect 24820 33940 24826 33992
rect 24949 33983 25007 33989
rect 24949 33949 24961 33983
rect 24995 33949 25007 33983
rect 24949 33943 25007 33949
rect 22244 33884 22508 33912
rect 22244 33872 22250 33884
rect 22278 33844 22284 33856
rect 21560 33816 22284 33844
rect 20993 33807 21051 33813
rect 22278 33804 22284 33816
rect 22336 33804 22342 33856
rect 22480 33844 22508 33884
rect 23014 33872 23020 33924
rect 23072 33912 23078 33924
rect 24964 33912 24992 33943
rect 25038 33940 25044 33992
rect 25096 33980 25102 33992
rect 25133 33983 25191 33989
rect 25133 33980 25145 33983
rect 25096 33952 25145 33980
rect 25096 33940 25102 33952
rect 25133 33949 25145 33952
rect 25179 33949 25191 33983
rect 25240 33980 25268 34020
rect 25866 34008 25872 34020
rect 25924 34008 25930 34060
rect 26528 34048 26556 34088
rect 26694 34076 26700 34088
rect 26752 34076 26758 34128
rect 31938 34116 31944 34128
rect 29012 34088 29684 34116
rect 29012 34060 29040 34088
rect 28905 34051 28963 34057
rect 26528 34020 28488 34048
rect 26053 33983 26111 33989
rect 26053 33980 26065 33983
rect 25240 33952 26065 33980
rect 25133 33943 25191 33949
rect 26053 33949 26065 33952
rect 26099 33949 26111 33983
rect 26053 33943 26111 33949
rect 26973 33983 27031 33989
rect 26973 33949 26985 33983
rect 27019 33980 27031 33983
rect 27338 33980 27344 33992
rect 27019 33952 27344 33980
rect 27019 33949 27031 33952
rect 26973 33943 27031 33949
rect 27338 33940 27344 33952
rect 27396 33940 27402 33992
rect 27525 33983 27583 33989
rect 27525 33949 27537 33983
rect 27571 33980 27583 33983
rect 27706 33980 27712 33992
rect 27571 33952 27712 33980
rect 27571 33949 27583 33952
rect 27525 33943 27583 33949
rect 27706 33940 27712 33952
rect 27764 33940 27770 33992
rect 25590 33912 25596 33924
rect 23072 33884 25596 33912
rect 23072 33872 23078 33884
rect 25590 33872 25596 33884
rect 25648 33912 25654 33924
rect 25777 33915 25835 33921
rect 25777 33912 25789 33915
rect 25648 33884 25789 33912
rect 25648 33872 25654 33884
rect 25777 33881 25789 33884
rect 25823 33881 25835 33915
rect 26697 33915 26755 33921
rect 26697 33912 26709 33915
rect 25777 33875 25835 33881
rect 25884 33884 26709 33912
rect 22738 33844 22744 33856
rect 22480 33816 22744 33844
rect 22738 33804 22744 33816
rect 22796 33804 22802 33856
rect 25682 33804 25688 33856
rect 25740 33844 25746 33856
rect 25884 33844 25912 33884
rect 26697 33881 26709 33884
rect 26743 33881 26755 33915
rect 26697 33875 26755 33881
rect 26786 33872 26792 33924
rect 26844 33912 26850 33924
rect 26881 33915 26939 33921
rect 26881 33912 26893 33915
rect 26844 33884 26893 33912
rect 26844 33872 26850 33884
rect 26881 33881 26893 33884
rect 26927 33881 26939 33915
rect 27890 33912 27896 33924
rect 27851 33884 27896 33912
rect 26881 33875 26939 33881
rect 27890 33872 27896 33884
rect 27948 33872 27954 33924
rect 28460 33912 28488 34020
rect 28905 34017 28917 34051
rect 28951 34048 28963 34051
rect 28994 34048 29000 34060
rect 28951 34020 29000 34048
rect 28951 34017 28963 34020
rect 28905 34011 28963 34017
rect 28994 34008 29000 34020
rect 29052 34008 29058 34060
rect 29089 34051 29147 34057
rect 29089 34017 29101 34051
rect 29135 34048 29147 34051
rect 29270 34048 29276 34060
rect 29135 34020 29276 34048
rect 29135 34017 29147 34020
rect 29089 34011 29147 34017
rect 29270 34008 29276 34020
rect 29328 34008 29334 34060
rect 29656 33992 29684 34088
rect 30116 34088 31944 34116
rect 29178 33940 29184 33992
rect 29236 33980 29242 33992
rect 29638 33980 29644 33992
rect 29236 33952 29281 33980
rect 29551 33952 29644 33980
rect 29236 33940 29242 33952
rect 29638 33940 29644 33952
rect 29696 33980 29702 33992
rect 29733 33983 29791 33989
rect 29733 33980 29745 33983
rect 29696 33952 29745 33980
rect 29696 33940 29702 33952
rect 29733 33949 29745 33952
rect 29779 33949 29791 33983
rect 29733 33943 29791 33949
rect 29881 33983 29939 33989
rect 29881 33949 29893 33983
rect 29927 33980 29939 33983
rect 30116 33980 30144 34088
rect 31938 34076 31944 34088
rect 31996 34116 32002 34128
rect 32968 34116 32996 34156
rect 35250 34144 35256 34156
rect 35308 34184 35314 34196
rect 35434 34184 35440 34196
rect 35308 34156 35440 34184
rect 35308 34144 35314 34156
rect 35434 34144 35440 34156
rect 35492 34144 35498 34196
rect 31996 34088 32996 34116
rect 31996 34076 32002 34088
rect 33042 34076 33048 34128
rect 33100 34116 33106 34128
rect 37826 34116 37832 34128
rect 33100 34088 37832 34116
rect 33100 34076 33106 34088
rect 37826 34076 37832 34088
rect 37884 34076 37890 34128
rect 36078 34048 36084 34060
rect 31496 34020 36084 34048
rect 29927 33952 30144 33980
rect 29927 33949 29939 33952
rect 29881 33943 29939 33949
rect 30190 33940 30196 33992
rect 30248 33989 30254 33992
rect 30248 33980 30256 33989
rect 31202 33980 31208 33992
rect 30248 33952 30293 33980
rect 31163 33952 31208 33980
rect 30248 33943 30256 33952
rect 30248 33940 30254 33943
rect 31202 33940 31208 33952
rect 31260 33940 31266 33992
rect 31294 33940 31300 33992
rect 31352 33980 31358 33992
rect 31496 33980 31524 34020
rect 36078 34008 36084 34020
rect 36136 34008 36142 34060
rect 31662 33980 31668 33992
rect 31720 33989 31726 33992
rect 31352 33952 31524 33980
rect 31628 33952 31668 33980
rect 31352 33940 31358 33952
rect 31662 33940 31668 33952
rect 31720 33943 31728 33989
rect 31720 33940 31726 33943
rect 37182 33940 37188 33992
rect 37240 33980 37246 33992
rect 37829 33983 37887 33989
rect 37829 33980 37841 33983
rect 37240 33952 37841 33980
rect 37240 33940 37246 33952
rect 37829 33949 37841 33952
rect 37875 33949 37887 33983
rect 37829 33943 37887 33949
rect 30006 33912 30012 33924
rect 28460 33884 29868 33912
rect 29967 33884 30012 33912
rect 25740 33816 25912 33844
rect 25740 33804 25746 33816
rect 26510 33804 26516 33856
rect 26568 33844 26574 33856
rect 26804 33844 26832 33872
rect 28718 33844 28724 33856
rect 26568 33816 26832 33844
rect 28679 33816 28724 33844
rect 26568 33804 26574 33816
rect 28718 33804 28724 33816
rect 28776 33804 28782 33856
rect 29840 33844 29868 33884
rect 30006 33872 30012 33884
rect 30064 33872 30070 33924
rect 30098 33872 30104 33924
rect 30156 33912 30162 33924
rect 30156 33884 30201 33912
rect 30156 33872 30162 33884
rect 31110 33872 31116 33924
rect 31168 33912 31174 33924
rect 31481 33915 31539 33921
rect 31481 33912 31493 33915
rect 31168 33884 31493 33912
rect 31168 33872 31174 33884
rect 31481 33881 31493 33884
rect 31527 33881 31539 33915
rect 31481 33875 31539 33881
rect 31573 33915 31631 33921
rect 31573 33881 31585 33915
rect 31619 33912 31631 33915
rect 34514 33912 34520 33924
rect 31619 33884 34520 33912
rect 31619 33881 31631 33884
rect 31573 33875 31631 33881
rect 31588 33844 31616 33875
rect 34514 33872 34520 33884
rect 34572 33872 34578 33924
rect 38102 33912 38108 33924
rect 38063 33884 38108 33912
rect 38102 33872 38108 33884
rect 38160 33872 38166 33924
rect 29840 33816 31616 33844
rect 32674 33804 32680 33856
rect 32732 33844 32738 33856
rect 35526 33844 35532 33856
rect 32732 33816 35532 33844
rect 32732 33804 32738 33816
rect 35526 33804 35532 33816
rect 35584 33804 35590 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 13541 33643 13599 33649
rect 13541 33609 13553 33643
rect 13587 33640 13599 33643
rect 13630 33640 13636 33652
rect 13587 33612 13636 33640
rect 13587 33609 13599 33612
rect 13541 33603 13599 33609
rect 13630 33600 13636 33612
rect 13688 33600 13694 33652
rect 14642 33640 14648 33652
rect 14603 33612 14648 33640
rect 14642 33600 14648 33612
rect 14700 33600 14706 33652
rect 16025 33643 16083 33649
rect 16025 33609 16037 33643
rect 16071 33640 16083 33643
rect 16206 33640 16212 33652
rect 16071 33612 16212 33640
rect 16071 33609 16083 33612
rect 16025 33603 16083 33609
rect 16206 33600 16212 33612
rect 16264 33600 16270 33652
rect 17494 33600 17500 33652
rect 17552 33640 17558 33652
rect 19061 33643 19119 33649
rect 19061 33640 19073 33643
rect 17552 33612 19073 33640
rect 17552 33600 17558 33612
rect 19061 33609 19073 33612
rect 19107 33609 19119 33643
rect 19061 33603 19119 33609
rect 19334 33600 19340 33652
rect 19392 33640 19398 33652
rect 20441 33643 20499 33649
rect 20441 33640 20453 33643
rect 19392 33612 20453 33640
rect 19392 33600 19398 33612
rect 20441 33609 20453 33612
rect 20487 33609 20499 33643
rect 20441 33603 20499 33609
rect 21361 33643 21419 33649
rect 21361 33609 21373 33643
rect 21407 33640 21419 33643
rect 21634 33640 21640 33652
rect 21407 33612 21640 33640
rect 21407 33609 21419 33612
rect 21361 33603 21419 33609
rect 21634 33600 21640 33612
rect 21692 33600 21698 33652
rect 22738 33600 22744 33652
rect 22796 33640 22802 33652
rect 24210 33640 24216 33652
rect 22796 33612 24216 33640
rect 22796 33600 22802 33612
rect 24210 33600 24216 33612
rect 24268 33600 24274 33652
rect 25501 33643 25559 33649
rect 25501 33609 25513 33643
rect 25547 33640 25559 33643
rect 27338 33640 27344 33652
rect 25547 33612 27344 33640
rect 25547 33609 25559 33612
rect 25501 33603 25559 33609
rect 27338 33600 27344 33612
rect 27396 33600 27402 33652
rect 28718 33600 28724 33652
rect 28776 33640 28782 33652
rect 31110 33640 31116 33652
rect 28776 33612 31116 33640
rect 28776 33600 28782 33612
rect 31110 33600 31116 33612
rect 31168 33600 31174 33652
rect 31665 33643 31723 33649
rect 31665 33609 31677 33643
rect 31711 33640 31723 33643
rect 32858 33640 32864 33652
rect 31711 33612 32864 33640
rect 31711 33609 31723 33612
rect 31665 33603 31723 33609
rect 32858 33600 32864 33612
rect 32916 33600 32922 33652
rect 35710 33640 35716 33652
rect 33152 33612 35716 33640
rect 7374 33572 7380 33584
rect 5368 33544 7380 33572
rect 5166 33464 5172 33516
rect 5224 33504 5230 33516
rect 5368 33513 5396 33544
rect 7374 33532 7380 33544
rect 7432 33572 7438 33584
rect 8478 33572 8484 33584
rect 7432 33544 8484 33572
rect 7432 33532 7438 33544
rect 8478 33532 8484 33544
rect 8536 33572 8542 33584
rect 9306 33572 9312 33584
rect 8536 33544 9312 33572
rect 8536 33532 8542 33544
rect 9306 33532 9312 33544
rect 9364 33572 9370 33584
rect 23382 33572 23388 33584
rect 9364 33544 10548 33572
rect 9364 33532 9370 33544
rect 5353 33507 5411 33513
rect 5353 33504 5365 33507
rect 5224 33476 5365 33504
rect 5224 33464 5230 33476
rect 5353 33473 5365 33476
rect 5399 33473 5411 33507
rect 5353 33467 5411 33473
rect 5445 33507 5503 33513
rect 5445 33473 5457 33507
rect 5491 33473 5503 33507
rect 5445 33467 5503 33473
rect 5905 33507 5963 33513
rect 5905 33473 5917 33507
rect 5951 33504 5963 33507
rect 6546 33504 6552 33516
rect 5951 33476 6552 33504
rect 5951 33473 5963 33476
rect 5905 33467 5963 33473
rect 5460 33436 5488 33467
rect 6546 33464 6552 33476
rect 6604 33464 6610 33516
rect 7006 33504 7012 33516
rect 6967 33476 7012 33504
rect 7006 33464 7012 33476
rect 7064 33464 7070 33516
rect 8110 33504 8116 33516
rect 8071 33476 8116 33504
rect 8110 33464 8116 33476
rect 8168 33464 8174 33516
rect 8297 33507 8355 33513
rect 8297 33473 8309 33507
rect 8343 33504 8355 33507
rect 8386 33504 8392 33516
rect 8343 33476 8392 33504
rect 8343 33473 8355 33476
rect 8297 33467 8355 33473
rect 8386 33464 8392 33476
rect 8444 33464 8450 33516
rect 10520 33513 10548 33544
rect 13188 33544 15792 33572
rect 10229 33507 10287 33513
rect 10229 33473 10241 33507
rect 10275 33473 10287 33507
rect 10229 33467 10287 33473
rect 10505 33507 10563 33513
rect 10505 33473 10517 33507
rect 10551 33473 10563 33507
rect 12066 33504 12072 33516
rect 12027 33476 12072 33504
rect 10505 33467 10563 33473
rect 7285 33439 7343 33445
rect 7285 33436 7297 33439
rect 5460 33408 7297 33436
rect 7285 33405 7297 33408
rect 7331 33436 7343 33439
rect 7466 33436 7472 33448
rect 7331 33408 7472 33436
rect 7331 33405 7343 33408
rect 7285 33399 7343 33405
rect 7466 33396 7472 33408
rect 7524 33396 7530 33448
rect 10244 33436 10272 33467
rect 12066 33464 12072 33476
rect 12124 33464 12130 33516
rect 12250 33504 12256 33516
rect 12211 33476 12256 33504
rect 12250 33464 12256 33476
rect 12308 33464 12314 33516
rect 13188 33513 13216 33544
rect 13173 33507 13231 33513
rect 13173 33473 13185 33507
rect 13219 33473 13231 33507
rect 13173 33467 13231 33473
rect 13265 33507 13323 33513
rect 13265 33473 13277 33507
rect 13311 33473 13323 33507
rect 13265 33467 13323 33473
rect 13357 33507 13415 33513
rect 13357 33473 13369 33507
rect 13403 33504 13415 33507
rect 14001 33507 14059 33513
rect 14001 33504 14013 33507
rect 13403 33476 14013 33504
rect 13403 33473 13415 33476
rect 13357 33467 13415 33473
rect 14001 33473 14013 33476
rect 14047 33504 14059 33507
rect 14182 33504 14188 33516
rect 14047 33476 14188 33504
rect 14047 33473 14059 33476
rect 14001 33467 14059 33473
rect 11330 33436 11336 33448
rect 10244 33408 11336 33436
rect 11330 33396 11336 33408
rect 11388 33396 11394 33448
rect 13280 33436 13308 33467
rect 14182 33464 14188 33476
rect 14240 33464 14246 33516
rect 14461 33507 14519 33513
rect 14461 33473 14473 33507
rect 14507 33504 14519 33507
rect 14550 33504 14556 33516
rect 14507 33476 14556 33504
rect 14507 33473 14519 33476
rect 14461 33467 14519 33473
rect 14550 33464 14556 33476
rect 14608 33504 14614 33516
rect 15010 33504 15016 33516
rect 14608 33476 15016 33504
rect 14608 33464 14614 33476
rect 15010 33464 15016 33476
rect 15068 33464 15074 33516
rect 15378 33504 15384 33516
rect 15339 33476 15384 33504
rect 15378 33464 15384 33476
rect 15436 33464 15442 33516
rect 13538 33436 13544 33448
rect 13280 33408 13544 33436
rect 13538 33396 13544 33408
rect 13596 33396 13602 33448
rect 14366 33436 14372 33448
rect 14327 33408 14372 33436
rect 14366 33396 14372 33408
rect 14424 33396 14430 33448
rect 14642 33396 14648 33448
rect 14700 33436 14706 33448
rect 15657 33439 15715 33445
rect 15657 33436 15669 33439
rect 14700 33408 15669 33436
rect 14700 33396 14706 33408
rect 15657 33405 15669 33408
rect 15703 33405 15715 33439
rect 15764 33436 15792 33544
rect 15856 33544 23388 33572
rect 15856 33513 15884 33544
rect 15841 33507 15899 33513
rect 15841 33473 15853 33507
rect 15887 33473 15899 33507
rect 17402 33504 17408 33516
rect 17363 33476 17408 33504
rect 15841 33467 15899 33473
rect 17402 33464 17408 33476
rect 17460 33464 17466 33516
rect 18230 33504 18236 33516
rect 17880 33476 18236 33504
rect 16942 33436 16948 33448
rect 15764 33408 16948 33436
rect 15657 33399 15715 33405
rect 16942 33396 16948 33408
rect 17000 33396 17006 33448
rect 17313 33439 17371 33445
rect 17313 33405 17325 33439
rect 17359 33436 17371 33439
rect 17770 33436 17776 33448
rect 17359 33408 17776 33436
rect 17359 33405 17371 33408
rect 17313 33399 17371 33405
rect 17770 33396 17776 33408
rect 17828 33396 17834 33448
rect 17880 33445 17908 33476
rect 18230 33464 18236 33476
rect 18288 33464 18294 33516
rect 19245 33507 19303 33513
rect 19245 33473 19257 33507
rect 19291 33473 19303 33507
rect 19245 33467 19303 33473
rect 17865 33439 17923 33445
rect 17865 33405 17877 33439
rect 17911 33405 17923 33439
rect 19150 33436 19156 33448
rect 17865 33399 17923 33405
rect 17972 33408 19156 33436
rect 12069 33371 12127 33377
rect 12069 33337 12081 33371
rect 12115 33368 12127 33371
rect 15194 33368 15200 33380
rect 12115 33340 15200 33368
rect 12115 33337 12127 33340
rect 12069 33331 12127 33337
rect 15194 33328 15200 33340
rect 15252 33328 15258 33380
rect 15838 33328 15844 33380
rect 15896 33368 15902 33380
rect 17494 33368 17500 33380
rect 15896 33340 17500 33368
rect 15896 33328 15902 33340
rect 17494 33328 17500 33340
rect 17552 33328 17558 33380
rect 6822 33260 6828 33312
rect 6880 33300 6886 33312
rect 8389 33303 8447 33309
rect 8389 33300 8401 33303
rect 6880 33272 8401 33300
rect 6880 33260 6886 33272
rect 8389 33269 8401 33272
rect 8435 33269 8447 33303
rect 8389 33263 8447 33269
rect 9950 33260 9956 33312
rect 10008 33300 10014 33312
rect 10045 33303 10103 33309
rect 10045 33300 10057 33303
rect 10008 33272 10057 33300
rect 10008 33260 10014 33272
rect 10045 33269 10057 33272
rect 10091 33269 10103 33303
rect 14090 33300 14096 33312
rect 14051 33272 14096 33300
rect 10045 33263 10103 33269
rect 14090 33260 14096 33272
rect 14148 33260 14154 33312
rect 14182 33260 14188 33312
rect 14240 33300 14246 33312
rect 14826 33300 14832 33312
rect 14240 33272 14832 33300
rect 14240 33260 14246 33272
rect 14826 33260 14832 33272
rect 14884 33260 14890 33312
rect 15470 33300 15476 33312
rect 15431 33272 15476 33300
rect 15470 33260 15476 33272
rect 15528 33260 15534 33312
rect 17773 33303 17831 33309
rect 17773 33269 17785 33303
rect 17819 33300 17831 33303
rect 17972 33300 18000 33408
rect 19150 33396 19156 33408
rect 19208 33396 19214 33448
rect 19260 33368 19288 33467
rect 19334 33464 19340 33516
rect 19392 33504 19398 33516
rect 19536 33513 19564 33544
rect 23382 33532 23388 33544
rect 23440 33532 23446 33584
rect 25130 33572 25136 33584
rect 24136 33544 25136 33572
rect 19521 33507 19579 33513
rect 19392 33476 19437 33504
rect 19392 33464 19398 33476
rect 19521 33473 19533 33507
rect 19567 33473 19579 33507
rect 19521 33467 19579 33473
rect 19613 33507 19671 33513
rect 19613 33473 19625 33507
rect 19659 33473 19671 33507
rect 19613 33467 19671 33473
rect 19426 33396 19432 33448
rect 19484 33436 19490 33448
rect 19628 33436 19656 33467
rect 19794 33464 19800 33516
rect 19852 33504 19858 33516
rect 20257 33507 20315 33513
rect 20257 33504 20269 33507
rect 19852 33476 20269 33504
rect 19852 33464 19858 33476
rect 20257 33473 20269 33476
rect 20303 33473 20315 33507
rect 20257 33467 20315 33473
rect 20346 33464 20352 33516
rect 20404 33504 20410 33516
rect 20533 33507 20591 33513
rect 20533 33504 20545 33507
rect 20404 33476 20545 33504
rect 20404 33464 20410 33476
rect 20533 33473 20545 33476
rect 20579 33473 20591 33507
rect 21266 33504 21272 33516
rect 21227 33476 21272 33504
rect 20533 33467 20591 33473
rect 21266 33464 21272 33476
rect 21324 33464 21330 33516
rect 22462 33464 22468 33516
rect 22520 33504 22526 33516
rect 22738 33504 22744 33516
rect 22520 33476 22565 33504
rect 22699 33476 22744 33504
rect 22520 33464 22526 33476
rect 22738 33464 22744 33476
rect 22796 33464 22802 33516
rect 24136 33504 24164 33544
rect 25130 33532 25136 33544
rect 25188 33572 25194 33584
rect 28905 33575 28963 33581
rect 28905 33572 28917 33575
rect 25188 33544 26280 33572
rect 25188 33532 25194 33544
rect 26252 33516 26280 33544
rect 27540 33544 28917 33572
rect 22848 33476 24164 33504
rect 22094 33436 22100 33448
rect 19484 33408 22100 33436
rect 19484 33396 19490 33408
rect 22094 33396 22100 33408
rect 22152 33396 22158 33448
rect 22557 33439 22615 33445
rect 22557 33405 22569 33439
rect 22603 33436 22615 33439
rect 22848 33436 22876 33476
rect 24210 33464 24216 33516
rect 24268 33504 24274 33516
rect 24268 33476 24313 33504
rect 24762 33494 24768 33516
rect 24268 33464 24274 33476
rect 24688 33466 24768 33494
rect 22603 33408 22876 33436
rect 22925 33439 22983 33445
rect 22603 33405 22615 33408
rect 22557 33399 22615 33405
rect 22925 33405 22937 33439
rect 22971 33405 22983 33439
rect 22925 33399 22983 33405
rect 23661 33439 23719 33445
rect 23661 33405 23673 33439
rect 23707 33436 23719 33439
rect 23750 33436 23756 33448
rect 23707 33408 23756 33436
rect 23707 33405 23719 33408
rect 23661 33399 23719 33405
rect 20346 33368 20352 33380
rect 19260 33340 20352 33368
rect 20346 33328 20352 33340
rect 20404 33328 20410 33380
rect 17819 33272 18000 33300
rect 18141 33303 18199 33309
rect 17819 33269 17831 33272
rect 17773 33263 17831 33269
rect 18141 33269 18153 33303
rect 18187 33300 18199 33303
rect 19242 33300 19248 33312
rect 18187 33272 19248 33300
rect 18187 33269 18199 33272
rect 18141 33263 18199 33269
rect 19242 33260 19248 33272
rect 19300 33260 19306 33312
rect 20073 33303 20131 33309
rect 20073 33269 20085 33303
rect 20119 33300 20131 33303
rect 20806 33300 20812 33312
rect 20119 33272 20812 33300
rect 20119 33269 20131 33272
rect 20073 33263 20131 33269
rect 20806 33260 20812 33272
rect 20864 33260 20870 33312
rect 20898 33260 20904 33312
rect 20956 33300 20962 33312
rect 21450 33300 21456 33312
rect 20956 33272 21456 33300
rect 20956 33260 20962 33272
rect 21450 33260 21456 33272
rect 21508 33300 21514 33312
rect 22940 33300 22968 33399
rect 23750 33396 23756 33408
rect 23808 33396 23814 33448
rect 24026 33436 24032 33448
rect 23987 33408 24032 33436
rect 24026 33396 24032 33408
rect 24084 33396 24090 33448
rect 24121 33439 24179 33445
rect 24121 33405 24133 33439
rect 24167 33436 24179 33439
rect 24688 33436 24716 33466
rect 24762 33464 24768 33466
rect 24820 33504 24826 33516
rect 24857 33507 24915 33513
rect 24857 33504 24869 33507
rect 24820 33476 24869 33504
rect 24820 33464 24826 33476
rect 24857 33473 24869 33476
rect 24903 33473 24915 33507
rect 26234 33504 26240 33516
rect 24857 33467 24915 33473
rect 25148 33476 26096 33504
rect 26147 33476 26240 33504
rect 25148 33436 25176 33476
rect 24167 33408 24716 33436
rect 24780 33408 25176 33436
rect 25225 33439 25283 33445
rect 24167 33405 24179 33408
rect 24121 33399 24179 33405
rect 23198 33328 23204 33380
rect 23256 33368 23262 33380
rect 24780 33368 24808 33408
rect 25225 33405 25237 33439
rect 25271 33405 25283 33439
rect 26068 33436 26096 33476
rect 26234 33464 26240 33476
rect 26292 33464 26298 33516
rect 26418 33504 26424 33516
rect 26379 33476 26424 33504
rect 26418 33464 26424 33476
rect 26476 33464 26482 33516
rect 27540 33513 27568 33544
rect 28905 33541 28917 33544
rect 28951 33541 28963 33575
rect 28905 33535 28963 33541
rect 30926 33532 30932 33584
rect 30984 33572 30990 33584
rect 31297 33575 31355 33581
rect 31297 33572 31309 33575
rect 30984 33544 31309 33572
rect 30984 33532 30990 33544
rect 31297 33541 31309 33544
rect 31343 33541 31355 33575
rect 31297 33535 31355 33541
rect 31386 33532 31392 33584
rect 31444 33572 31450 33584
rect 32674 33572 32680 33584
rect 31444 33544 32680 33572
rect 31444 33532 31450 33544
rect 32674 33532 32680 33544
rect 32732 33532 32738 33584
rect 33152 33581 33180 33612
rect 35710 33600 35716 33612
rect 35768 33600 35774 33652
rect 36081 33643 36139 33649
rect 36081 33609 36093 33643
rect 36127 33640 36139 33643
rect 36630 33640 36636 33652
rect 36127 33612 36636 33640
rect 36127 33609 36139 33612
rect 36081 33603 36139 33609
rect 36630 33600 36636 33612
rect 36688 33600 36694 33652
rect 33137 33575 33195 33581
rect 33137 33541 33149 33575
rect 33183 33541 33195 33575
rect 33137 33535 33195 33541
rect 33229 33575 33287 33581
rect 33229 33541 33241 33575
rect 33275 33572 33287 33575
rect 33686 33572 33692 33584
rect 33275 33544 33692 33572
rect 33275 33541 33287 33544
rect 33229 33535 33287 33541
rect 33686 33532 33692 33544
rect 33744 33532 33750 33584
rect 34698 33581 34704 33584
rect 34697 33535 34704 33581
rect 34756 33572 34762 33584
rect 34756 33544 34797 33572
rect 34698 33532 34704 33535
rect 34756 33532 34762 33544
rect 27525 33507 27583 33513
rect 27525 33504 27537 33507
rect 26528 33476 27537 33504
rect 26528 33436 26556 33476
rect 27525 33473 27537 33476
rect 27571 33473 27583 33507
rect 27525 33467 27583 33473
rect 27614 33464 27620 33516
rect 27672 33504 27678 33516
rect 28721 33507 28779 33513
rect 28721 33504 28733 33507
rect 27672 33476 28733 33504
rect 27672 33464 27678 33476
rect 28721 33473 28733 33476
rect 28767 33473 28779 33507
rect 28721 33467 28779 33473
rect 29733 33507 29791 33513
rect 29733 33473 29745 33507
rect 29779 33473 29791 33507
rect 31018 33504 31024 33516
rect 30979 33476 31024 33504
rect 29733 33467 29791 33473
rect 26068 33408 26556 33436
rect 25225 33399 25283 33405
rect 23256 33340 24808 33368
rect 23256 33328 23262 33340
rect 24854 33328 24860 33380
rect 24912 33368 24918 33380
rect 25240 33368 25268 33399
rect 26878 33396 26884 33448
rect 26936 33436 26942 33448
rect 27801 33439 27859 33445
rect 27801 33436 27813 33439
rect 26936 33408 27813 33436
rect 26936 33396 26942 33408
rect 27801 33405 27813 33408
rect 27847 33405 27859 33439
rect 27801 33399 27859 33405
rect 27982 33396 27988 33448
rect 28040 33436 28046 33448
rect 28997 33439 29055 33445
rect 28997 33436 29009 33439
rect 28040 33408 29009 33436
rect 28040 33396 28046 33408
rect 28997 33405 29009 33408
rect 29043 33405 29055 33439
rect 28997 33399 29055 33405
rect 24912 33340 25268 33368
rect 26513 33371 26571 33377
rect 24912 33328 24918 33340
rect 26513 33337 26525 33371
rect 26559 33368 26571 33371
rect 27430 33368 27436 33380
rect 26559 33340 27436 33368
rect 26559 33337 26571 33340
rect 26513 33331 26571 33337
rect 27430 33328 27436 33340
rect 27488 33368 27494 33380
rect 29086 33368 29092 33380
rect 27488 33340 29092 33368
rect 27488 33328 27494 33340
rect 29086 33328 29092 33340
rect 29144 33368 29150 33380
rect 29748 33368 29776 33467
rect 31018 33464 31024 33476
rect 31076 33464 31082 33516
rect 31114 33507 31172 33513
rect 31114 33473 31126 33507
rect 31160 33473 31172 33507
rect 31114 33467 31172 33473
rect 29822 33396 29828 33448
rect 29880 33436 29886 33448
rect 30009 33439 30067 33445
rect 30009 33436 30021 33439
rect 29880 33408 30021 33436
rect 29880 33396 29886 33408
rect 30009 33405 30021 33408
rect 30055 33405 30067 33439
rect 30009 33399 30067 33405
rect 30742 33396 30748 33448
rect 30800 33436 30806 33448
rect 31128 33436 31156 33467
rect 31478 33464 31484 33516
rect 31536 33513 31542 33516
rect 31536 33504 31544 33513
rect 32858 33504 32864 33516
rect 31536 33476 31581 33504
rect 32819 33476 32864 33504
rect 31536 33467 31544 33476
rect 31536 33464 31542 33467
rect 32858 33464 32864 33476
rect 32916 33464 32922 33516
rect 32954 33507 33012 33513
rect 32954 33473 32966 33507
rect 33000 33504 33012 33507
rect 33042 33504 33048 33516
rect 33000 33476 33048 33504
rect 33000 33473 33012 33476
rect 32954 33467 33012 33473
rect 30800 33408 31156 33436
rect 30800 33396 30806 33408
rect 29144 33340 29776 33368
rect 29144 33328 29150 33340
rect 29914 33328 29920 33380
rect 29972 33368 29978 33380
rect 32968 33368 32996 33467
rect 33042 33464 33048 33476
rect 33100 33464 33106 33516
rect 33367 33507 33425 33513
rect 33367 33473 33379 33507
rect 33413 33504 33425 33507
rect 34330 33504 34336 33516
rect 33413 33476 34336 33504
rect 33413 33473 33425 33476
rect 33367 33467 33425 33473
rect 34330 33464 34336 33476
rect 34388 33464 34394 33516
rect 34422 33464 34428 33516
rect 34480 33504 34486 33516
rect 34606 33513 34612 33516
rect 34563 33507 34612 33513
rect 34480 33476 34525 33504
rect 34480 33464 34486 33476
rect 34563 33473 34575 33507
rect 34609 33473 34612 33507
rect 34563 33467 34612 33473
rect 34606 33464 34612 33467
rect 34664 33464 34670 33516
rect 34793 33507 34851 33513
rect 34793 33473 34805 33507
rect 34839 33504 34851 33507
rect 34882 33504 34888 33516
rect 34839 33476 34888 33504
rect 34839 33473 34851 33476
rect 34793 33467 34851 33473
rect 34882 33464 34888 33476
rect 34940 33464 34946 33516
rect 35437 33507 35495 33513
rect 35437 33504 35449 33507
rect 34992 33476 35449 33504
rect 34992 33377 35020 33476
rect 35437 33473 35449 33476
rect 35483 33473 35495 33507
rect 35437 33467 35495 33473
rect 35530 33507 35588 33513
rect 35530 33473 35542 33507
rect 35576 33473 35588 33507
rect 35710 33504 35716 33516
rect 35671 33476 35716 33504
rect 35530 33467 35588 33473
rect 35250 33396 35256 33448
rect 35308 33436 35314 33448
rect 35544 33436 35572 33467
rect 35710 33464 35716 33476
rect 35768 33464 35774 33516
rect 35805 33507 35863 33513
rect 35805 33473 35817 33507
rect 35851 33473 35863 33507
rect 35805 33467 35863 33473
rect 35308 33408 35572 33436
rect 35308 33396 35314 33408
rect 35618 33396 35624 33448
rect 35676 33436 35682 33448
rect 35820 33436 35848 33467
rect 35894 33464 35900 33516
rect 35952 33513 35958 33516
rect 35952 33504 35960 33513
rect 36170 33504 36176 33516
rect 35952 33476 36176 33504
rect 35952 33467 35960 33476
rect 35952 33464 35958 33467
rect 36170 33464 36176 33476
rect 36228 33464 36234 33516
rect 37826 33504 37832 33516
rect 37787 33476 37832 33504
rect 37826 33464 37832 33476
rect 37884 33464 37890 33516
rect 35676 33408 35848 33436
rect 35676 33396 35682 33408
rect 36354 33396 36360 33448
rect 36412 33436 36418 33448
rect 37182 33436 37188 33448
rect 36412 33408 37188 33436
rect 36412 33396 36418 33408
rect 37182 33396 37188 33408
rect 37240 33436 37246 33448
rect 37921 33439 37979 33445
rect 37921 33436 37933 33439
rect 37240 33408 37933 33436
rect 37240 33396 37246 33408
rect 37921 33405 37933 33408
rect 37967 33405 37979 33439
rect 37921 33399 37979 33405
rect 38010 33396 38016 33448
rect 38068 33436 38074 33448
rect 38068 33408 38113 33436
rect 38068 33396 38074 33408
rect 29972 33340 32996 33368
rect 34977 33371 35035 33377
rect 29972 33328 29978 33340
rect 34977 33337 34989 33371
rect 35023 33337 35035 33371
rect 37734 33368 37740 33380
rect 34977 33331 35035 33337
rect 36832 33340 37740 33368
rect 21508 33272 22968 33300
rect 21508 33260 21514 33272
rect 23750 33260 23756 33312
rect 23808 33300 23814 33312
rect 24995 33303 25053 33309
rect 24995 33300 25007 33303
rect 23808 33272 25007 33300
rect 23808 33260 23814 33272
rect 24995 33269 25007 33272
rect 25041 33269 25053 33303
rect 24995 33263 25053 33269
rect 25133 33303 25191 33309
rect 25133 33269 25145 33303
rect 25179 33300 25191 33303
rect 25774 33300 25780 33312
rect 25179 33272 25780 33300
rect 25179 33269 25191 33272
rect 25133 33263 25191 33269
rect 25774 33260 25780 33272
rect 25832 33260 25838 33312
rect 33505 33303 33563 33309
rect 33505 33269 33517 33303
rect 33551 33300 33563 33303
rect 36832 33300 36860 33340
rect 37734 33328 37740 33340
rect 37792 33328 37798 33380
rect 33551 33272 36860 33300
rect 33551 33269 33563 33272
rect 33505 33263 33563 33269
rect 37090 33260 37096 33312
rect 37148 33300 37154 33312
rect 37461 33303 37519 33309
rect 37461 33300 37473 33303
rect 37148 33272 37473 33300
rect 37148 33260 37154 33272
rect 37461 33269 37473 33272
rect 37507 33269 37519 33303
rect 37461 33263 37519 33269
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 6825 33099 6883 33105
rect 6825 33065 6837 33099
rect 6871 33096 6883 33099
rect 10226 33096 10232 33108
rect 6871 33068 10232 33096
rect 6871 33065 6883 33068
rect 6825 33059 6883 33065
rect 10226 33056 10232 33068
rect 10284 33056 10290 33108
rect 10873 33099 10931 33105
rect 10873 33065 10885 33099
rect 10919 33065 10931 33099
rect 10873 33059 10931 33065
rect 12069 33099 12127 33105
rect 12069 33065 12081 33099
rect 12115 33096 12127 33099
rect 13538 33096 13544 33108
rect 12115 33068 13544 33096
rect 12115 33065 12127 33068
rect 12069 33059 12127 33065
rect 7745 33031 7803 33037
rect 7745 32997 7757 33031
rect 7791 33028 7803 33031
rect 8110 33028 8116 33040
rect 7791 33000 8116 33028
rect 7791 32997 7803 33000
rect 7745 32991 7803 32997
rect 8110 32988 8116 33000
rect 8168 33028 8174 33040
rect 8297 33031 8355 33037
rect 8297 33028 8309 33031
rect 8168 33000 8309 33028
rect 8168 32988 8174 33000
rect 8297 32997 8309 33000
rect 8343 32997 8355 33031
rect 8297 32991 8355 32997
rect 9674 32988 9680 33040
rect 9732 33028 9738 33040
rect 10888 33028 10916 33059
rect 13538 33056 13544 33068
rect 13596 33056 13602 33108
rect 13722 33056 13728 33108
rect 13780 33096 13786 33108
rect 15654 33096 15660 33108
rect 13780 33068 15660 33096
rect 13780 33056 13786 33068
rect 15654 33056 15660 33068
rect 15712 33056 15718 33108
rect 15838 33096 15844 33108
rect 15799 33068 15844 33096
rect 15838 33056 15844 33068
rect 15896 33056 15902 33108
rect 15930 33056 15936 33108
rect 15988 33096 15994 33108
rect 16025 33099 16083 33105
rect 16025 33096 16037 33099
rect 15988 33068 16037 33096
rect 15988 33056 15994 33068
rect 16025 33065 16037 33068
rect 16071 33065 16083 33099
rect 16025 33059 16083 33065
rect 17589 33099 17647 33105
rect 17589 33065 17601 33099
rect 17635 33065 17647 33099
rect 17589 33059 17647 33065
rect 17773 33099 17831 33105
rect 17773 33065 17785 33099
rect 17819 33096 17831 33099
rect 18046 33096 18052 33108
rect 17819 33068 18052 33096
rect 17819 33065 17831 33068
rect 17773 33059 17831 33065
rect 9732 33000 10916 33028
rect 11333 33031 11391 33037
rect 9732 32988 9738 33000
rect 11333 32997 11345 33031
rect 11379 33028 11391 33031
rect 17604 33028 17632 33059
rect 18046 33056 18052 33068
rect 18104 33056 18110 33108
rect 18138 33056 18144 33108
rect 18196 33096 18202 33108
rect 18322 33096 18328 33108
rect 18196 33068 18328 33096
rect 18196 33056 18202 33068
rect 18322 33056 18328 33068
rect 18380 33056 18386 33108
rect 20162 33056 20168 33108
rect 20220 33096 20226 33108
rect 20346 33096 20352 33108
rect 20220 33068 20352 33096
rect 20220 33056 20226 33068
rect 20346 33056 20352 33068
rect 20404 33056 20410 33108
rect 20530 33056 20536 33108
rect 20588 33096 20594 33108
rect 22646 33096 22652 33108
rect 20588 33068 22652 33096
rect 20588 33056 20594 33068
rect 22646 33056 22652 33068
rect 22704 33056 22710 33108
rect 25222 33096 25228 33108
rect 25183 33068 25228 33096
rect 25222 33056 25228 33068
rect 25280 33056 25286 33108
rect 30377 33099 30435 33105
rect 30377 33065 30389 33099
rect 30423 33096 30435 33099
rect 30650 33096 30656 33108
rect 30423 33068 30656 33096
rect 30423 33065 30435 33068
rect 30377 33059 30435 33065
rect 30650 33056 30656 33068
rect 30708 33056 30714 33108
rect 31202 33056 31208 33108
rect 31260 33096 31266 33108
rect 31481 33099 31539 33105
rect 31481 33096 31493 33099
rect 31260 33068 31493 33096
rect 31260 33056 31266 33068
rect 31481 33065 31493 33068
rect 31527 33065 31539 33099
rect 31481 33059 31539 33065
rect 32493 33099 32551 33105
rect 32493 33065 32505 33099
rect 32539 33096 32551 33099
rect 32858 33096 32864 33108
rect 32539 33068 32864 33096
rect 32539 33065 32551 33068
rect 32493 33059 32551 33065
rect 32858 33056 32864 33068
rect 32916 33056 32922 33108
rect 35710 33056 35716 33108
rect 35768 33096 35774 33108
rect 36354 33096 36360 33108
rect 35768 33068 36032 33096
rect 36315 33068 36360 33096
rect 35768 33056 35774 33068
rect 20714 33028 20720 33040
rect 11379 33000 16436 33028
rect 17604 33000 20720 33028
rect 11379 32997 11391 33000
rect 11333 32991 11391 32997
rect 4614 32960 4620 32972
rect 4448 32932 4620 32960
rect 4448 32901 4476 32932
rect 4614 32920 4620 32932
rect 4672 32960 4678 32972
rect 5350 32960 5356 32972
rect 4672 32932 5356 32960
rect 4672 32920 4678 32932
rect 5350 32920 5356 32932
rect 5408 32920 5414 32972
rect 5810 32920 5816 32972
rect 5868 32960 5874 32972
rect 5868 32932 8248 32960
rect 5868 32920 5874 32932
rect 4433 32895 4491 32901
rect 4433 32861 4445 32895
rect 4479 32861 4491 32895
rect 4433 32855 4491 32861
rect 4522 32852 4528 32904
rect 4580 32892 4586 32904
rect 5166 32892 5172 32904
rect 4580 32864 5172 32892
rect 4580 32852 4586 32864
rect 5166 32852 5172 32864
rect 5224 32852 5230 32904
rect 5258 32852 5264 32904
rect 5316 32892 5322 32904
rect 6733 32895 6791 32901
rect 5316 32864 5361 32892
rect 5316 32852 5322 32864
rect 6733 32861 6745 32895
rect 6779 32861 6791 32895
rect 6733 32855 6791 32861
rect 6917 32895 6975 32901
rect 6917 32861 6929 32895
rect 6963 32892 6975 32895
rect 7374 32892 7380 32904
rect 6963 32864 7380 32892
rect 6963 32861 6975 32864
rect 6917 32855 6975 32861
rect 4706 32824 4712 32836
rect 4667 32796 4712 32824
rect 4706 32784 4712 32796
rect 4764 32784 4770 32836
rect 5718 32824 5724 32836
rect 5679 32796 5724 32824
rect 5718 32784 5724 32796
rect 5776 32784 5782 32836
rect 6748 32824 6776 32855
rect 7374 32852 7380 32864
rect 7432 32852 7438 32904
rect 7561 32895 7619 32901
rect 7561 32861 7573 32895
rect 7607 32892 7619 32895
rect 7742 32892 7748 32904
rect 7607 32864 7748 32892
rect 7607 32861 7619 32864
rect 7561 32855 7619 32861
rect 7742 32852 7748 32864
rect 7800 32852 7806 32904
rect 8220 32901 8248 32932
rect 8386 32920 8392 32972
rect 8444 32960 8450 32972
rect 8481 32963 8539 32969
rect 8481 32960 8493 32963
rect 8444 32932 8493 32960
rect 8444 32920 8450 32932
rect 8481 32929 8493 32932
rect 8527 32960 8539 32963
rect 9766 32960 9772 32972
rect 8527 32932 9772 32960
rect 8527 32929 8539 32932
rect 8481 32923 8539 32929
rect 9766 32920 9772 32932
rect 9824 32920 9830 32972
rect 10045 32963 10103 32969
rect 10045 32929 10057 32963
rect 10091 32960 10103 32963
rect 10134 32960 10140 32972
rect 10091 32932 10140 32960
rect 10091 32929 10103 32932
rect 10045 32923 10103 32929
rect 10134 32920 10140 32932
rect 10192 32960 10198 32972
rect 10965 32963 11023 32969
rect 10192 32932 10916 32960
rect 10192 32920 10198 32932
rect 8205 32895 8263 32901
rect 8205 32861 8217 32895
rect 8251 32861 8263 32895
rect 8205 32855 8263 32861
rect 9214 32852 9220 32904
rect 9272 32892 9278 32904
rect 9677 32895 9735 32901
rect 9677 32892 9689 32895
rect 9272 32864 9689 32892
rect 9272 32852 9278 32864
rect 9677 32861 9689 32864
rect 9723 32861 9735 32895
rect 9858 32892 9864 32904
rect 9819 32864 9864 32892
rect 9677 32855 9735 32861
rect 9858 32852 9864 32864
rect 9916 32852 9922 32904
rect 9953 32895 10011 32901
rect 9953 32861 9965 32895
rect 9999 32861 10011 32895
rect 10226 32892 10232 32904
rect 10187 32864 10232 32892
rect 9953 32855 10011 32861
rect 7466 32824 7472 32836
rect 6748 32796 7472 32824
rect 7466 32784 7472 32796
rect 7524 32784 7530 32836
rect 9968 32824 9996 32855
rect 10226 32852 10232 32864
rect 10284 32852 10290 32904
rect 10888 32892 10916 32932
rect 10965 32929 10977 32963
rect 11011 32960 11023 32963
rect 11238 32960 11244 32972
rect 11011 32932 11244 32960
rect 11011 32929 11023 32932
rect 10965 32923 11023 32929
rect 11238 32920 11244 32932
rect 11296 32920 11302 32972
rect 12437 32963 12495 32969
rect 12437 32960 12449 32963
rect 11348 32932 12449 32960
rect 11146 32892 11152 32904
rect 10888 32864 11008 32892
rect 11107 32864 11152 32892
rect 9968 32796 10548 32824
rect 8481 32759 8539 32765
rect 8481 32725 8493 32759
rect 8527 32756 8539 32759
rect 9582 32756 9588 32768
rect 8527 32728 9588 32756
rect 8527 32725 8539 32728
rect 8481 32719 8539 32725
rect 9582 32716 9588 32728
rect 9640 32716 9646 32768
rect 10410 32756 10416 32768
rect 10371 32728 10416 32756
rect 10410 32716 10416 32728
rect 10468 32716 10474 32768
rect 10520 32756 10548 32796
rect 10594 32784 10600 32836
rect 10652 32824 10658 32836
rect 10873 32827 10931 32833
rect 10873 32824 10885 32827
rect 10652 32796 10885 32824
rect 10652 32784 10658 32796
rect 10873 32793 10885 32796
rect 10919 32793 10931 32827
rect 10980 32824 11008 32864
rect 11146 32852 11152 32864
rect 11204 32852 11210 32904
rect 11348 32824 11376 32932
rect 12437 32929 12449 32932
rect 12483 32929 12495 32963
rect 12437 32923 12495 32929
rect 13354 32920 13360 32972
rect 13412 32960 13418 32972
rect 15013 32963 15071 32969
rect 15013 32960 15025 32963
rect 13412 32932 15025 32960
rect 13412 32920 13418 32932
rect 15013 32929 15025 32932
rect 15059 32929 15071 32963
rect 15013 32923 15071 32929
rect 15378 32920 15384 32972
rect 15436 32960 15442 32972
rect 15749 32963 15807 32969
rect 15749 32960 15761 32963
rect 15436 32932 15761 32960
rect 15436 32920 15442 32932
rect 15749 32929 15761 32932
rect 15795 32929 15807 32963
rect 15749 32923 15807 32929
rect 12250 32892 12256 32904
rect 12211 32864 12256 32892
rect 12250 32852 12256 32864
rect 12308 32852 12314 32904
rect 12345 32895 12403 32901
rect 12345 32861 12357 32895
rect 12391 32861 12403 32895
rect 12526 32892 12532 32904
rect 12487 32864 12532 32892
rect 12345 32855 12403 32861
rect 10980 32796 11376 32824
rect 10873 32787 10931 32793
rect 11974 32784 11980 32836
rect 12032 32824 12038 32836
rect 12360 32824 12388 32855
rect 12526 32852 12532 32864
rect 12584 32852 12590 32904
rect 13538 32892 13544 32904
rect 13499 32864 13544 32892
rect 13538 32852 13544 32864
rect 13596 32852 13602 32904
rect 13722 32892 13728 32904
rect 13683 32864 13728 32892
rect 13722 32852 13728 32864
rect 13780 32852 13786 32904
rect 15102 32852 15108 32904
rect 15160 32892 15166 32904
rect 15657 32895 15715 32901
rect 15657 32892 15669 32895
rect 15160 32864 15669 32892
rect 15160 32852 15166 32864
rect 15657 32861 15669 32864
rect 15703 32861 15715 32895
rect 16408 32892 16436 33000
rect 20714 32988 20720 33000
rect 20772 32988 20778 33040
rect 22738 33028 22744 33040
rect 22699 33000 22744 33028
rect 22738 32988 22744 33000
rect 22796 32988 22802 33040
rect 23382 32988 23388 33040
rect 23440 33028 23446 33040
rect 25409 33031 25467 33037
rect 25409 33028 25421 33031
rect 23440 33000 25421 33028
rect 23440 32988 23446 33000
rect 25409 32997 25421 33000
rect 25455 32997 25467 33031
rect 25409 32991 25467 32997
rect 26234 32988 26240 33040
rect 26292 32988 26298 33040
rect 30190 33028 30196 33040
rect 27448 33000 30196 33028
rect 17497 32963 17555 32969
rect 17497 32929 17509 32963
rect 17543 32960 17555 32963
rect 17770 32960 17776 32972
rect 17543 32932 17776 32960
rect 17543 32929 17555 32932
rect 17497 32923 17555 32929
rect 17770 32920 17776 32932
rect 17828 32920 17834 32972
rect 18509 32963 18567 32969
rect 18509 32929 18521 32963
rect 18555 32929 18567 32963
rect 20993 32963 21051 32969
rect 18509 32923 18567 32929
rect 19720 32932 20668 32960
rect 17586 32892 17592 32904
rect 16408 32864 17448 32892
rect 17547 32864 17592 32892
rect 15657 32855 15715 32861
rect 12802 32824 12808 32836
rect 12032 32796 12808 32824
rect 12032 32784 12038 32796
rect 12802 32784 12808 32796
rect 12860 32784 12866 32836
rect 13814 32784 13820 32836
rect 13872 32824 13878 32836
rect 14277 32827 14335 32833
rect 14277 32824 14289 32827
rect 13872 32796 14289 32824
rect 13872 32784 13878 32796
rect 14277 32793 14289 32796
rect 14323 32793 14335 32827
rect 14277 32787 14335 32793
rect 15194 32784 15200 32836
rect 15252 32824 15258 32836
rect 17313 32827 17371 32833
rect 17313 32824 17325 32827
rect 15252 32796 17325 32824
rect 15252 32784 15258 32796
rect 17313 32793 17325 32796
rect 17359 32793 17371 32827
rect 17420 32824 17448 32864
rect 17586 32852 17592 32864
rect 17644 32852 17650 32904
rect 17862 32852 17868 32904
rect 17920 32892 17926 32904
rect 18233 32895 18291 32901
rect 18233 32892 18245 32895
rect 17920 32864 18245 32892
rect 17920 32852 17926 32864
rect 18233 32861 18245 32864
rect 18279 32861 18291 32895
rect 18233 32855 18291 32861
rect 18138 32824 18144 32836
rect 17420 32796 18144 32824
rect 17313 32787 17371 32793
rect 18138 32784 18144 32796
rect 18196 32824 18202 32836
rect 18524 32824 18552 32923
rect 19720 32901 19748 32932
rect 19705 32895 19763 32901
rect 19705 32861 19717 32895
rect 19751 32861 19763 32895
rect 19705 32855 19763 32861
rect 19889 32895 19947 32901
rect 19889 32861 19901 32895
rect 19935 32892 19947 32895
rect 20162 32892 20168 32904
rect 19935 32864 20168 32892
rect 19935 32861 19947 32864
rect 19889 32855 19947 32861
rect 20162 32852 20168 32864
rect 20220 32852 20226 32904
rect 20530 32892 20536 32904
rect 20491 32864 20536 32892
rect 20530 32852 20536 32864
rect 20588 32852 20594 32904
rect 20640 32901 20668 32932
rect 20993 32929 21005 32963
rect 21039 32960 21051 32963
rect 21634 32960 21640 32972
rect 21039 32932 21640 32960
rect 21039 32929 21051 32932
rect 20993 32923 21051 32929
rect 21634 32920 21640 32932
rect 21692 32920 21698 32972
rect 22462 32960 22468 32972
rect 21928 32932 22468 32960
rect 20625 32895 20683 32901
rect 20625 32861 20637 32895
rect 20671 32892 20683 32895
rect 20714 32892 20720 32904
rect 20671 32864 20720 32892
rect 20671 32861 20683 32864
rect 20625 32855 20683 32861
rect 20714 32852 20720 32864
rect 20772 32852 20778 32904
rect 21928 32901 21956 32932
rect 22462 32920 22468 32932
rect 22520 32960 22526 32972
rect 23014 32960 23020 32972
rect 22520 32932 23020 32960
rect 22520 32920 22526 32932
rect 21913 32895 21971 32901
rect 21913 32861 21925 32895
rect 21959 32861 21971 32895
rect 21913 32855 21971 32861
rect 22005 32895 22063 32901
rect 22005 32861 22017 32895
rect 22051 32892 22063 32895
rect 22554 32892 22560 32904
rect 22051 32864 22560 32892
rect 22051 32861 22063 32864
rect 22005 32855 22063 32861
rect 20898 32824 20904 32836
rect 18196 32796 18552 32824
rect 20859 32796 20904 32824
rect 18196 32784 18202 32796
rect 20898 32784 20904 32796
rect 20956 32824 20962 32836
rect 22020 32824 22048 32855
rect 22554 32852 22560 32864
rect 22612 32852 22618 32904
rect 22664 32901 22692 32932
rect 23014 32920 23020 32932
rect 23072 32920 23078 32972
rect 24765 32963 24823 32969
rect 24765 32929 24777 32963
rect 24811 32960 24823 32963
rect 24946 32960 24952 32972
rect 24811 32932 24952 32960
rect 24811 32929 24823 32932
rect 24765 32923 24823 32929
rect 24946 32920 24952 32932
rect 25004 32920 25010 32972
rect 26252 32960 26280 32988
rect 27448 32969 27476 33000
rect 30190 32988 30196 33000
rect 30248 32988 30254 33040
rect 30944 33000 35849 33028
rect 26160 32932 26280 32960
rect 27433 32963 27491 32969
rect 22649 32895 22707 32901
rect 22649 32861 22661 32895
rect 22695 32861 22707 32895
rect 22649 32855 22707 32861
rect 22925 32895 22983 32901
rect 22925 32861 22937 32895
rect 22971 32892 22983 32895
rect 23566 32892 23572 32904
rect 22971 32864 23572 32892
rect 22971 32861 22983 32864
rect 22925 32855 22983 32861
rect 23566 32852 23572 32864
rect 23624 32852 23630 32904
rect 23842 32852 23848 32904
rect 23900 32892 23906 32904
rect 24857 32895 24915 32901
rect 24857 32892 24869 32895
rect 23900 32864 24869 32892
rect 23900 32852 23906 32864
rect 24857 32861 24869 32864
rect 24903 32861 24915 32895
rect 24857 32855 24915 32861
rect 25225 32895 25283 32901
rect 25225 32861 25237 32895
rect 25271 32892 25283 32895
rect 25958 32892 25964 32904
rect 25271 32864 25964 32892
rect 25271 32861 25283 32864
rect 25225 32855 25283 32861
rect 25958 32852 25964 32864
rect 26016 32852 26022 32904
rect 26160 32901 26188 32932
rect 27433 32929 27445 32963
rect 27479 32929 27491 32963
rect 28718 32960 28724 32972
rect 28679 32932 28724 32960
rect 27433 32923 27491 32929
rect 28718 32920 28724 32932
rect 28776 32920 28782 32972
rect 26145 32895 26203 32901
rect 26145 32861 26157 32895
rect 26191 32861 26203 32895
rect 26145 32855 26203 32861
rect 26234 32852 26240 32904
rect 26292 32892 26298 32904
rect 26789 32895 26847 32901
rect 26789 32892 26801 32895
rect 26292 32864 26801 32892
rect 26292 32852 26298 32864
rect 26789 32861 26801 32864
rect 26835 32861 26847 32895
rect 26789 32855 26847 32861
rect 27893 32895 27951 32901
rect 27893 32861 27905 32895
rect 27939 32892 27951 32895
rect 27982 32892 27988 32904
rect 27939 32864 27988 32892
rect 27939 32861 27951 32864
rect 27893 32855 27951 32861
rect 20956 32796 22048 32824
rect 22189 32827 22247 32833
rect 20956 32784 20962 32796
rect 22189 32793 22201 32827
rect 22235 32824 22247 32827
rect 22738 32824 22744 32836
rect 22235 32796 22744 32824
rect 22235 32793 22247 32796
rect 22189 32787 22247 32793
rect 22738 32784 22744 32796
rect 22796 32784 22802 32836
rect 25682 32784 25688 32836
rect 25740 32824 25746 32836
rect 27908 32824 27936 32855
rect 27982 32852 27988 32864
rect 28040 32852 28046 32904
rect 28166 32852 28172 32904
rect 28224 32892 28230 32904
rect 28261 32895 28319 32901
rect 28261 32892 28273 32895
rect 28224 32864 28273 32892
rect 28224 32852 28230 32864
rect 28261 32861 28273 32864
rect 28307 32861 28319 32895
rect 28261 32855 28319 32861
rect 28813 32895 28871 32901
rect 28813 32861 28825 32895
rect 28859 32892 28871 32895
rect 28902 32892 28908 32904
rect 28859 32864 28908 32892
rect 28859 32861 28871 32864
rect 28813 32855 28871 32861
rect 28902 32852 28908 32864
rect 28960 32852 28966 32904
rect 29914 32901 29920 32904
rect 29733 32895 29791 32901
rect 29733 32861 29745 32895
rect 29779 32861 29791 32895
rect 29733 32855 29791 32861
rect 29881 32895 29920 32901
rect 29881 32861 29893 32895
rect 29881 32855 29920 32861
rect 25740 32796 27936 32824
rect 25740 32784 25746 32796
rect 11054 32756 11060 32768
rect 10520 32728 11060 32756
rect 11054 32716 11060 32728
rect 11112 32716 11118 32768
rect 13725 32759 13783 32765
rect 13725 32725 13737 32759
rect 13771 32756 13783 32759
rect 14182 32756 14188 32768
rect 13771 32728 14188 32756
rect 13771 32725 13783 32728
rect 13725 32719 13783 32725
rect 14182 32716 14188 32728
rect 14240 32716 14246 32768
rect 15654 32716 15660 32768
rect 15712 32756 15718 32768
rect 18414 32756 18420 32768
rect 15712 32728 18420 32756
rect 15712 32716 15718 32728
rect 18414 32716 18420 32728
rect 18472 32716 18478 32768
rect 18509 32759 18567 32765
rect 18509 32725 18521 32759
rect 18555 32756 18567 32759
rect 18690 32756 18696 32768
rect 18555 32728 18696 32756
rect 18555 32725 18567 32728
rect 18509 32719 18567 32725
rect 18690 32716 18696 32728
rect 18748 32716 18754 32768
rect 19426 32716 19432 32768
rect 19484 32756 19490 32768
rect 19794 32756 19800 32768
rect 19484 32728 19800 32756
rect 19484 32716 19490 32728
rect 19794 32716 19800 32728
rect 19852 32716 19858 32768
rect 19978 32716 19984 32768
rect 20036 32756 20042 32768
rect 20349 32759 20407 32765
rect 20349 32756 20361 32759
rect 20036 32728 20361 32756
rect 20036 32716 20042 32728
rect 20349 32725 20361 32728
rect 20395 32725 20407 32759
rect 20349 32719 20407 32725
rect 21266 32716 21272 32768
rect 21324 32756 21330 32768
rect 21634 32756 21640 32768
rect 21324 32728 21640 32756
rect 21324 32716 21330 32728
rect 21634 32716 21640 32728
rect 21692 32716 21698 32768
rect 21913 32759 21971 32765
rect 21913 32725 21925 32759
rect 21959 32756 21971 32759
rect 22646 32756 22652 32768
rect 21959 32728 22652 32756
rect 21959 32725 21971 32728
rect 21913 32719 21971 32725
rect 22646 32716 22652 32728
rect 22704 32716 22710 32768
rect 23106 32756 23112 32768
rect 23067 32728 23112 32756
rect 23106 32716 23112 32728
rect 23164 32716 23170 32768
rect 24210 32716 24216 32768
rect 24268 32756 24274 32768
rect 24762 32756 24768 32768
rect 24268 32728 24768 32756
rect 24268 32716 24274 32728
rect 24762 32716 24768 32728
rect 24820 32716 24826 32768
rect 26970 32716 26976 32768
rect 27028 32756 27034 32768
rect 29748 32756 29776 32855
rect 29914 32852 29920 32855
rect 29972 32852 29978 32904
rect 30098 32892 30104 32904
rect 30059 32864 30104 32892
rect 30098 32852 30104 32864
rect 30156 32852 30162 32904
rect 30213 32901 30241 32988
rect 30198 32895 30256 32901
rect 30198 32861 30210 32895
rect 30244 32892 30256 32895
rect 30244 32864 30328 32892
rect 30244 32861 30256 32864
rect 30198 32855 30256 32861
rect 30009 32827 30067 32833
rect 30009 32793 30021 32827
rect 30055 32793 30067 32827
rect 30009 32787 30067 32793
rect 29822 32756 29828 32768
rect 27028 32728 29828 32756
rect 27028 32716 27034 32728
rect 29822 32716 29828 32728
rect 29880 32716 29886 32768
rect 30024 32756 30052 32787
rect 30300 32768 30328 32864
rect 30374 32852 30380 32904
rect 30432 32892 30438 32904
rect 30944 32901 30972 33000
rect 31496 32972 31524 33000
rect 31478 32920 31484 32972
rect 31536 32920 31542 32972
rect 32122 32920 32128 32972
rect 32180 32960 32186 32972
rect 32180 32932 32260 32960
rect 32180 32920 32186 32932
rect 30837 32895 30895 32901
rect 30837 32892 30849 32895
rect 30432 32864 30849 32892
rect 30432 32852 30438 32864
rect 30837 32861 30849 32864
rect 30883 32861 30895 32895
rect 30837 32855 30895 32861
rect 30930 32895 30988 32901
rect 30930 32861 30942 32895
rect 30976 32861 30988 32895
rect 30930 32855 30988 32861
rect 31294 32852 31300 32904
rect 31352 32901 31358 32904
rect 31352 32892 31360 32901
rect 31938 32892 31944 32904
rect 31352 32864 31397 32892
rect 31899 32864 31944 32892
rect 31352 32855 31360 32864
rect 31352 32852 31358 32855
rect 31938 32852 31944 32864
rect 31996 32852 32002 32904
rect 32232 32901 32260 32932
rect 32217 32895 32275 32901
rect 32217 32861 32229 32895
rect 32263 32861 32275 32895
rect 32217 32855 32275 32861
rect 32306 32852 32312 32904
rect 32364 32892 32370 32904
rect 32364 32864 32409 32892
rect 32364 32852 32370 32864
rect 34514 32852 34520 32904
rect 34572 32892 34578 32904
rect 35158 32892 35164 32904
rect 34572 32864 35164 32892
rect 34572 32852 34578 32864
rect 35158 32852 35164 32864
rect 35216 32852 35222 32904
rect 35434 32852 35440 32904
rect 35492 32892 35498 32904
rect 35821 32901 35849 33000
rect 36004 32901 36032 33068
rect 36354 33056 36360 33068
rect 36412 33056 36418 33108
rect 36262 32988 36268 33040
rect 36320 32988 36326 33040
rect 36280 32960 36308 32988
rect 36817 32963 36875 32969
rect 36817 32960 36829 32963
rect 36280 32932 36829 32960
rect 36817 32929 36829 32932
rect 36863 32929 36875 32963
rect 36817 32923 36875 32929
rect 35713 32895 35771 32901
rect 35713 32892 35725 32895
rect 35492 32864 35725 32892
rect 35492 32852 35498 32864
rect 35713 32861 35725 32864
rect 35759 32861 35771 32895
rect 35713 32855 35771 32861
rect 35806 32895 35864 32901
rect 35806 32861 35818 32895
rect 35852 32861 35864 32895
rect 35806 32855 35864 32861
rect 35989 32895 36047 32901
rect 35989 32861 36001 32895
rect 36035 32861 36047 32895
rect 35989 32855 36047 32861
rect 31113 32827 31171 32833
rect 31113 32793 31125 32827
rect 31159 32793 31171 32827
rect 31113 32787 31171 32793
rect 31205 32827 31263 32833
rect 31205 32793 31217 32827
rect 31251 32824 31263 32827
rect 31251 32796 31616 32824
rect 31251 32793 31263 32796
rect 31205 32787 31263 32793
rect 30098 32756 30104 32768
rect 30024 32728 30104 32756
rect 30098 32716 30104 32728
rect 30156 32716 30162 32768
rect 30282 32716 30288 32768
rect 30340 32716 30346 32768
rect 31128 32756 31156 32787
rect 31294 32756 31300 32768
rect 31128 32728 31300 32756
rect 31294 32716 31300 32728
rect 31352 32716 31358 32768
rect 31588 32756 31616 32796
rect 31754 32784 31760 32836
rect 31812 32824 31818 32836
rect 32125 32827 32183 32833
rect 32125 32824 32137 32827
rect 31812 32796 32137 32824
rect 31812 32784 31818 32796
rect 32125 32793 32137 32796
rect 32171 32793 32183 32827
rect 32125 32787 32183 32793
rect 34882 32756 34888 32768
rect 31588 32728 34888 32756
rect 34882 32716 34888 32728
rect 34940 32716 34946 32768
rect 35821 32756 35849 32855
rect 36170 32852 36176 32904
rect 36228 32901 36234 32904
rect 37090 32901 37096 32904
rect 36228 32892 36236 32901
rect 37084 32892 37096 32901
rect 36228 32864 36273 32892
rect 37051 32864 37096 32892
rect 36228 32855 36236 32864
rect 37084 32855 37096 32864
rect 36228 32852 36234 32855
rect 37090 32852 37096 32855
rect 37148 32852 37154 32904
rect 36078 32824 36084 32836
rect 36039 32796 36084 32824
rect 36078 32784 36084 32796
rect 36136 32784 36142 32836
rect 37826 32756 37832 32768
rect 35821 32728 37832 32756
rect 37826 32716 37832 32728
rect 37884 32756 37890 32768
rect 38197 32759 38255 32765
rect 38197 32756 38209 32759
rect 37884 32728 38209 32756
rect 37884 32716 37890 32728
rect 38197 32725 38209 32728
rect 38243 32725 38255 32759
rect 38197 32719 38255 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 9125 32555 9183 32561
rect 9125 32521 9137 32555
rect 9171 32552 9183 32555
rect 9214 32552 9220 32564
rect 9171 32524 9220 32552
rect 9171 32521 9183 32524
rect 9125 32515 9183 32521
rect 9214 32512 9220 32524
rect 9272 32512 9278 32564
rect 9582 32552 9588 32564
rect 9543 32524 9588 32552
rect 9582 32512 9588 32524
rect 9640 32512 9646 32564
rect 10410 32512 10416 32564
rect 10468 32552 10474 32564
rect 12161 32555 12219 32561
rect 12161 32552 12173 32555
rect 10468 32524 12173 32552
rect 10468 32512 10474 32524
rect 12161 32521 12173 32524
rect 12207 32521 12219 32555
rect 12161 32515 12219 32521
rect 13173 32555 13231 32561
rect 13173 32521 13185 32555
rect 13219 32552 13231 32555
rect 13219 32524 14320 32552
rect 13219 32521 13231 32524
rect 13173 32515 13231 32521
rect 4706 32444 4712 32496
rect 4764 32484 4770 32496
rect 6549 32487 6607 32493
rect 6549 32484 6561 32487
rect 4764 32456 6561 32484
rect 4764 32444 4770 32456
rect 4614 32416 4620 32428
rect 4575 32388 4620 32416
rect 4614 32376 4620 32388
rect 4672 32376 4678 32428
rect 5552 32425 5580 32456
rect 6549 32453 6561 32456
rect 6595 32453 6607 32487
rect 6549 32447 6607 32453
rect 7742 32444 7748 32496
rect 7800 32484 7806 32496
rect 8202 32484 8208 32496
rect 7800 32456 8208 32484
rect 7800 32444 7806 32456
rect 8202 32444 8208 32456
rect 8260 32444 8266 32496
rect 8386 32484 8392 32496
rect 8347 32456 8392 32484
rect 8386 32444 8392 32456
rect 8444 32444 8450 32496
rect 11793 32487 11851 32493
rect 9140 32456 9812 32484
rect 5537 32419 5595 32425
rect 5537 32385 5549 32419
rect 5583 32385 5595 32419
rect 5537 32379 5595 32385
rect 5718 32376 5724 32428
rect 5776 32416 5782 32428
rect 5997 32419 6055 32425
rect 5997 32416 6009 32419
rect 5776 32388 6009 32416
rect 5776 32376 5782 32388
rect 5997 32385 6009 32388
rect 6043 32416 6055 32419
rect 6733 32419 6791 32425
rect 6733 32416 6745 32419
rect 6043 32388 6745 32416
rect 6043 32385 6055 32388
rect 5997 32379 6055 32385
rect 6733 32385 6745 32388
rect 6779 32385 6791 32419
rect 6733 32379 6791 32385
rect 6914 32376 6920 32428
rect 6972 32416 6978 32428
rect 9140 32416 9168 32456
rect 6972 32388 9168 32416
rect 6972 32376 6978 32388
rect 9214 32376 9220 32428
rect 9272 32416 9278 32428
rect 9401 32419 9459 32425
rect 9401 32416 9413 32419
rect 9272 32388 9413 32416
rect 9272 32376 9278 32388
rect 9401 32385 9413 32388
rect 9447 32385 9459 32419
rect 9401 32379 9459 32385
rect 9490 32376 9496 32428
rect 9548 32416 9554 32428
rect 9784 32416 9812 32456
rect 11793 32453 11805 32487
rect 11839 32484 11851 32487
rect 11882 32484 11888 32496
rect 11839 32456 11888 32484
rect 11839 32453 11851 32456
rect 11793 32447 11851 32453
rect 11882 32444 11888 32456
rect 11940 32444 11946 32496
rect 11977 32487 12035 32493
rect 11977 32453 11989 32487
rect 12023 32484 12035 32487
rect 12250 32484 12256 32496
rect 12023 32456 12256 32484
rect 12023 32453 12035 32456
rect 11977 32447 12035 32453
rect 12250 32444 12256 32456
rect 12308 32444 12314 32496
rect 14182 32484 14188 32496
rect 14143 32456 14188 32484
rect 14182 32444 14188 32456
rect 14240 32444 14246 32496
rect 14292 32484 14320 32524
rect 14366 32512 14372 32564
rect 14424 32552 14430 32564
rect 14645 32555 14703 32561
rect 14645 32552 14657 32555
rect 14424 32524 14657 32552
rect 14424 32512 14430 32524
rect 14645 32521 14657 32524
rect 14691 32521 14703 32555
rect 14645 32515 14703 32521
rect 16298 32512 16304 32564
rect 16356 32552 16362 32564
rect 20438 32552 20444 32564
rect 16356 32524 20444 32552
rect 16356 32512 16362 32524
rect 20438 32512 20444 32524
rect 20496 32512 20502 32564
rect 20714 32552 20720 32564
rect 20675 32524 20720 32552
rect 20714 32512 20720 32524
rect 20772 32512 20778 32564
rect 20898 32512 20904 32564
rect 20956 32552 20962 32564
rect 20956 32524 21956 32552
rect 20956 32512 20962 32524
rect 16850 32484 16856 32496
rect 14292 32456 16856 32484
rect 16850 32444 16856 32456
rect 16908 32444 16914 32496
rect 19702 32484 19708 32496
rect 16960 32456 19708 32484
rect 9861 32419 9919 32425
rect 9861 32416 9873 32419
rect 9548 32388 9593 32416
rect 9784 32388 9873 32416
rect 9548 32376 9554 32388
rect 9861 32385 9873 32388
rect 9907 32385 9919 32419
rect 9861 32379 9919 32385
rect 4433 32351 4491 32357
rect 4433 32317 4445 32351
rect 4479 32348 4491 32351
rect 4522 32348 4528 32360
rect 4479 32320 4528 32348
rect 4479 32317 4491 32320
rect 4433 32311 4491 32317
rect 4522 32308 4528 32320
rect 4580 32308 4586 32360
rect 5629 32351 5687 32357
rect 5629 32317 5641 32351
rect 5675 32317 5687 32351
rect 5629 32311 5687 32317
rect 4801 32283 4859 32289
rect 4801 32249 4813 32283
rect 4847 32280 4859 32283
rect 5442 32280 5448 32292
rect 4847 32252 5448 32280
rect 4847 32249 4859 32252
rect 4801 32243 4859 32249
rect 5442 32240 5448 32252
rect 5500 32240 5506 32292
rect 5644 32280 5672 32311
rect 6454 32308 6460 32360
rect 6512 32348 6518 32360
rect 9508 32348 9536 32376
rect 6512 32320 9536 32348
rect 9876 32348 9904 32379
rect 10226 32376 10232 32428
rect 10284 32416 10290 32428
rect 10321 32419 10379 32425
rect 10321 32416 10333 32419
rect 10284 32388 10333 32416
rect 10284 32376 10290 32388
rect 10321 32385 10333 32388
rect 10367 32385 10379 32419
rect 10321 32379 10379 32385
rect 12066 32376 12072 32428
rect 12124 32416 12130 32428
rect 12805 32419 12863 32425
rect 12805 32416 12817 32419
rect 12124 32388 12169 32416
rect 12268 32388 12817 32416
rect 12124 32376 12130 32388
rect 10505 32351 10563 32357
rect 10505 32348 10517 32351
rect 9876 32320 10517 32348
rect 6512 32308 6518 32320
rect 10505 32317 10517 32320
rect 10551 32348 10563 32351
rect 11974 32348 11980 32360
rect 10551 32320 11980 32348
rect 10551 32317 10563 32320
rect 10505 32311 10563 32317
rect 11974 32308 11980 32320
rect 12032 32308 12038 32360
rect 12158 32308 12164 32360
rect 12216 32348 12222 32360
rect 12268 32348 12296 32388
rect 12805 32385 12817 32388
rect 12851 32385 12863 32419
rect 12805 32379 12863 32385
rect 14461 32419 14519 32425
rect 14461 32385 14473 32419
rect 14507 32416 14519 32419
rect 14550 32416 14556 32428
rect 14507 32388 14556 32416
rect 14507 32385 14519 32388
rect 14461 32379 14519 32385
rect 14550 32376 14556 32388
rect 14608 32376 14614 32428
rect 14918 32376 14924 32428
rect 14976 32416 14982 32428
rect 15289 32419 15347 32425
rect 15289 32416 15301 32419
rect 14976 32388 15301 32416
rect 14976 32376 14982 32388
rect 15289 32385 15301 32388
rect 15335 32416 15347 32419
rect 16025 32419 16083 32425
rect 15335 32388 15976 32416
rect 15335 32385 15347 32388
rect 15289 32379 15347 32385
rect 12216 32320 12296 32348
rect 12345 32351 12403 32357
rect 12216 32308 12222 32320
rect 12345 32317 12357 32351
rect 12391 32348 12403 32351
rect 12618 32348 12624 32360
rect 12391 32320 12624 32348
rect 12391 32317 12403 32320
rect 12345 32311 12403 32317
rect 12618 32308 12624 32320
rect 12676 32308 12682 32360
rect 12894 32348 12900 32360
rect 12855 32320 12900 32348
rect 12894 32308 12900 32320
rect 12952 32308 12958 32360
rect 14366 32348 14372 32360
rect 14327 32320 14372 32348
rect 14366 32308 14372 32320
rect 14424 32308 14430 32360
rect 14826 32308 14832 32360
rect 14884 32348 14890 32360
rect 15105 32351 15163 32357
rect 15105 32348 15117 32351
rect 14884 32320 15117 32348
rect 14884 32308 14890 32320
rect 15105 32317 15117 32320
rect 15151 32317 15163 32351
rect 15378 32348 15384 32360
rect 15339 32320 15384 32348
rect 15105 32311 15163 32317
rect 15378 32308 15384 32320
rect 15436 32308 15442 32360
rect 15470 32308 15476 32360
rect 15528 32348 15534 32360
rect 15948 32348 15976 32388
rect 16025 32385 16037 32419
rect 16071 32416 16083 32419
rect 16298 32416 16304 32428
rect 16071 32388 16304 32416
rect 16071 32385 16083 32388
rect 16025 32379 16083 32385
rect 16298 32376 16304 32388
rect 16356 32376 16362 32428
rect 16960 32348 16988 32456
rect 19702 32444 19708 32456
rect 19760 32444 19766 32496
rect 20346 32444 20352 32496
rect 20404 32444 20410 32496
rect 20622 32444 20628 32496
rect 20680 32484 20686 32496
rect 21818 32484 21824 32496
rect 20680 32456 21824 32484
rect 20680 32444 20686 32456
rect 17310 32416 17316 32428
rect 17271 32388 17316 32416
rect 17310 32376 17316 32388
rect 17368 32376 17374 32428
rect 17420 32388 17632 32416
rect 15528 32320 15573 32348
rect 15948 32320 16988 32348
rect 17221 32351 17279 32357
rect 15528 32308 15534 32320
rect 17221 32317 17233 32351
rect 17267 32348 17279 32351
rect 17420 32348 17448 32388
rect 17267 32320 17448 32348
rect 17604 32348 17632 32388
rect 17678 32376 17684 32428
rect 17736 32416 17742 32428
rect 17957 32419 18015 32425
rect 17957 32416 17969 32419
rect 17736 32388 17969 32416
rect 17736 32376 17742 32388
rect 17957 32385 17969 32388
rect 18003 32385 18015 32419
rect 18138 32416 18144 32428
rect 18099 32388 18144 32416
rect 17957 32379 18015 32385
rect 18138 32376 18144 32388
rect 18196 32376 18202 32428
rect 20364 32416 20392 32444
rect 20533 32419 20591 32425
rect 20533 32416 20545 32419
rect 20364 32388 20545 32416
rect 20533 32385 20545 32388
rect 20579 32416 20591 32419
rect 20898 32416 20904 32428
rect 20579 32388 20904 32416
rect 20579 32385 20591 32388
rect 20533 32379 20591 32385
rect 20898 32376 20904 32388
rect 20956 32376 20962 32428
rect 21284 32425 21312 32456
rect 21818 32444 21824 32456
rect 21876 32444 21882 32496
rect 21269 32419 21327 32425
rect 21269 32385 21281 32419
rect 21315 32385 21327 32419
rect 21269 32379 21327 32385
rect 21453 32419 21511 32425
rect 21453 32385 21465 32419
rect 21499 32385 21511 32419
rect 21928 32416 21956 32524
rect 22278 32512 22284 32564
rect 22336 32512 22342 32564
rect 25958 32552 25964 32564
rect 25919 32524 25964 32552
rect 25958 32512 25964 32524
rect 26016 32512 26022 32564
rect 30837 32555 30895 32561
rect 30837 32521 30849 32555
rect 30883 32552 30895 32555
rect 31018 32552 31024 32564
rect 30883 32524 31024 32552
rect 30883 32521 30895 32524
rect 30837 32515 30895 32521
rect 31018 32512 31024 32524
rect 31076 32512 31082 32564
rect 32306 32512 32312 32564
rect 32364 32552 32370 32564
rect 34790 32552 34796 32564
rect 32364 32524 34796 32552
rect 32364 32512 32370 32524
rect 34790 32512 34796 32524
rect 34848 32552 34854 32564
rect 35250 32552 35256 32564
rect 34848 32524 35256 32552
rect 34848 32512 34854 32524
rect 35250 32512 35256 32524
rect 35308 32512 35314 32564
rect 35434 32552 35440 32564
rect 35395 32524 35440 32552
rect 35434 32512 35440 32524
rect 35492 32512 35498 32564
rect 22296 32425 22324 32512
rect 26142 32444 26148 32496
rect 26200 32484 26206 32496
rect 27522 32484 27528 32496
rect 26200 32456 27528 32484
rect 26200 32444 26206 32456
rect 22005 32419 22063 32425
rect 22005 32416 22017 32419
rect 21928 32388 22017 32416
rect 21453 32379 21511 32385
rect 22005 32385 22017 32388
rect 22051 32385 22063 32419
rect 22005 32379 22063 32385
rect 22281 32419 22339 32425
rect 22281 32385 22293 32419
rect 22327 32416 22339 32419
rect 22830 32416 22836 32428
rect 22327 32388 22836 32416
rect 22327 32385 22339 32388
rect 22281 32379 22339 32385
rect 19978 32348 19984 32360
rect 17604 32320 19984 32348
rect 17267 32317 17279 32320
rect 17221 32311 17279 32317
rect 19978 32308 19984 32320
rect 20036 32308 20042 32360
rect 20349 32351 20407 32357
rect 20349 32317 20361 32351
rect 20395 32348 20407 32351
rect 21174 32348 21180 32360
rect 20395 32320 21180 32348
rect 20395 32317 20407 32320
rect 20349 32311 20407 32317
rect 21174 32308 21180 32320
rect 21232 32308 21238 32360
rect 21468 32348 21496 32379
rect 22830 32376 22836 32388
rect 22888 32376 22894 32428
rect 23014 32376 23020 32428
rect 23072 32416 23078 32428
rect 23109 32419 23167 32425
rect 23109 32416 23121 32419
rect 23072 32388 23121 32416
rect 23072 32376 23078 32388
rect 23109 32385 23121 32388
rect 23155 32385 23167 32419
rect 23109 32379 23167 32385
rect 23293 32419 23351 32425
rect 23293 32385 23305 32419
rect 23339 32416 23351 32419
rect 24118 32416 24124 32428
rect 23339 32388 24124 32416
rect 23339 32385 23351 32388
rect 23293 32379 23351 32385
rect 24118 32376 24124 32388
rect 24176 32376 24182 32428
rect 24210 32376 24216 32428
rect 24268 32416 24274 32428
rect 24397 32419 24455 32425
rect 24268 32388 24313 32416
rect 24268 32376 24274 32388
rect 24397 32385 24409 32419
rect 24443 32416 24455 32419
rect 25038 32416 25044 32428
rect 24443 32388 25044 32416
rect 24443 32385 24455 32388
rect 24397 32379 24455 32385
rect 25038 32376 25044 32388
rect 25096 32376 25102 32428
rect 25682 32376 25688 32428
rect 25740 32416 25746 32428
rect 25869 32419 25927 32425
rect 25869 32416 25881 32419
rect 25740 32388 25881 32416
rect 25740 32376 25746 32388
rect 25869 32385 25881 32388
rect 25915 32385 25927 32419
rect 25869 32379 25927 32385
rect 26234 32376 26240 32428
rect 26292 32416 26298 32428
rect 27172 32425 27200 32456
rect 27522 32444 27528 32456
rect 27580 32484 27586 32496
rect 27580 32456 28948 32484
rect 27580 32444 27586 32456
rect 26329 32419 26387 32425
rect 26329 32416 26341 32419
rect 26292 32388 26341 32416
rect 26292 32376 26298 32388
rect 26329 32385 26341 32388
rect 26375 32385 26387 32419
rect 26329 32379 26387 32385
rect 27157 32419 27215 32425
rect 27157 32385 27169 32419
rect 27203 32385 27215 32419
rect 27157 32379 27215 32385
rect 27341 32419 27399 32425
rect 27341 32385 27353 32419
rect 27387 32385 27399 32419
rect 28442 32416 28448 32428
rect 28403 32388 28448 32416
rect 27341 32379 27399 32385
rect 21468 32320 22304 32348
rect 6730 32280 6736 32292
rect 5644 32252 6736 32280
rect 6730 32240 6736 32252
rect 6788 32240 6794 32292
rect 8202 32240 8208 32292
rect 8260 32280 8266 32292
rect 8573 32283 8631 32289
rect 8573 32280 8585 32283
rect 8260 32252 8585 32280
rect 8260 32240 8266 32252
rect 8573 32249 8585 32252
rect 8619 32280 8631 32283
rect 10318 32280 10324 32292
rect 8619 32252 10324 32280
rect 8619 32249 8631 32252
rect 8573 32243 8631 32249
rect 10318 32240 10324 32252
rect 10376 32280 10382 32292
rect 10376 32252 11192 32280
rect 10376 32240 10382 32252
rect 6638 32172 6644 32224
rect 6696 32212 6702 32224
rect 6825 32215 6883 32221
rect 6825 32212 6837 32215
rect 6696 32184 6837 32212
rect 6696 32172 6702 32184
rect 6825 32181 6837 32184
rect 6871 32181 6883 32215
rect 6825 32175 6883 32181
rect 8294 32172 8300 32224
rect 8352 32212 8358 32224
rect 9674 32212 9680 32224
rect 8352 32184 9680 32212
rect 8352 32172 8358 32184
rect 9674 32172 9680 32184
rect 9732 32172 9738 32224
rect 9769 32215 9827 32221
rect 9769 32181 9781 32215
rect 9815 32212 9827 32215
rect 11054 32212 11060 32224
rect 9815 32184 11060 32212
rect 9815 32181 9827 32184
rect 9769 32175 9827 32181
rect 11054 32172 11060 32184
rect 11112 32172 11118 32224
rect 11164 32212 11192 32252
rect 11514 32240 11520 32292
rect 11572 32280 11578 32292
rect 11572 32252 13124 32280
rect 11572 32240 11578 32252
rect 12342 32212 12348 32224
rect 11164 32184 12348 32212
rect 12342 32172 12348 32184
rect 12400 32172 12406 32224
rect 12802 32212 12808 32224
rect 12763 32184 12808 32212
rect 12802 32172 12808 32184
rect 12860 32172 12866 32224
rect 13096 32212 13124 32252
rect 14016 32252 14320 32280
rect 14016 32212 14044 32252
rect 14182 32212 14188 32224
rect 13096 32184 14044 32212
rect 14143 32184 14188 32212
rect 14182 32172 14188 32184
rect 14240 32172 14246 32224
rect 14292 32212 14320 32252
rect 18414 32240 18420 32292
rect 18472 32280 18478 32292
rect 21818 32280 21824 32292
rect 18472 32252 21824 32280
rect 18472 32240 18478 32252
rect 21818 32240 21824 32252
rect 21876 32240 21882 32292
rect 15470 32212 15476 32224
rect 14292 32184 15476 32212
rect 15470 32172 15476 32184
rect 15528 32172 15534 32224
rect 16206 32212 16212 32224
rect 16167 32184 16212 32212
rect 16206 32172 16212 32184
rect 16264 32172 16270 32224
rect 16942 32212 16948 32224
rect 16903 32184 16948 32212
rect 16942 32172 16948 32184
rect 17000 32212 17006 32224
rect 17402 32212 17408 32224
rect 17000 32184 17408 32212
rect 17000 32172 17006 32184
rect 17402 32172 17408 32184
rect 17460 32172 17466 32224
rect 17494 32172 17500 32224
rect 17552 32212 17558 32224
rect 18049 32215 18107 32221
rect 17552 32184 17597 32212
rect 17552 32172 17558 32184
rect 18049 32181 18061 32215
rect 18095 32212 18107 32215
rect 18506 32212 18512 32224
rect 18095 32184 18512 32212
rect 18095 32181 18107 32184
rect 18049 32175 18107 32181
rect 18506 32172 18512 32184
rect 18564 32172 18570 32224
rect 18782 32172 18788 32224
rect 18840 32212 18846 32224
rect 21266 32212 21272 32224
rect 18840 32184 21272 32212
rect 18840 32172 18846 32184
rect 21266 32172 21272 32184
rect 21324 32172 21330 32224
rect 22276 32212 22304 32320
rect 22370 32308 22376 32360
rect 22428 32348 22434 32360
rect 24857 32351 24915 32357
rect 22428 32320 22473 32348
rect 22428 32308 22434 32320
rect 24857 32317 24869 32351
rect 24903 32317 24915 32351
rect 27356 32348 27384 32379
rect 28442 32376 28448 32388
rect 28500 32376 28506 32428
rect 28810 32416 28816 32428
rect 28771 32388 28816 32416
rect 28810 32376 28816 32388
rect 28868 32376 28874 32428
rect 28920 32425 28948 32456
rect 30098 32444 30104 32496
rect 30156 32484 30162 32496
rect 30469 32487 30527 32493
rect 30469 32484 30481 32487
rect 30156 32456 30481 32484
rect 30156 32444 30162 32456
rect 30469 32453 30481 32456
rect 30515 32453 30527 32487
rect 30469 32447 30527 32453
rect 30558 32487 30616 32493
rect 30558 32453 30570 32487
rect 30604 32484 30616 32487
rect 31662 32484 31668 32496
rect 30604 32456 31668 32484
rect 30604 32453 30616 32456
rect 30558 32447 30616 32453
rect 31662 32444 31668 32456
rect 31720 32484 31726 32496
rect 34514 32484 34520 32496
rect 31720 32456 34520 32484
rect 31720 32444 31726 32456
rect 34514 32444 34520 32456
rect 34572 32444 34578 32496
rect 34606 32444 34612 32496
rect 34664 32484 34670 32496
rect 35069 32487 35127 32493
rect 35069 32484 35081 32487
rect 34664 32456 35081 32484
rect 34664 32444 34670 32456
rect 35069 32453 35081 32456
rect 35115 32453 35127 32487
rect 35069 32447 35127 32453
rect 35158 32444 35164 32496
rect 35216 32484 35222 32496
rect 35802 32484 35808 32496
rect 35216 32456 35808 32484
rect 35216 32444 35222 32456
rect 35802 32444 35808 32456
rect 35860 32444 35866 32496
rect 28905 32419 28963 32425
rect 28905 32385 28917 32419
rect 28951 32385 28963 32419
rect 28905 32379 28963 32385
rect 29638 32376 29644 32428
rect 29696 32416 29702 32428
rect 30190 32416 30196 32428
rect 29696 32388 30196 32416
rect 29696 32376 29702 32388
rect 30190 32376 30196 32388
rect 30248 32376 30254 32428
rect 30286 32419 30344 32425
rect 30286 32385 30298 32419
rect 30332 32385 30344 32419
rect 30286 32379 30344 32385
rect 28258 32348 28264 32360
rect 27356 32320 28264 32348
rect 24857 32311 24915 32317
rect 23014 32240 23020 32292
rect 23072 32280 23078 32292
rect 24872 32280 24900 32311
rect 28258 32308 28264 32320
rect 28316 32348 28322 32360
rect 28353 32351 28411 32357
rect 28353 32348 28365 32351
rect 28316 32320 28365 32348
rect 28316 32308 28322 32320
rect 28353 32317 28365 32320
rect 28399 32317 28411 32351
rect 28353 32311 28411 32317
rect 29730 32308 29736 32360
rect 29788 32348 29794 32360
rect 30301 32348 30329 32379
rect 30374 32376 30380 32428
rect 30432 32416 30438 32428
rect 30658 32419 30716 32425
rect 30658 32416 30670 32419
rect 30432 32388 30670 32416
rect 30432 32376 30438 32388
rect 30658 32385 30670 32388
rect 30704 32416 30716 32419
rect 31202 32416 31208 32428
rect 30704 32388 31208 32416
rect 30704 32385 30716 32388
rect 30658 32379 30716 32385
rect 31202 32376 31208 32388
rect 31260 32376 31266 32428
rect 32858 32376 32864 32428
rect 32916 32416 32922 32428
rect 33025 32419 33083 32425
rect 33025 32416 33037 32419
rect 32916 32388 33037 32416
rect 32916 32376 32922 32388
rect 33025 32385 33037 32388
rect 33071 32385 33083 32419
rect 34882 32416 34888 32428
rect 34843 32388 34888 32416
rect 33025 32379 33083 32385
rect 34882 32376 34888 32388
rect 34940 32376 34946 32428
rect 35250 32416 35256 32428
rect 35211 32388 35256 32416
rect 35250 32376 35256 32388
rect 35308 32376 35314 32428
rect 37826 32416 37832 32428
rect 37787 32388 37832 32416
rect 37826 32376 37832 32388
rect 37884 32376 37890 32428
rect 32582 32348 32588 32360
rect 29788 32320 32588 32348
rect 29788 32308 29794 32320
rect 32582 32308 32588 32320
rect 32640 32308 32646 32360
rect 32766 32348 32772 32360
rect 32727 32320 32772 32348
rect 32766 32308 32772 32320
rect 32824 32308 32830 32360
rect 34900 32348 34928 32376
rect 35618 32348 35624 32360
rect 34900 32320 35624 32348
rect 35618 32308 35624 32320
rect 35676 32308 35682 32360
rect 38102 32348 38108 32360
rect 38063 32320 38108 32348
rect 38102 32308 38108 32320
rect 38160 32308 38166 32360
rect 28166 32280 28172 32292
rect 23072 32252 28172 32280
rect 23072 32240 23078 32252
rect 28166 32240 28172 32252
rect 28224 32240 28230 32292
rect 28718 32240 28724 32292
rect 28776 32280 28782 32292
rect 32306 32280 32312 32292
rect 28776 32252 32312 32280
rect 28776 32240 28782 32252
rect 32306 32240 32312 32252
rect 32364 32240 32370 32292
rect 35710 32240 35716 32292
rect 35768 32280 35774 32292
rect 36078 32280 36084 32292
rect 35768 32252 36084 32280
rect 35768 32240 35774 32252
rect 36078 32240 36084 32252
rect 36136 32240 36142 32292
rect 23290 32212 23296 32224
rect 22276 32184 23296 32212
rect 23290 32172 23296 32184
rect 23348 32172 23354 32224
rect 23385 32215 23443 32221
rect 23385 32181 23397 32215
rect 23431 32212 23443 32215
rect 25682 32212 25688 32224
rect 23431 32184 25688 32212
rect 23431 32181 23443 32184
rect 23385 32175 23443 32181
rect 25682 32172 25688 32184
rect 25740 32172 25746 32224
rect 27154 32212 27160 32224
rect 27115 32184 27160 32212
rect 27154 32172 27160 32184
rect 27212 32172 27218 32224
rect 27893 32215 27951 32221
rect 27893 32181 27905 32215
rect 27939 32212 27951 32215
rect 31386 32212 31392 32224
rect 27939 32184 31392 32212
rect 27939 32181 27951 32184
rect 27893 32175 27951 32181
rect 31386 32172 31392 32184
rect 31444 32212 31450 32224
rect 31570 32212 31576 32224
rect 31444 32184 31576 32212
rect 31444 32172 31450 32184
rect 31570 32172 31576 32184
rect 31628 32172 31634 32224
rect 34146 32212 34152 32224
rect 34107 32184 34152 32212
rect 34146 32172 34152 32184
rect 34204 32212 34210 32224
rect 36170 32212 36176 32224
rect 34204 32184 36176 32212
rect 34204 32172 34210 32184
rect 36170 32172 36176 32184
rect 36228 32172 36234 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 6454 32008 6460 32020
rect 6415 31980 6460 32008
rect 6454 31968 6460 31980
rect 6512 31968 6518 32020
rect 6546 31968 6552 32020
rect 6604 32008 6610 32020
rect 8294 32008 8300 32020
rect 6604 31980 8300 32008
rect 6604 31968 6610 31980
rect 4249 31943 4307 31949
rect 4249 31909 4261 31943
rect 4295 31940 4307 31943
rect 4890 31940 4896 31952
rect 4295 31912 4896 31940
rect 4295 31909 4307 31912
rect 4249 31903 4307 31909
rect 4890 31900 4896 31912
rect 4948 31900 4954 31952
rect 4706 31872 4712 31884
rect 4264 31844 4712 31872
rect 4264 31813 4292 31844
rect 4706 31832 4712 31844
rect 4764 31872 4770 31884
rect 5534 31872 5540 31884
rect 4764 31844 4936 31872
rect 4764 31832 4770 31844
rect 4908 31813 4936 31844
rect 5092 31844 5540 31872
rect 4065 31807 4123 31813
rect 4065 31773 4077 31807
rect 4111 31804 4123 31807
rect 4249 31807 4307 31813
rect 4111 31776 4200 31804
rect 4111 31773 4123 31776
rect 4065 31767 4123 31773
rect 4172 31736 4200 31776
rect 4249 31773 4261 31807
rect 4295 31773 4307 31807
rect 4801 31807 4859 31813
rect 4801 31804 4813 31807
rect 4249 31767 4307 31773
rect 4356 31776 4813 31804
rect 4356 31736 4384 31776
rect 4801 31773 4813 31776
rect 4847 31773 4859 31807
rect 4908 31807 4971 31813
rect 4908 31776 4925 31807
rect 4801 31767 4859 31773
rect 4913 31773 4925 31776
rect 4959 31773 4971 31807
rect 5092 31798 5120 31844
rect 5534 31832 5540 31844
rect 5592 31832 5598 31884
rect 4913 31767 4971 31773
rect 5000 31770 5120 31798
rect 5353 31807 5411 31813
rect 5353 31773 5365 31807
rect 5399 31804 5411 31807
rect 5626 31804 5632 31816
rect 5399 31776 5632 31804
rect 5399 31773 5411 31776
rect 4172 31708 4384 31736
rect 4816 31736 4844 31767
rect 5000 31736 5028 31770
rect 5353 31767 5411 31773
rect 5626 31764 5632 31776
rect 5684 31804 5690 31816
rect 5810 31804 5816 31816
rect 5684 31776 5816 31804
rect 5684 31764 5690 31776
rect 5810 31764 5816 31776
rect 5868 31764 5874 31816
rect 6656 31813 6684 31980
rect 8294 31968 8300 31980
rect 8352 31968 8358 32020
rect 9217 32011 9275 32017
rect 9217 31977 9229 32011
rect 9263 32008 9275 32011
rect 9858 32008 9864 32020
rect 9263 31980 9864 32008
rect 9263 31977 9275 31980
rect 9217 31971 9275 31977
rect 9858 31968 9864 31980
rect 9916 31968 9922 32020
rect 10134 32008 10140 32020
rect 10095 31980 10140 32008
rect 10134 31968 10140 31980
rect 10192 31968 10198 32020
rect 11514 32008 11520 32020
rect 11475 31980 11520 32008
rect 11514 31968 11520 31980
rect 11572 31968 11578 32020
rect 11716 31980 12296 32008
rect 6822 31940 6828 31952
rect 6783 31912 6828 31940
rect 6822 31900 6828 31912
rect 6880 31900 6886 31952
rect 9585 31875 9643 31881
rect 6748 31844 9352 31872
rect 6748 31816 6776 31844
rect 6641 31807 6699 31813
rect 6641 31773 6653 31807
rect 6687 31773 6699 31807
rect 6641 31767 6699 31773
rect 6730 31764 6736 31816
rect 6788 31804 6794 31816
rect 6917 31807 6975 31813
rect 6788 31776 6833 31804
rect 6788 31764 6794 31776
rect 6917 31773 6929 31807
rect 6963 31804 6975 31807
rect 7006 31804 7012 31816
rect 6963 31776 7012 31804
rect 6963 31773 6975 31776
rect 6917 31767 6975 31773
rect 7006 31764 7012 31776
rect 7064 31764 7070 31816
rect 8036 31813 8064 31844
rect 7929 31807 7987 31813
rect 7929 31804 7941 31807
rect 7116 31776 7941 31804
rect 4816 31708 5028 31736
rect 6638 31628 6644 31680
rect 6696 31668 6702 31680
rect 7116 31668 7144 31776
rect 7929 31773 7941 31776
rect 7975 31773 7987 31807
rect 7929 31767 7987 31773
rect 8021 31807 8079 31813
rect 8021 31773 8033 31807
rect 8067 31773 8079 31807
rect 8202 31804 8208 31816
rect 8163 31776 8208 31804
rect 8021 31767 8079 31773
rect 8202 31764 8208 31776
rect 8260 31764 8266 31816
rect 8294 31764 8300 31816
rect 8352 31804 8358 31816
rect 8352 31776 8397 31804
rect 8352 31764 8358 31776
rect 6696 31640 7144 31668
rect 6696 31628 6702 31640
rect 7650 31628 7656 31680
rect 7708 31668 7714 31680
rect 7745 31671 7803 31677
rect 7745 31668 7757 31671
rect 7708 31640 7757 31668
rect 7708 31628 7714 31640
rect 7745 31637 7757 31640
rect 7791 31637 7803 31671
rect 9324 31668 9352 31844
rect 9585 31841 9597 31875
rect 9631 31872 9643 31875
rect 10042 31872 10048 31884
rect 9631 31844 10048 31872
rect 9631 31841 9643 31844
rect 9585 31835 9643 31841
rect 10042 31832 10048 31844
rect 10100 31832 10106 31884
rect 11716 31872 11744 31980
rect 11974 31940 11980 31952
rect 10796 31844 11744 31872
rect 9401 31807 9459 31813
rect 9401 31773 9413 31807
rect 9447 31773 9459 31807
rect 9401 31767 9459 31773
rect 9677 31807 9735 31813
rect 9677 31773 9689 31807
rect 9723 31804 9735 31807
rect 9766 31804 9772 31816
rect 9723 31776 9772 31804
rect 9723 31773 9735 31776
rect 9677 31767 9735 31773
rect 9416 31736 9444 31767
rect 9766 31764 9772 31776
rect 9824 31764 9830 31816
rect 9950 31764 9956 31816
rect 10008 31804 10014 31816
rect 10226 31804 10232 31816
rect 10008 31776 10232 31804
rect 10008 31764 10014 31776
rect 10226 31764 10232 31776
rect 10284 31804 10290 31816
rect 10321 31807 10379 31813
rect 10321 31804 10333 31807
rect 10284 31776 10333 31804
rect 10284 31764 10290 31776
rect 10321 31773 10333 31776
rect 10367 31773 10379 31807
rect 10594 31804 10600 31816
rect 10555 31776 10600 31804
rect 10321 31767 10379 31773
rect 10594 31764 10600 31776
rect 10652 31764 10658 31816
rect 10796 31736 10824 31844
rect 11716 31816 11744 31844
rect 11808 31912 11980 31940
rect 11698 31804 11704 31816
rect 11611 31776 11704 31804
rect 11698 31764 11704 31776
rect 11756 31764 11762 31816
rect 11808 31813 11836 31912
rect 11974 31900 11980 31912
rect 12032 31900 12038 31952
rect 12268 31872 12296 31980
rect 12342 31968 12348 32020
rect 12400 32008 12406 32020
rect 12529 32011 12587 32017
rect 12529 32008 12541 32011
rect 12400 31980 12541 32008
rect 12400 31968 12406 31980
rect 12529 31977 12541 31980
rect 12575 31977 12587 32011
rect 14918 32008 14924 32020
rect 14879 31980 14924 32008
rect 12529 31971 12587 31977
rect 14918 31968 14924 31980
rect 14976 31968 14982 32020
rect 15102 32008 15108 32020
rect 15063 31980 15108 32008
rect 15102 31968 15108 31980
rect 15160 31968 15166 32020
rect 15194 31968 15200 32020
rect 15252 32008 15258 32020
rect 15565 32011 15623 32017
rect 15565 32008 15577 32011
rect 15252 31980 15577 32008
rect 15252 31968 15258 31980
rect 15565 31977 15577 31980
rect 15611 31977 15623 32011
rect 17402 32008 17408 32020
rect 15565 31971 15623 31977
rect 17144 31980 17408 32008
rect 17144 31940 17172 31980
rect 17402 31968 17408 31980
rect 17460 31968 17466 32020
rect 19613 32011 19671 32017
rect 19613 31977 19625 32011
rect 19659 31977 19671 32011
rect 19613 31971 19671 31977
rect 19797 32011 19855 32017
rect 19797 31977 19809 32011
rect 19843 32008 19855 32011
rect 21726 32008 21732 32020
rect 19843 31980 21732 32008
rect 19843 31977 19855 31980
rect 19797 31971 19855 31977
rect 15488 31912 17172 31940
rect 15488 31872 15516 31912
rect 17218 31900 17224 31952
rect 17276 31940 17282 31952
rect 18877 31943 18935 31949
rect 18877 31940 18889 31943
rect 17276 31912 18889 31940
rect 17276 31900 17282 31912
rect 18877 31909 18889 31912
rect 18923 31909 18935 31943
rect 18877 31903 18935 31909
rect 19058 31900 19064 31952
rect 19116 31940 19122 31952
rect 19628 31940 19656 31971
rect 21726 31968 21732 31980
rect 21784 31968 21790 32020
rect 22830 31968 22836 32020
rect 22888 32008 22894 32020
rect 22888 31980 23520 32008
rect 22888 31968 22894 31980
rect 23382 31940 23388 31952
rect 19116 31912 19564 31940
rect 19628 31912 23388 31940
rect 19116 31900 19122 31912
rect 17494 31872 17500 31884
rect 12268 31844 12572 31872
rect 11793 31807 11851 31813
rect 11793 31773 11805 31807
rect 11839 31773 11851 31807
rect 11793 31767 11851 31773
rect 11977 31807 12035 31813
rect 11977 31773 11989 31807
rect 12023 31773 12035 31807
rect 11977 31767 12035 31773
rect 12069 31807 12127 31813
rect 12069 31773 12081 31807
rect 12115 31798 12127 31807
rect 12342 31804 12348 31816
rect 12176 31798 12348 31804
rect 12115 31776 12348 31798
rect 12115 31773 12204 31776
rect 12069 31770 12204 31773
rect 12069 31767 12127 31770
rect 9416 31708 10824 31736
rect 11146 31696 11152 31748
rect 11204 31736 11210 31748
rect 11514 31736 11520 31748
rect 11204 31708 11520 31736
rect 11204 31696 11210 31708
rect 11514 31696 11520 31708
rect 11572 31736 11578 31748
rect 11992 31736 12020 31767
rect 12342 31764 12348 31776
rect 12400 31764 12406 31816
rect 12544 31813 12572 31844
rect 14660 31844 15516 31872
rect 15580 31844 17500 31872
rect 12529 31807 12587 31813
rect 12529 31773 12541 31807
rect 12575 31773 12587 31807
rect 12529 31767 12587 31773
rect 12618 31764 12624 31816
rect 12676 31804 12682 31816
rect 12894 31804 12900 31816
rect 12676 31776 12721 31804
rect 12820 31776 12900 31804
rect 12676 31764 12682 31776
rect 12820 31736 12848 31776
rect 12894 31764 12900 31776
rect 12952 31764 12958 31816
rect 14660 31813 14688 31844
rect 14645 31807 14703 31813
rect 14645 31773 14657 31807
rect 14691 31773 14703 31807
rect 14826 31804 14832 31816
rect 14739 31776 14832 31804
rect 14645 31767 14703 31773
rect 11572 31708 12848 31736
rect 11572 31696 11578 31708
rect 14550 31696 14556 31748
rect 14608 31736 14614 31748
rect 14752 31736 14780 31776
rect 14826 31764 14832 31776
rect 14884 31764 14890 31816
rect 15580 31813 15608 31844
rect 17494 31832 17500 31844
rect 17552 31832 17558 31884
rect 18782 31872 18788 31884
rect 18524 31844 18788 31872
rect 14921 31807 14979 31813
rect 14921 31773 14933 31807
rect 14967 31804 14979 31807
rect 15565 31807 15623 31813
rect 14967 31776 15516 31804
rect 14967 31773 14979 31776
rect 14921 31767 14979 31773
rect 14608 31708 14780 31736
rect 15488 31736 15516 31776
rect 15565 31773 15577 31807
rect 15611 31773 15623 31807
rect 15565 31767 15623 31773
rect 15657 31807 15715 31813
rect 15657 31773 15669 31807
rect 15703 31804 15715 31807
rect 15746 31804 15752 31816
rect 15703 31776 15752 31804
rect 15703 31773 15715 31776
rect 15657 31767 15715 31773
rect 15672 31736 15700 31767
rect 15746 31764 15752 31776
rect 15804 31764 15810 31816
rect 16942 31804 16948 31816
rect 16903 31776 16948 31804
rect 16942 31764 16948 31776
rect 17000 31764 17006 31816
rect 17310 31804 17316 31816
rect 17271 31776 17316 31804
rect 17310 31764 17316 31776
rect 17368 31764 17374 31816
rect 17405 31807 17463 31813
rect 17405 31773 17417 31807
rect 17451 31804 17463 31807
rect 17954 31804 17960 31816
rect 17451 31776 17960 31804
rect 17451 31773 17463 31776
rect 17405 31767 17463 31773
rect 17954 31764 17960 31776
rect 18012 31804 18018 31816
rect 18414 31804 18420 31816
rect 18012 31776 18420 31804
rect 18012 31764 18018 31776
rect 18414 31764 18420 31776
rect 18472 31764 18478 31816
rect 18524 31813 18552 31844
rect 18782 31832 18788 31844
rect 18840 31832 18846 31884
rect 18966 31832 18972 31884
rect 19024 31872 19030 31884
rect 19536 31872 19564 31912
rect 23382 31900 23388 31912
rect 23440 31900 23446 31952
rect 23492 31940 23520 31980
rect 23658 31968 23664 32020
rect 23716 32008 23722 32020
rect 24118 32008 24124 32020
rect 23716 31980 24124 32008
rect 23716 31968 23722 31980
rect 24118 31968 24124 31980
rect 24176 32008 24182 32020
rect 24765 32011 24823 32017
rect 24765 32008 24777 32011
rect 24176 31980 24777 32008
rect 24176 31968 24182 31980
rect 24765 31977 24777 31980
rect 24811 31977 24823 32011
rect 24765 31971 24823 31977
rect 25314 31968 25320 32020
rect 25372 32008 25378 32020
rect 25777 32011 25835 32017
rect 25777 32008 25789 32011
rect 25372 31980 25789 32008
rect 25372 31968 25378 31980
rect 25777 31977 25789 31980
rect 25823 32008 25835 32011
rect 26878 32008 26884 32020
rect 25823 31980 26884 32008
rect 25823 31977 25835 31980
rect 25777 31971 25835 31977
rect 26878 31968 26884 31980
rect 26936 31968 26942 32020
rect 28442 31968 28448 32020
rect 28500 32008 28506 32020
rect 29733 32011 29791 32017
rect 29733 32008 29745 32011
rect 28500 31980 29745 32008
rect 28500 31968 28506 31980
rect 29733 31977 29745 31980
rect 29779 31977 29791 32011
rect 29733 31971 29791 31977
rect 32769 32011 32827 32017
rect 32769 31977 32781 32011
rect 32815 32008 32827 32011
rect 32858 32008 32864 32020
rect 32815 31980 32864 32008
rect 32815 31977 32827 31980
rect 32769 31971 32827 31977
rect 32858 31968 32864 31980
rect 32916 31968 32922 32020
rect 35897 32011 35955 32017
rect 35897 31977 35909 32011
rect 35943 32008 35955 32011
rect 37826 32008 37832 32020
rect 35943 31980 37832 32008
rect 35943 31977 35955 31980
rect 35897 31971 35955 31977
rect 37826 31968 37832 31980
rect 37884 31968 37890 32020
rect 28810 31940 28816 31952
rect 23492 31912 28816 31940
rect 21637 31875 21695 31881
rect 19024 31844 19472 31872
rect 19536 31844 21312 31872
rect 19024 31832 19030 31844
rect 18509 31807 18567 31813
rect 18509 31773 18521 31807
rect 18555 31773 18567 31807
rect 18690 31804 18696 31816
rect 18651 31776 18696 31804
rect 18509 31767 18567 31773
rect 18690 31764 18696 31776
rect 18748 31764 18754 31816
rect 19444 31813 19472 31844
rect 19429 31807 19487 31813
rect 19429 31773 19441 31807
rect 19475 31773 19487 31807
rect 19429 31767 19487 31773
rect 19613 31807 19671 31813
rect 19613 31773 19625 31807
rect 19659 31773 19671 31807
rect 19613 31767 19671 31773
rect 15488 31708 15700 31736
rect 14608 31696 14614 31708
rect 15838 31696 15844 31748
rect 15896 31736 15902 31748
rect 19628 31736 19656 31767
rect 20438 31764 20444 31816
rect 20496 31804 20502 31816
rect 20714 31804 20720 31816
rect 20496 31776 20720 31804
rect 20496 31764 20502 31776
rect 20714 31764 20720 31776
rect 20772 31764 20778 31816
rect 21284 31813 21312 31844
rect 21637 31841 21649 31875
rect 21683 31872 21695 31875
rect 22462 31872 22468 31884
rect 21683 31844 22468 31872
rect 21683 31841 21695 31844
rect 21637 31835 21695 31841
rect 22462 31832 22468 31844
rect 22520 31832 22526 31884
rect 23198 31872 23204 31884
rect 22940 31844 23204 31872
rect 21269 31807 21327 31813
rect 21269 31773 21281 31807
rect 21315 31804 21327 31807
rect 21315 31776 21404 31804
rect 21315 31773 21327 31776
rect 21269 31767 21327 31773
rect 15896 31708 19656 31736
rect 15896 31696 15902 31708
rect 9858 31668 9864 31680
rect 9324 31640 9864 31668
rect 7745 31631 7803 31637
rect 9858 31628 9864 31640
rect 9916 31668 9922 31680
rect 10505 31671 10563 31677
rect 10505 31668 10517 31671
rect 9916 31640 10517 31668
rect 9916 31628 9922 31640
rect 10505 31637 10517 31640
rect 10551 31637 10563 31671
rect 10505 31631 10563 31637
rect 10594 31628 10600 31680
rect 10652 31668 10658 31680
rect 12618 31668 12624 31680
rect 10652 31640 12624 31668
rect 10652 31628 10658 31640
rect 12618 31628 12624 31640
rect 12676 31628 12682 31680
rect 12802 31628 12808 31680
rect 12860 31668 12866 31680
rect 12897 31671 12955 31677
rect 12897 31668 12909 31671
rect 12860 31640 12909 31668
rect 12860 31628 12866 31640
rect 12897 31637 12909 31640
rect 12943 31637 12955 31671
rect 12897 31631 12955 31637
rect 15010 31628 15016 31680
rect 15068 31668 15074 31680
rect 15933 31671 15991 31677
rect 15933 31668 15945 31671
rect 15068 31640 15945 31668
rect 15068 31628 15074 31640
rect 15933 31637 15945 31640
rect 15979 31637 15991 31671
rect 15933 31631 15991 31637
rect 18966 31628 18972 31680
rect 19024 31668 19030 31680
rect 19334 31668 19340 31680
rect 19024 31640 19340 31668
rect 19024 31628 19030 31640
rect 19334 31628 19340 31640
rect 19392 31628 19398 31680
rect 19978 31628 19984 31680
rect 20036 31668 20042 31680
rect 21269 31671 21327 31677
rect 21269 31668 21281 31671
rect 20036 31640 21281 31668
rect 20036 31628 20042 31640
rect 21269 31637 21281 31640
rect 21315 31637 21327 31671
rect 21376 31668 21404 31776
rect 21542 31764 21548 31816
rect 21600 31804 21606 31816
rect 21910 31804 21916 31816
rect 21600 31776 21916 31804
rect 21600 31764 21606 31776
rect 21910 31764 21916 31776
rect 21968 31764 21974 31816
rect 22940 31813 22968 31844
rect 23198 31832 23204 31844
rect 23256 31832 23262 31884
rect 23290 31832 23296 31884
rect 23348 31872 23354 31884
rect 25498 31872 25504 31884
rect 23348 31844 25504 31872
rect 23348 31832 23354 31844
rect 25498 31832 25504 31844
rect 25556 31872 25562 31884
rect 26697 31875 26755 31881
rect 25556 31844 26464 31872
rect 25556 31832 25562 31844
rect 22925 31807 22983 31813
rect 22925 31773 22937 31807
rect 22971 31773 22983 31807
rect 23474 31804 23480 31816
rect 22925 31767 22983 31773
rect 23400 31776 23480 31804
rect 21726 31696 21732 31748
rect 21784 31736 21790 31748
rect 22370 31736 22376 31748
rect 21784 31708 22376 31736
rect 21784 31696 21790 31708
rect 22370 31696 22376 31708
rect 22428 31696 22434 31748
rect 22554 31696 22560 31748
rect 22612 31736 22618 31748
rect 23293 31739 23351 31745
rect 23293 31736 23305 31739
rect 22612 31708 23305 31736
rect 22612 31696 22618 31708
rect 23293 31705 23305 31708
rect 23339 31705 23351 31739
rect 23293 31699 23351 31705
rect 23400 31668 23428 31776
rect 23474 31764 23480 31776
rect 23532 31804 23538 31816
rect 24673 31807 24731 31813
rect 23532 31776 24624 31804
rect 23532 31764 23538 31776
rect 24596 31736 24624 31776
rect 24673 31773 24685 31807
rect 24719 31804 24731 31807
rect 24854 31804 24860 31816
rect 24719 31776 24860 31804
rect 24719 31773 24731 31776
rect 24673 31767 24731 31773
rect 24854 31764 24860 31776
rect 24912 31764 24918 31816
rect 24949 31807 25007 31813
rect 24949 31773 24961 31807
rect 24995 31804 25007 31807
rect 25590 31804 25596 31816
rect 24995 31776 25029 31804
rect 25551 31776 25596 31804
rect 24995 31773 25007 31776
rect 24949 31767 25007 31773
rect 24964 31736 24992 31767
rect 25590 31764 25596 31776
rect 25648 31764 25654 31816
rect 25774 31804 25780 31816
rect 25735 31776 25780 31804
rect 25774 31764 25780 31776
rect 25832 31764 25838 31816
rect 26436 31804 26464 31844
rect 26697 31841 26709 31875
rect 26743 31872 26755 31875
rect 26743 31844 27016 31872
rect 26743 31841 26755 31844
rect 26697 31835 26755 31841
rect 26878 31804 26884 31816
rect 26436 31776 26556 31804
rect 26839 31776 26884 31804
rect 24596 31708 24992 31736
rect 25406 31696 25412 31748
rect 25464 31736 25470 31748
rect 26234 31736 26240 31748
rect 25464 31708 26240 31736
rect 25464 31696 25470 31708
rect 26234 31696 26240 31708
rect 26292 31736 26298 31748
rect 26418 31736 26424 31748
rect 26292 31708 26424 31736
rect 26292 31696 26298 31708
rect 26418 31696 26424 31708
rect 26476 31696 26482 31748
rect 21376 31640 23428 31668
rect 21269 31631 21327 31637
rect 25038 31628 25044 31680
rect 25096 31668 25102 31680
rect 25866 31668 25872 31680
rect 25096 31640 25872 31668
rect 25096 31628 25102 31640
rect 25866 31628 25872 31640
rect 25924 31628 25930 31680
rect 25961 31671 26019 31677
rect 25961 31637 25973 31671
rect 26007 31668 26019 31671
rect 26050 31668 26056 31680
rect 26007 31640 26056 31668
rect 26007 31637 26019 31640
rect 25961 31631 26019 31637
rect 26050 31628 26056 31640
rect 26108 31628 26114 31680
rect 26528 31668 26556 31776
rect 26878 31764 26884 31776
rect 26936 31764 26942 31816
rect 26988 31804 27016 31844
rect 27522 31832 27528 31884
rect 27580 31872 27586 31884
rect 27617 31875 27675 31881
rect 27617 31872 27629 31875
rect 27580 31844 27629 31872
rect 27580 31832 27586 31844
rect 27617 31841 27629 31844
rect 27663 31841 27675 31875
rect 27617 31835 27675 31841
rect 27706 31804 27712 31816
rect 26988 31776 27712 31804
rect 27706 31764 27712 31776
rect 27764 31764 27770 31816
rect 28184 31813 28212 31912
rect 28810 31900 28816 31912
rect 28868 31900 28874 31952
rect 28994 31940 29000 31952
rect 28955 31912 29000 31940
rect 28994 31900 29000 31912
rect 29052 31900 29058 31952
rect 32033 31943 32091 31949
rect 32033 31909 32045 31943
rect 32079 31909 32091 31943
rect 32033 31903 32091 31909
rect 28258 31832 28264 31884
rect 28316 31872 28322 31884
rect 32048 31872 32076 31903
rect 35710 31900 35716 31952
rect 35768 31900 35774 31952
rect 35728 31872 35756 31900
rect 28316 31844 28382 31872
rect 29012 31844 29960 31872
rect 32048 31844 32812 31872
rect 28316 31832 28322 31844
rect 28169 31807 28227 31813
rect 28169 31773 28181 31807
rect 28215 31773 28227 31807
rect 28169 31767 28227 31773
rect 28629 31807 28687 31813
rect 28629 31773 28641 31807
rect 28675 31773 28687 31807
rect 29012 31804 29040 31844
rect 28629 31767 28687 31773
rect 28966 31776 29040 31804
rect 26786 31696 26792 31748
rect 26844 31736 26850 31748
rect 28644 31736 28672 31767
rect 28966 31748 28994 31776
rect 29086 31764 29092 31816
rect 29144 31804 29150 31816
rect 29932 31813 29960 31844
rect 29733 31807 29791 31813
rect 29733 31804 29745 31807
rect 29144 31776 29745 31804
rect 29144 31764 29150 31776
rect 29733 31773 29745 31776
rect 29779 31773 29791 31807
rect 29733 31767 29791 31773
rect 29917 31807 29975 31813
rect 29917 31773 29929 31807
rect 29963 31773 29975 31807
rect 32217 31807 32275 31813
rect 32217 31804 32229 31807
rect 29917 31767 29975 31773
rect 32140 31776 32229 31804
rect 26844 31708 28672 31736
rect 26844 31696 26850 31708
rect 28902 31696 28908 31748
rect 28960 31708 28994 31748
rect 32030 31736 32036 31748
rect 31991 31708 32036 31736
rect 28960 31696 28966 31708
rect 32030 31696 32036 31708
rect 32088 31696 32094 31748
rect 32140 31680 32168 31776
rect 32217 31773 32229 31776
rect 32263 31773 32275 31807
rect 32217 31767 32275 31773
rect 32309 31807 32367 31813
rect 32309 31773 32321 31807
rect 32355 31804 32367 31807
rect 32490 31804 32496 31816
rect 32355 31776 32496 31804
rect 32355 31773 32367 31776
rect 32309 31767 32367 31773
rect 32490 31764 32496 31776
rect 32548 31764 32554 31816
rect 32784 31813 32812 31844
rect 35544 31844 35756 31872
rect 32769 31807 32827 31813
rect 32769 31773 32781 31807
rect 32815 31773 32827 31807
rect 32950 31804 32956 31816
rect 32911 31776 32956 31804
rect 32769 31767 32827 31773
rect 32950 31764 32956 31776
rect 33008 31764 33014 31816
rect 35250 31804 35256 31816
rect 35211 31776 35256 31804
rect 35250 31764 35256 31776
rect 35308 31764 35314 31816
rect 35346 31807 35404 31813
rect 35346 31773 35358 31807
rect 35392 31773 35404 31807
rect 35346 31767 35404 31773
rect 32582 31696 32588 31748
rect 32640 31736 32646 31748
rect 35361 31736 35389 31767
rect 35434 31764 35440 31816
rect 35492 31764 35498 31816
rect 35544 31813 35572 31844
rect 36262 31832 36268 31884
rect 36320 31872 36326 31884
rect 36357 31875 36415 31881
rect 36357 31872 36369 31875
rect 36320 31844 36369 31872
rect 36320 31832 36326 31844
rect 36357 31841 36369 31844
rect 36403 31841 36415 31875
rect 36357 31835 36415 31841
rect 35529 31807 35587 31813
rect 35529 31773 35541 31807
rect 35575 31773 35587 31807
rect 35529 31767 35587 31773
rect 35621 31807 35679 31813
rect 35621 31773 35633 31807
rect 35667 31804 35679 31807
rect 35759 31807 35817 31813
rect 35667 31776 35701 31804
rect 35667 31773 35679 31776
rect 35621 31767 35679 31773
rect 35759 31773 35771 31807
rect 35805 31804 35817 31807
rect 35894 31804 35900 31816
rect 35805 31776 35900 31804
rect 35805 31773 35817 31776
rect 35759 31767 35817 31773
rect 32640 31708 35389 31736
rect 35452 31736 35480 31764
rect 35636 31736 35664 31767
rect 35894 31764 35900 31776
rect 35952 31764 35958 31816
rect 36624 31807 36682 31813
rect 36624 31773 36636 31807
rect 36670 31804 36682 31807
rect 37458 31804 37464 31816
rect 36670 31776 37464 31804
rect 36670 31773 36682 31776
rect 36624 31767 36682 31773
rect 37458 31764 37464 31776
rect 37516 31764 37522 31816
rect 35452 31708 35664 31736
rect 32640 31696 32646 31708
rect 27065 31671 27123 31677
rect 27065 31668 27077 31671
rect 26528 31640 27077 31668
rect 27065 31637 27077 31640
rect 27111 31668 27123 31671
rect 28626 31668 28632 31680
rect 27111 31640 28632 31668
rect 27111 31637 27123 31640
rect 27065 31631 27123 31637
rect 28626 31628 28632 31640
rect 28684 31628 28690 31680
rect 32122 31628 32128 31680
rect 32180 31628 32186 31680
rect 35361 31668 35389 31708
rect 37734 31668 37740 31680
rect 35361 31640 37740 31668
rect 37734 31628 37740 31640
rect 37792 31628 37798 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 7193 31467 7251 31473
rect 7193 31433 7205 31467
rect 7239 31464 7251 31467
rect 11882 31464 11888 31476
rect 7239 31436 11888 31464
rect 7239 31433 7251 31436
rect 7193 31427 7251 31433
rect 11882 31424 11888 31436
rect 11940 31424 11946 31476
rect 12161 31467 12219 31473
rect 12161 31433 12173 31467
rect 12207 31464 12219 31467
rect 12805 31467 12863 31473
rect 12805 31464 12817 31467
rect 12207 31436 12817 31464
rect 12207 31433 12219 31436
rect 12161 31427 12219 31433
rect 12805 31433 12817 31436
rect 12851 31433 12863 31467
rect 12805 31427 12863 31433
rect 12894 31424 12900 31476
rect 12952 31464 12958 31476
rect 14737 31467 14795 31473
rect 12952 31436 14688 31464
rect 12952 31424 12958 31436
rect 7834 31396 7840 31408
rect 7392 31368 7840 31396
rect 5353 31331 5411 31337
rect 5353 31297 5365 31331
rect 5399 31328 5411 31331
rect 5442 31328 5448 31340
rect 5399 31300 5448 31328
rect 5399 31297 5411 31300
rect 5353 31291 5411 31297
rect 5442 31288 5448 31300
rect 5500 31288 5506 31340
rect 5534 31288 5540 31340
rect 5592 31328 5598 31340
rect 6638 31328 6644 31340
rect 5592 31300 6644 31328
rect 5592 31288 5598 31300
rect 6638 31288 6644 31300
rect 6696 31288 6702 31340
rect 7392 31337 7420 31368
rect 7834 31356 7840 31368
rect 7892 31356 7898 31408
rect 8205 31399 8263 31405
rect 8205 31365 8217 31399
rect 8251 31396 8263 31399
rect 9122 31396 9128 31408
rect 8251 31368 9128 31396
rect 8251 31365 8263 31368
rect 8205 31359 8263 31365
rect 9122 31356 9128 31368
rect 9180 31396 9186 31408
rect 13630 31396 13636 31408
rect 9180 31368 13636 31396
rect 9180 31356 9186 31368
rect 13630 31356 13636 31368
rect 13688 31356 13694 31408
rect 14001 31399 14059 31405
rect 14001 31365 14013 31399
rect 14047 31396 14059 31399
rect 14047 31368 14596 31396
rect 14047 31365 14059 31368
rect 14001 31359 14059 31365
rect 14568 31340 14596 31368
rect 7377 31331 7435 31337
rect 7377 31297 7389 31331
rect 7423 31297 7435 31331
rect 7650 31328 7656 31340
rect 7611 31300 7656 31328
rect 7377 31291 7435 31297
rect 7650 31288 7656 31300
rect 7708 31288 7714 31340
rect 10137 31331 10195 31337
rect 10137 31297 10149 31331
rect 10183 31328 10195 31331
rect 10318 31328 10324 31340
rect 10183 31300 10324 31328
rect 10183 31297 10195 31300
rect 10137 31291 10195 31297
rect 10318 31288 10324 31300
rect 10376 31288 10382 31340
rect 10413 31331 10471 31337
rect 10413 31297 10425 31331
rect 10459 31328 10471 31331
rect 10594 31328 10600 31340
rect 10459 31300 10600 31328
rect 10459 31297 10471 31300
rect 10413 31291 10471 31297
rect 10594 31288 10600 31300
rect 10652 31288 10658 31340
rect 11790 31328 11796 31340
rect 11751 31300 11796 31328
rect 11790 31288 11796 31300
rect 11848 31288 11854 31340
rect 11977 31331 12035 31337
rect 11977 31297 11989 31331
rect 12023 31328 12035 31331
rect 12342 31328 12348 31340
rect 12023 31300 12348 31328
rect 12023 31297 12035 31300
rect 11977 31291 12035 31297
rect 7469 31263 7527 31269
rect 7469 31229 7481 31263
rect 7515 31260 7527 31263
rect 8202 31260 8208 31272
rect 7515 31232 8208 31260
rect 7515 31229 7527 31232
rect 7469 31223 7527 31229
rect 8202 31220 8208 31232
rect 8260 31220 8266 31272
rect 9033 31263 9091 31269
rect 9033 31229 9045 31263
rect 9079 31260 9091 31263
rect 9582 31260 9588 31272
rect 9079 31232 9588 31260
rect 9079 31229 9091 31232
rect 9033 31223 9091 31229
rect 9582 31220 9588 31232
rect 9640 31220 9646 31272
rect 10229 31263 10287 31269
rect 10229 31229 10241 31263
rect 10275 31229 10287 31263
rect 10229 31223 10287 31229
rect 7561 31195 7619 31201
rect 7561 31161 7573 31195
rect 7607 31192 7619 31195
rect 7926 31192 7932 31204
rect 7607 31164 7932 31192
rect 7607 31161 7619 31164
rect 7561 31155 7619 31161
rect 7926 31152 7932 31164
rect 7984 31152 7990 31204
rect 10244 31192 10272 31223
rect 11054 31220 11060 31272
rect 11112 31260 11118 31272
rect 11992 31260 12020 31291
rect 12342 31288 12348 31300
rect 12400 31288 12406 31340
rect 12434 31288 12440 31340
rect 12492 31328 12498 31340
rect 12621 31331 12679 31337
rect 12621 31328 12633 31331
rect 12492 31300 12633 31328
rect 12492 31288 12498 31300
rect 12621 31297 12633 31300
rect 12667 31297 12679 31331
rect 12621 31291 12679 31297
rect 12897 31331 12955 31337
rect 12897 31297 12909 31331
rect 12943 31297 12955 31331
rect 12897 31291 12955 31297
rect 11112 31232 12020 31260
rect 11112 31220 11118 31232
rect 12250 31220 12256 31272
rect 12308 31260 12314 31272
rect 12912 31260 12940 31291
rect 12986 31288 12992 31340
rect 13044 31328 13050 31340
rect 14277 31331 14335 31337
rect 14277 31328 14289 31331
rect 13044 31300 14289 31328
rect 13044 31288 13050 31300
rect 14277 31297 14289 31300
rect 14323 31297 14335 31331
rect 14550 31328 14556 31340
rect 14511 31300 14556 31328
rect 14277 31291 14335 31297
rect 14550 31288 14556 31300
rect 14608 31288 14614 31340
rect 14660 31328 14688 31436
rect 14737 31433 14749 31467
rect 14783 31464 14795 31467
rect 15378 31464 15384 31476
rect 14783 31436 15384 31464
rect 14783 31433 14795 31436
rect 14737 31427 14795 31433
rect 15378 31424 15384 31436
rect 15436 31424 15442 31476
rect 17402 31424 17408 31476
rect 17460 31464 17466 31476
rect 17497 31467 17555 31473
rect 17497 31464 17509 31467
rect 17460 31436 17509 31464
rect 17460 31424 17466 31436
rect 17497 31433 17509 31436
rect 17543 31433 17555 31467
rect 18874 31464 18880 31476
rect 18835 31436 18880 31464
rect 17497 31427 17555 31433
rect 18874 31424 18880 31436
rect 18932 31424 18938 31476
rect 19978 31464 19984 31476
rect 18984 31436 19984 31464
rect 16850 31396 16856 31408
rect 16811 31368 16856 31396
rect 16850 31356 16856 31368
rect 16908 31356 16914 31408
rect 16942 31356 16948 31408
rect 17000 31396 17006 31408
rect 18984 31396 19012 31436
rect 19978 31424 19984 31436
rect 20036 31424 20042 31476
rect 22002 31424 22008 31476
rect 22060 31464 22066 31476
rect 22281 31467 22339 31473
rect 22281 31464 22293 31467
rect 22060 31436 22293 31464
rect 22060 31424 22066 31436
rect 22281 31433 22293 31436
rect 22327 31433 22339 31467
rect 22281 31427 22339 31433
rect 23566 31424 23572 31476
rect 23624 31464 23630 31476
rect 25590 31464 25596 31476
rect 23624 31436 25596 31464
rect 23624 31424 23630 31436
rect 25590 31424 25596 31436
rect 25648 31464 25654 31476
rect 27430 31464 27436 31476
rect 25648 31436 27436 31464
rect 25648 31424 25654 31436
rect 27430 31424 27436 31436
rect 27488 31464 27494 31476
rect 27890 31464 27896 31476
rect 27488 31436 27896 31464
rect 27488 31424 27494 31436
rect 27890 31424 27896 31436
rect 27948 31424 27954 31476
rect 28258 31424 28264 31476
rect 28316 31464 28322 31476
rect 28629 31467 28687 31473
rect 28629 31464 28641 31467
rect 28316 31436 28641 31464
rect 28316 31424 28322 31436
rect 28629 31433 28641 31436
rect 28675 31433 28687 31467
rect 28629 31427 28687 31433
rect 30742 31424 30748 31476
rect 30800 31464 30806 31476
rect 31297 31467 31355 31473
rect 30800 31436 31248 31464
rect 30800 31424 30806 31436
rect 17000 31368 19012 31396
rect 17000 31356 17006 31368
rect 15289 31331 15347 31337
rect 15289 31328 15301 31331
rect 14660 31300 15301 31328
rect 15289 31297 15301 31300
rect 15335 31328 15347 31331
rect 16206 31328 16212 31340
rect 15335 31300 16212 31328
rect 15335 31297 15347 31300
rect 15289 31291 15347 31297
rect 16206 31288 16212 31300
rect 16264 31288 16270 31340
rect 17328 31337 17356 31368
rect 19150 31356 19156 31408
rect 19208 31396 19214 31408
rect 19518 31396 19524 31408
rect 19208 31368 19524 31396
rect 19208 31356 19214 31368
rect 19518 31356 19524 31368
rect 19576 31396 19582 31408
rect 19576 31368 20484 31396
rect 19576 31356 19582 31368
rect 17313 31331 17371 31337
rect 17313 31297 17325 31331
rect 17359 31297 17371 31331
rect 17313 31291 17371 31297
rect 18233 31331 18291 31337
rect 18233 31297 18245 31331
rect 18279 31297 18291 31331
rect 18506 31328 18512 31340
rect 18467 31300 18512 31328
rect 18233 31291 18291 31297
rect 14461 31263 14519 31269
rect 12308 31232 12940 31260
rect 13740 31232 14412 31260
rect 12308 31220 12314 31232
rect 11882 31192 11888 31204
rect 10244 31164 11888 31192
rect 11882 31152 11888 31164
rect 11940 31152 11946 31204
rect 12621 31195 12679 31201
rect 12621 31161 12633 31195
rect 12667 31192 12679 31195
rect 13740 31192 13768 31232
rect 12667 31164 13768 31192
rect 12667 31161 12679 31164
rect 12621 31155 12679 31161
rect 13814 31152 13820 31204
rect 13872 31192 13878 31204
rect 14384 31192 14412 31232
rect 14461 31229 14473 31263
rect 14507 31260 14519 31263
rect 15378 31260 15384 31272
rect 14507 31232 15384 31260
rect 14507 31229 14519 31232
rect 14461 31223 14519 31229
rect 15378 31220 15384 31232
rect 15436 31220 15442 31272
rect 15470 31220 15476 31272
rect 15528 31260 15534 31272
rect 17218 31260 17224 31272
rect 15528 31232 15573 31260
rect 17131 31232 17224 31260
rect 15528 31220 15534 31232
rect 17218 31220 17224 31232
rect 17276 31260 17282 31272
rect 17402 31260 17408 31272
rect 17276 31232 17408 31260
rect 17276 31220 17282 31232
rect 17402 31220 17408 31232
rect 17460 31220 17466 31272
rect 18248 31260 18276 31291
rect 18506 31288 18512 31300
rect 18564 31288 18570 31340
rect 18693 31331 18751 31337
rect 18693 31297 18705 31331
rect 18739 31328 18751 31331
rect 18782 31328 18788 31340
rect 18739 31300 18788 31328
rect 18739 31297 18751 31300
rect 18693 31291 18751 31297
rect 18782 31288 18788 31300
rect 18840 31288 18846 31340
rect 18966 31288 18972 31340
rect 19024 31328 19030 31340
rect 19613 31331 19671 31337
rect 19613 31328 19625 31331
rect 19024 31300 19625 31328
rect 19024 31288 19030 31300
rect 19613 31297 19625 31300
rect 19659 31297 19671 31331
rect 19613 31291 19671 31297
rect 19705 31331 19763 31337
rect 19705 31297 19717 31331
rect 19751 31328 19763 31331
rect 20254 31328 20260 31340
rect 19751 31300 20260 31328
rect 19751 31297 19763 31300
rect 19705 31291 19763 31297
rect 20254 31288 20260 31300
rect 20312 31288 20318 31340
rect 20456 31337 20484 31368
rect 21284 31368 22324 31396
rect 21284 31337 21312 31368
rect 22296 31340 22324 31368
rect 22370 31356 22376 31408
rect 22428 31396 22434 31408
rect 28994 31396 29000 31408
rect 22428 31368 26280 31396
rect 22428 31356 22434 31368
rect 20441 31331 20499 31337
rect 20441 31297 20453 31331
rect 20487 31297 20499 31331
rect 20441 31291 20499 31297
rect 21269 31331 21327 31337
rect 21269 31297 21281 31331
rect 21315 31297 21327 31331
rect 21450 31328 21456 31340
rect 21411 31300 21456 31328
rect 21269 31291 21327 31297
rect 21450 31288 21456 31300
rect 21508 31288 21514 31340
rect 22278 31328 22284 31340
rect 22239 31300 22284 31328
rect 22278 31288 22284 31300
rect 22336 31288 22342 31340
rect 22572 31337 22600 31368
rect 22557 31331 22615 31337
rect 22557 31297 22569 31331
rect 22603 31297 22615 31331
rect 23658 31328 23664 31340
rect 23619 31300 23664 31328
rect 22557 31291 22615 31297
rect 23658 31288 23664 31300
rect 23716 31288 23722 31340
rect 23750 31288 23756 31340
rect 23808 31328 23814 31340
rect 23937 31331 23995 31337
rect 23937 31328 23949 31331
rect 23808 31300 23949 31328
rect 23808 31288 23814 31300
rect 23937 31297 23949 31300
rect 23983 31297 23995 31331
rect 25406 31328 25412 31340
rect 23937 31291 23995 31297
rect 24320 31300 25412 31328
rect 19429 31263 19487 31269
rect 19429 31260 19441 31263
rect 18248 31232 19441 31260
rect 19429 31229 19441 31232
rect 19475 31229 19487 31263
rect 19429 31223 19487 31229
rect 19797 31263 19855 31269
rect 19797 31229 19809 31263
rect 19843 31229 19855 31263
rect 19797 31223 19855 31229
rect 15838 31192 15844 31204
rect 13872 31164 14320 31192
rect 14384 31164 15844 31192
rect 13872 31152 13878 31164
rect 5534 31084 5540 31136
rect 5592 31124 5598 31136
rect 5629 31127 5687 31133
rect 5629 31124 5641 31127
rect 5592 31096 5641 31124
rect 5592 31084 5598 31096
rect 5629 31093 5641 31096
rect 5675 31093 5687 31127
rect 5629 31087 5687 31093
rect 6086 31084 6092 31136
rect 6144 31124 6150 31136
rect 9766 31124 9772 31136
rect 6144 31096 9772 31124
rect 6144 31084 6150 31096
rect 9766 31084 9772 31096
rect 9824 31124 9830 31136
rect 10413 31127 10471 31133
rect 10413 31124 10425 31127
rect 9824 31096 10425 31124
rect 9824 31084 9830 31096
rect 10413 31093 10425 31096
rect 10459 31124 10471 31127
rect 10502 31124 10508 31136
rect 10459 31096 10508 31124
rect 10459 31093 10471 31096
rect 10413 31087 10471 31093
rect 10502 31084 10508 31096
rect 10560 31084 10566 31136
rect 10597 31127 10655 31133
rect 10597 31093 10609 31127
rect 10643 31124 10655 31127
rect 11698 31124 11704 31136
rect 10643 31096 11704 31124
rect 10643 31093 10655 31096
rect 10597 31087 10655 31093
rect 11698 31084 11704 31096
rect 11756 31084 11762 31136
rect 14292 31133 14320 31164
rect 15838 31152 15844 31164
rect 15896 31152 15902 31204
rect 17586 31192 17592 31204
rect 17328 31164 17592 31192
rect 17328 31133 17356 31164
rect 17586 31152 17592 31164
rect 17644 31152 17650 31204
rect 19812 31192 19840 31223
rect 19886 31220 19892 31272
rect 19944 31260 19950 31272
rect 20717 31263 20775 31269
rect 19944 31232 19989 31260
rect 19944 31220 19950 31232
rect 20717 31229 20729 31263
rect 20763 31260 20775 31263
rect 21542 31260 21548 31272
rect 20763 31232 21548 31260
rect 20763 31229 20775 31232
rect 20717 31223 20775 31229
rect 21542 31220 21548 31232
rect 21600 31220 21606 31272
rect 24320 31260 24348 31300
rect 25406 31288 25412 31300
rect 25464 31288 25470 31340
rect 25590 31288 25596 31340
rect 25648 31328 25654 31340
rect 25685 31331 25743 31337
rect 25685 31328 25697 31331
rect 25648 31300 25697 31328
rect 25648 31288 25654 31300
rect 25685 31297 25697 31300
rect 25731 31297 25743 31331
rect 25685 31291 25743 31297
rect 25777 31331 25835 31337
rect 25777 31297 25789 31331
rect 25823 31297 25835 31331
rect 25777 31291 25835 31297
rect 22066 31232 24348 31260
rect 24397 31263 24455 31269
rect 20162 31192 20168 31204
rect 19812 31164 20168 31192
rect 20162 31152 20168 31164
rect 20220 31192 20226 31204
rect 22066 31192 22094 31232
rect 24397 31229 24409 31263
rect 24443 31229 24455 31263
rect 24397 31223 24455 31229
rect 20220 31164 22094 31192
rect 20220 31152 20226 31164
rect 23474 31152 23480 31204
rect 23532 31192 23538 31204
rect 23753 31195 23811 31201
rect 23753 31192 23765 31195
rect 23532 31164 23765 31192
rect 23532 31152 23538 31164
rect 23753 31161 23765 31164
rect 23799 31161 23811 31195
rect 23753 31155 23811 31161
rect 24302 31152 24308 31204
rect 24360 31192 24366 31204
rect 24412 31192 24440 31223
rect 25222 31220 25228 31272
rect 25280 31260 25286 31272
rect 25792 31260 25820 31291
rect 25866 31288 25872 31340
rect 25924 31328 25930 31340
rect 26029 31331 26087 31337
rect 25924 31300 25969 31328
rect 25924 31288 25930 31300
rect 26029 31297 26041 31331
rect 26075 31328 26087 31331
rect 26252 31328 26280 31368
rect 28966 31356 29000 31396
rect 29052 31356 29058 31408
rect 30558 31356 30564 31408
rect 30616 31396 30622 31408
rect 31021 31399 31079 31405
rect 31021 31396 31033 31399
rect 30616 31368 31033 31396
rect 30616 31356 30622 31368
rect 31021 31365 31033 31368
rect 31067 31365 31079 31399
rect 31220 31396 31248 31436
rect 31297 31433 31309 31467
rect 31343 31464 31355 31467
rect 32030 31464 32036 31476
rect 31343 31436 32036 31464
rect 31343 31433 31355 31436
rect 31297 31427 31355 31433
rect 32030 31424 32036 31436
rect 32088 31464 32094 31476
rect 32493 31467 32551 31473
rect 32493 31464 32505 31467
rect 32088 31436 32505 31464
rect 32088 31424 32094 31436
rect 32493 31433 32505 31436
rect 32539 31433 32551 31467
rect 32493 31427 32551 31433
rect 32677 31467 32735 31473
rect 32677 31433 32689 31467
rect 32723 31464 32735 31467
rect 32950 31464 32956 31476
rect 32723 31436 32956 31464
rect 32723 31433 32735 31436
rect 32677 31427 32735 31433
rect 32950 31424 32956 31436
rect 33008 31424 33014 31476
rect 35069 31467 35127 31473
rect 35069 31433 35081 31467
rect 35115 31464 35127 31467
rect 35250 31464 35256 31476
rect 35115 31436 35256 31464
rect 35115 31433 35127 31436
rect 35069 31427 35127 31433
rect 35250 31424 35256 31436
rect 35308 31424 35314 31476
rect 35342 31424 35348 31476
rect 35400 31464 35406 31476
rect 35618 31464 35624 31476
rect 35400 31436 35624 31464
rect 35400 31424 35406 31436
rect 35618 31424 35624 31436
rect 35676 31424 35682 31476
rect 37458 31464 37464 31476
rect 37419 31436 37464 31464
rect 37458 31424 37464 31436
rect 37516 31424 37522 31476
rect 37826 31424 37832 31476
rect 37884 31464 37890 31476
rect 37921 31467 37979 31473
rect 37921 31464 37933 31467
rect 37884 31436 37933 31464
rect 37884 31424 37890 31436
rect 37921 31433 37933 31436
rect 37967 31433 37979 31467
rect 37921 31427 37979 31433
rect 31220 31368 31754 31396
rect 31021 31359 31079 31365
rect 27246 31328 27252 31340
rect 26075 31297 26090 31328
rect 26252 31300 27252 31328
rect 26029 31291 26090 31297
rect 25280 31232 25820 31260
rect 25280 31220 25286 31232
rect 24360 31164 24440 31192
rect 25792 31192 25820 31232
rect 25958 31192 25964 31204
rect 25792 31164 25964 31192
rect 24360 31152 24366 31164
rect 25958 31152 25964 31164
rect 26016 31152 26022 31204
rect 26062 31136 26090 31291
rect 27246 31288 27252 31300
rect 27304 31288 27310 31340
rect 27430 31328 27436 31340
rect 27391 31300 27436 31328
rect 27430 31288 27436 31300
rect 27488 31288 27494 31340
rect 28537 31331 28595 31337
rect 28537 31328 28549 31331
rect 27540 31300 28549 31328
rect 26878 31220 26884 31272
rect 26936 31260 26942 31272
rect 27540 31260 27568 31300
rect 28537 31297 28549 31300
rect 28583 31297 28595 31331
rect 28537 31291 28595 31297
rect 28626 31288 28632 31340
rect 28684 31328 28690 31340
rect 28721 31331 28779 31337
rect 28721 31328 28733 31331
rect 28684 31300 28733 31328
rect 28684 31288 28690 31300
rect 28721 31297 28733 31300
rect 28767 31328 28779 31331
rect 28966 31328 28994 31356
rect 28767 31300 28994 31328
rect 28767 31297 28779 31300
rect 28721 31291 28779 31297
rect 29178 31288 29184 31340
rect 29236 31328 29242 31340
rect 29365 31331 29423 31337
rect 29365 31328 29377 31331
rect 29236 31300 29377 31328
rect 29236 31288 29242 31300
rect 29365 31297 29377 31300
rect 29411 31297 29423 31331
rect 29365 31291 29423 31297
rect 29549 31331 29607 31337
rect 29549 31297 29561 31331
rect 29595 31297 29607 31331
rect 30650 31328 30656 31340
rect 30611 31300 30656 31328
rect 29549 31291 29607 31297
rect 26936 31232 27568 31260
rect 26936 31220 26942 31232
rect 27614 31220 27620 31272
rect 27672 31260 27678 31272
rect 27709 31263 27767 31269
rect 27709 31260 27721 31263
rect 27672 31232 27721 31260
rect 27672 31220 27678 31232
rect 27709 31229 27721 31232
rect 27755 31229 27767 31263
rect 27709 31223 27767 31229
rect 27890 31220 27896 31272
rect 27948 31260 27954 31272
rect 28902 31260 28908 31272
rect 27948 31232 28908 31260
rect 27948 31220 27954 31232
rect 28902 31220 28908 31232
rect 28960 31220 28966 31272
rect 26418 31152 26424 31204
rect 26476 31192 26482 31204
rect 29564 31192 29592 31291
rect 30650 31288 30656 31300
rect 30708 31288 30714 31340
rect 30742 31288 30748 31340
rect 30800 31328 30806 31340
rect 30926 31328 30932 31340
rect 30800 31300 30845 31328
rect 30887 31300 30932 31328
rect 30800 31288 30806 31300
rect 30926 31288 30932 31300
rect 30984 31288 30990 31340
rect 31036 31260 31064 31359
rect 31159 31331 31217 31337
rect 31159 31297 31171 31331
rect 31205 31328 31217 31331
rect 31570 31328 31576 31340
rect 31205 31300 31576 31328
rect 31205 31297 31217 31300
rect 31159 31291 31217 31297
rect 31570 31288 31576 31300
rect 31628 31288 31634 31340
rect 31726 31328 31754 31368
rect 32122 31356 32128 31408
rect 32180 31396 32186 31408
rect 32309 31399 32367 31405
rect 32309 31396 32321 31399
rect 32180 31368 32321 31396
rect 32180 31356 32186 31368
rect 32309 31365 32321 31368
rect 32355 31365 32367 31399
rect 32309 31359 32367 31365
rect 34606 31356 34612 31408
rect 34664 31396 34670 31408
rect 34701 31399 34759 31405
rect 34701 31396 34713 31399
rect 34664 31368 34713 31396
rect 34664 31356 34670 31368
rect 34701 31365 34713 31368
rect 34747 31365 34759 31399
rect 34701 31359 34759 31365
rect 34793 31399 34851 31405
rect 34793 31365 34805 31399
rect 34839 31396 34851 31399
rect 35526 31396 35532 31408
rect 34839 31368 35532 31396
rect 34839 31365 34851 31368
rect 34793 31359 34851 31365
rect 35526 31356 35532 31368
rect 35584 31356 35590 31408
rect 34146 31328 34152 31340
rect 31726 31300 34152 31328
rect 34146 31288 34152 31300
rect 34204 31288 34210 31340
rect 34514 31328 34520 31340
rect 34475 31300 34520 31328
rect 34514 31288 34520 31300
rect 34572 31288 34578 31340
rect 34882 31328 34888 31340
rect 34843 31300 34888 31328
rect 34882 31288 34888 31300
rect 34940 31328 34946 31340
rect 35434 31328 35440 31340
rect 34940 31300 35440 31328
rect 34940 31288 34946 31300
rect 35434 31288 35440 31300
rect 35492 31288 35498 31340
rect 37734 31288 37740 31340
rect 37792 31328 37798 31340
rect 37829 31331 37887 31337
rect 37829 31328 37841 31331
rect 37792 31300 37841 31328
rect 37792 31288 37798 31300
rect 37829 31297 37841 31300
rect 37875 31297 37887 31331
rect 37829 31291 37887 31297
rect 34606 31260 34612 31272
rect 31036 31232 34612 31260
rect 34606 31220 34612 31232
rect 34664 31220 34670 31272
rect 38010 31260 38016 31272
rect 37971 31232 38016 31260
rect 38010 31220 38016 31232
rect 38068 31220 38074 31272
rect 26476 31164 29592 31192
rect 29641 31195 29699 31201
rect 26476 31152 26482 31164
rect 29641 31161 29653 31195
rect 29687 31192 29699 31195
rect 35986 31192 35992 31204
rect 29687 31164 31754 31192
rect 29687 31161 29699 31164
rect 29641 31155 29699 31161
rect 14277 31127 14335 31133
rect 14277 31093 14289 31127
rect 14323 31093 14335 31127
rect 14277 31087 14335 31093
rect 17313 31127 17371 31133
rect 17313 31093 17325 31127
rect 17359 31093 17371 31127
rect 17313 31087 17371 31093
rect 17494 31084 17500 31136
rect 17552 31124 17558 31136
rect 18325 31127 18383 31133
rect 18325 31124 18337 31127
rect 17552 31096 18337 31124
rect 17552 31084 17558 31096
rect 18325 31093 18337 31096
rect 18371 31093 18383 31127
rect 18325 31087 18383 31093
rect 18782 31084 18788 31136
rect 18840 31124 18846 31136
rect 20898 31124 20904 31136
rect 18840 31096 20904 31124
rect 18840 31084 18846 31096
rect 20898 31084 20904 31096
rect 20956 31084 20962 31136
rect 21269 31127 21327 31133
rect 21269 31093 21281 31127
rect 21315 31124 21327 31127
rect 22554 31124 22560 31136
rect 21315 31096 22560 31124
rect 21315 31093 21327 31096
rect 21269 31087 21327 31093
rect 22554 31084 22560 31096
rect 22612 31084 22618 31136
rect 25406 31124 25412 31136
rect 25367 31096 25412 31124
rect 25406 31084 25412 31096
rect 25464 31084 25470 31136
rect 26050 31084 26056 31136
rect 26108 31084 26114 31136
rect 31726 31124 31754 31164
rect 32324 31164 35992 31192
rect 32324 31124 32352 31164
rect 35986 31152 35992 31164
rect 36044 31152 36050 31204
rect 32490 31124 32496 31136
rect 31726 31096 32352 31124
rect 32451 31096 32496 31124
rect 32490 31084 32496 31096
rect 32548 31084 32554 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 6546 30920 6552 30932
rect 6507 30892 6552 30920
rect 6546 30880 6552 30892
rect 6604 30880 6610 30932
rect 7006 30920 7012 30932
rect 6967 30892 7012 30920
rect 7006 30880 7012 30892
rect 7064 30880 7070 30932
rect 7926 30920 7932 30932
rect 7887 30892 7932 30920
rect 7926 30880 7932 30892
rect 7984 30880 7990 30932
rect 9398 30880 9404 30932
rect 9456 30920 9462 30932
rect 10226 30920 10232 30932
rect 9456 30892 10232 30920
rect 9456 30880 9462 30892
rect 10226 30880 10232 30892
rect 10284 30880 10290 30932
rect 11425 30923 11483 30929
rect 11425 30889 11437 30923
rect 11471 30920 11483 30923
rect 12066 30920 12072 30932
rect 11471 30892 12072 30920
rect 11471 30889 11483 30892
rect 11425 30883 11483 30889
rect 12066 30880 12072 30892
rect 12124 30880 12130 30932
rect 12713 30923 12771 30929
rect 12713 30889 12725 30923
rect 12759 30920 12771 30923
rect 12986 30920 12992 30932
rect 12759 30892 12992 30920
rect 12759 30889 12771 30892
rect 12713 30883 12771 30889
rect 12986 30880 12992 30892
rect 13044 30880 13050 30932
rect 13541 30923 13599 30929
rect 13541 30889 13553 30923
rect 13587 30920 13599 30923
rect 14182 30920 14188 30932
rect 13587 30892 14188 30920
rect 13587 30889 13599 30892
rect 13541 30883 13599 30889
rect 14182 30880 14188 30892
rect 14240 30880 14246 30932
rect 15010 30880 15016 30932
rect 15068 30920 15074 30932
rect 17865 30923 17923 30929
rect 15068 30892 16528 30920
rect 15068 30880 15074 30892
rect 6914 30852 6920 30864
rect 5920 30824 6920 30852
rect 5920 30784 5948 30824
rect 6914 30812 6920 30824
rect 6972 30852 6978 30864
rect 7374 30852 7380 30864
rect 6972 30824 7380 30852
rect 6972 30812 6978 30824
rect 7374 30812 7380 30824
rect 7432 30812 7438 30864
rect 10594 30852 10600 30864
rect 9784 30824 10600 30852
rect 6638 30784 6644 30796
rect 5828 30756 5948 30784
rect 6599 30756 6644 30784
rect 5828 30725 5856 30756
rect 6638 30744 6644 30756
rect 6696 30744 6702 30796
rect 7190 30784 7196 30796
rect 6840 30756 7196 30784
rect 6840 30725 6868 30756
rect 7190 30744 7196 30756
rect 7248 30784 7254 30796
rect 8202 30784 8208 30796
rect 7248 30756 8208 30784
rect 7248 30744 7254 30756
rect 8202 30744 8208 30756
rect 8260 30784 8266 30796
rect 8389 30787 8447 30793
rect 8389 30784 8401 30787
rect 8260 30756 8401 30784
rect 8260 30744 8266 30756
rect 8389 30753 8401 30756
rect 8435 30753 8447 30787
rect 8389 30747 8447 30753
rect 5077 30719 5135 30725
rect 5077 30685 5089 30719
rect 5123 30716 5135 30719
rect 5813 30719 5871 30725
rect 5123 30688 5764 30716
rect 5123 30685 5135 30688
rect 5077 30679 5135 30685
rect 4890 30648 4896 30660
rect 4851 30620 4896 30648
rect 4890 30608 4896 30620
rect 4948 30608 4954 30660
rect 5258 30648 5264 30660
rect 5219 30620 5264 30648
rect 5258 30608 5264 30620
rect 5316 30608 5322 30660
rect 5736 30648 5764 30688
rect 5813 30685 5825 30719
rect 5859 30685 5871 30719
rect 5997 30719 6055 30725
rect 5997 30716 6009 30719
rect 5813 30679 5871 30685
rect 5920 30688 6009 30716
rect 5920 30648 5948 30688
rect 5997 30685 6009 30688
rect 6043 30716 6055 30719
rect 6825 30719 6883 30725
rect 6043 30688 6684 30716
rect 6043 30685 6055 30688
rect 5997 30679 6055 30685
rect 6086 30648 6092 30660
rect 5736 30620 5948 30648
rect 6047 30620 6092 30648
rect 6086 30608 6092 30620
rect 6144 30608 6150 30660
rect 6549 30651 6607 30657
rect 6549 30617 6561 30651
rect 6595 30617 6607 30651
rect 6656 30648 6684 30688
rect 6825 30685 6837 30719
rect 6871 30685 6883 30719
rect 8110 30716 8116 30728
rect 8071 30688 8116 30716
rect 6825 30679 6883 30685
rect 8110 30676 8116 30688
rect 8168 30676 8174 30728
rect 8297 30719 8355 30725
rect 8297 30685 8309 30719
rect 8343 30685 8355 30719
rect 8297 30679 8355 30685
rect 7558 30648 7564 30660
rect 6656 30620 7564 30648
rect 6549 30611 6607 30617
rect 6564 30580 6592 30611
rect 7558 30608 7564 30620
rect 7616 30608 7622 30660
rect 7926 30608 7932 30660
rect 7984 30648 7990 30660
rect 8312 30648 8340 30679
rect 9214 30676 9220 30728
rect 9272 30716 9278 30728
rect 9784 30725 9812 30824
rect 10594 30812 10600 30824
rect 10652 30812 10658 30864
rect 12434 30812 12440 30864
rect 12492 30852 12498 30864
rect 15470 30852 15476 30864
rect 12492 30824 12940 30852
rect 12492 30812 12498 30824
rect 10321 30787 10379 30793
rect 10321 30753 10333 30787
rect 10367 30784 10379 30787
rect 11054 30784 11060 30796
rect 10367 30756 11060 30784
rect 10367 30753 10379 30756
rect 10321 30747 10379 30753
rect 11054 30744 11060 30756
rect 11112 30744 11118 30796
rect 11716 30756 12756 30784
rect 11716 30728 11744 30756
rect 9769 30719 9827 30725
rect 9769 30716 9781 30719
rect 9272 30688 9781 30716
rect 9272 30676 9278 30688
rect 9769 30685 9781 30688
rect 9815 30685 9827 30719
rect 9953 30719 10011 30725
rect 9953 30716 9965 30719
rect 9769 30679 9827 30685
rect 9876 30688 9965 30716
rect 7984 30620 8340 30648
rect 7984 30608 7990 30620
rect 9876 30592 9904 30688
rect 9953 30685 9965 30688
rect 9999 30685 10011 30719
rect 11698 30716 11704 30728
rect 11659 30688 11704 30716
rect 9953 30679 10011 30685
rect 11698 30676 11704 30688
rect 11756 30676 11762 30728
rect 11974 30676 11980 30728
rect 12032 30716 12038 30728
rect 12069 30719 12127 30725
rect 12069 30716 12081 30719
rect 12032 30688 12081 30716
rect 12032 30676 12038 30688
rect 12069 30685 12081 30688
rect 12115 30685 12127 30719
rect 12069 30679 12127 30685
rect 12161 30719 12219 30725
rect 12161 30685 12173 30719
rect 12207 30716 12219 30719
rect 12342 30716 12348 30728
rect 12207 30688 12348 30716
rect 12207 30685 12219 30688
rect 12161 30679 12219 30685
rect 12342 30676 12348 30688
rect 12400 30676 12406 30728
rect 12728 30725 12756 30756
rect 12912 30725 12940 30824
rect 13372 30824 15476 30852
rect 13372 30728 13400 30824
rect 13633 30787 13691 30793
rect 13633 30753 13645 30787
rect 13679 30784 13691 30787
rect 13722 30784 13728 30796
rect 13679 30756 13728 30784
rect 13679 30753 13691 30756
rect 13633 30747 13691 30753
rect 13722 30744 13728 30756
rect 13780 30744 13786 30796
rect 12713 30719 12771 30725
rect 12713 30685 12725 30719
rect 12759 30685 12771 30719
rect 12713 30679 12771 30685
rect 12897 30719 12955 30725
rect 12897 30685 12909 30719
rect 12943 30716 12955 30719
rect 13354 30716 13360 30728
rect 12943 30688 13360 30716
rect 12943 30685 12955 30688
rect 12897 30679 12955 30685
rect 13354 30676 13360 30688
rect 13412 30676 13418 30728
rect 13449 30719 13507 30725
rect 13449 30685 13461 30719
rect 13495 30685 13507 30719
rect 13449 30679 13507 30685
rect 11885 30651 11943 30657
rect 11885 30617 11897 30651
rect 11931 30648 11943 30651
rect 12802 30648 12808 30660
rect 11931 30620 12808 30648
rect 11931 30617 11943 30620
rect 11885 30611 11943 30617
rect 12802 30608 12808 30620
rect 12860 30648 12866 30660
rect 13464 30648 13492 30679
rect 15010 30676 15016 30728
rect 15068 30716 15074 30728
rect 15304 30725 15332 30824
rect 15470 30812 15476 30824
rect 15528 30812 15534 30864
rect 16500 30852 16528 30892
rect 17865 30889 17877 30923
rect 17911 30920 17923 30923
rect 19334 30920 19340 30932
rect 17911 30892 19340 30920
rect 17911 30889 17923 30892
rect 17865 30883 17923 30889
rect 19334 30880 19340 30892
rect 19392 30880 19398 30932
rect 19702 30920 19708 30932
rect 19663 30892 19708 30920
rect 19702 30880 19708 30892
rect 19760 30880 19766 30932
rect 20438 30920 20444 30932
rect 20399 30892 20444 30920
rect 20438 30880 20444 30892
rect 20496 30880 20502 30932
rect 20898 30880 20904 30932
rect 20956 30920 20962 30932
rect 22002 30920 22008 30932
rect 20956 30892 22008 30920
rect 20956 30880 20962 30892
rect 22002 30880 22008 30892
rect 22060 30880 22066 30932
rect 22278 30880 22284 30932
rect 22336 30920 22342 30932
rect 25038 30920 25044 30932
rect 22336 30892 25044 30920
rect 22336 30880 22342 30892
rect 25038 30880 25044 30892
rect 25096 30880 25102 30932
rect 28261 30923 28319 30929
rect 28261 30889 28273 30923
rect 28307 30920 28319 30923
rect 29638 30920 29644 30932
rect 28307 30892 29644 30920
rect 28307 30889 28319 30892
rect 28261 30883 28319 30889
rect 29638 30880 29644 30892
rect 29696 30880 29702 30932
rect 31110 30880 31116 30932
rect 31168 30920 31174 30932
rect 34238 30920 34244 30932
rect 31168 30892 34244 30920
rect 31168 30880 31174 30892
rect 34238 30880 34244 30892
rect 34296 30880 34302 30932
rect 25406 30852 25412 30864
rect 16500 30824 19840 30852
rect 17773 30787 17831 30793
rect 17773 30753 17785 30787
rect 17819 30784 17831 30787
rect 17819 30756 18000 30784
rect 17819 30753 17831 30756
rect 17773 30747 17831 30753
rect 15105 30719 15163 30725
rect 15105 30716 15117 30719
rect 15068 30688 15117 30716
rect 15068 30676 15074 30688
rect 15105 30685 15117 30688
rect 15151 30685 15163 30719
rect 15105 30679 15163 30685
rect 15289 30719 15347 30725
rect 15289 30685 15301 30719
rect 15335 30685 15347 30719
rect 15289 30679 15347 30685
rect 15381 30719 15439 30725
rect 15381 30685 15393 30719
rect 15427 30685 15439 30719
rect 15381 30679 15439 30685
rect 12860 30620 13492 30648
rect 12860 30608 12866 30620
rect 13538 30608 13544 30660
rect 13596 30648 13602 30660
rect 15396 30648 15424 30679
rect 15470 30676 15476 30728
rect 15528 30716 15534 30728
rect 15657 30719 15715 30725
rect 15528 30688 15573 30716
rect 15528 30676 15534 30688
rect 15657 30685 15669 30719
rect 15703 30716 15715 30719
rect 15838 30716 15844 30728
rect 15703 30688 15844 30716
rect 15703 30685 15715 30688
rect 15657 30679 15715 30685
rect 15838 30676 15844 30688
rect 15896 30716 15902 30728
rect 16393 30719 16451 30725
rect 16393 30716 16405 30719
rect 15896 30688 16405 30716
rect 15896 30676 15902 30688
rect 16393 30685 16405 30688
rect 16439 30685 16451 30719
rect 16574 30716 16580 30728
rect 16535 30688 16580 30716
rect 16393 30679 16451 30685
rect 16574 30676 16580 30688
rect 16632 30676 16638 30728
rect 17218 30676 17224 30728
rect 17276 30716 17282 30728
rect 17865 30719 17923 30725
rect 17865 30716 17877 30719
rect 17276 30688 17877 30716
rect 17276 30676 17282 30688
rect 17865 30685 17877 30688
rect 17911 30685 17923 30719
rect 17865 30679 17923 30685
rect 13596 30620 15424 30648
rect 16761 30651 16819 30657
rect 13596 30608 13602 30620
rect 16761 30617 16773 30651
rect 16807 30648 16819 30651
rect 17494 30648 17500 30660
rect 16807 30620 17500 30648
rect 16807 30617 16819 30620
rect 16761 30611 16819 30617
rect 17494 30608 17500 30620
rect 17552 30608 17558 30660
rect 17586 30608 17592 30660
rect 17644 30648 17650 30660
rect 17972 30648 18000 30756
rect 18690 30744 18696 30796
rect 18748 30784 18754 30796
rect 19521 30787 19579 30793
rect 19521 30784 19533 30787
rect 18748 30756 19533 30784
rect 18748 30744 18754 30756
rect 19521 30753 19533 30756
rect 19567 30753 19579 30787
rect 19812 30784 19840 30824
rect 20088 30824 25412 30852
rect 20088 30784 20116 30824
rect 25406 30812 25412 30824
rect 25464 30812 25470 30864
rect 25866 30812 25872 30864
rect 25924 30852 25930 30864
rect 26237 30855 26295 30861
rect 26237 30852 26249 30855
rect 25924 30824 26249 30852
rect 25924 30812 25930 30824
rect 26237 30821 26249 30824
rect 26283 30821 26295 30855
rect 26237 30815 26295 30821
rect 19812 30756 20116 30784
rect 19521 30747 19579 30753
rect 20438 30744 20444 30796
rect 20496 30784 20502 30796
rect 20625 30787 20683 30793
rect 20625 30784 20637 30787
rect 20496 30756 20637 30784
rect 20496 30744 20502 30756
rect 20625 30753 20637 30756
rect 20671 30753 20683 30787
rect 20625 30747 20683 30753
rect 21450 30744 21456 30796
rect 21508 30784 21514 30796
rect 23014 30784 23020 30796
rect 21508 30756 23020 30784
rect 21508 30744 21514 30756
rect 19705 30719 19763 30725
rect 19705 30685 19717 30719
rect 19751 30716 19763 30719
rect 19978 30716 19984 30728
rect 19751 30688 19984 30716
rect 19751 30685 19763 30688
rect 19705 30679 19763 30685
rect 19978 30676 19984 30688
rect 20036 30676 20042 30728
rect 20349 30719 20407 30725
rect 20349 30685 20361 30719
rect 20395 30716 20407 30719
rect 20530 30716 20536 30728
rect 20395 30688 20536 30716
rect 20395 30685 20407 30688
rect 20349 30679 20407 30685
rect 20530 30676 20536 30688
rect 20588 30676 20594 30728
rect 22278 30716 22284 30728
rect 22239 30688 22284 30716
rect 22278 30676 22284 30688
rect 22336 30676 22342 30728
rect 22664 30725 22692 30756
rect 23014 30744 23020 30756
rect 23072 30744 23078 30796
rect 23198 30744 23204 30796
rect 23256 30784 23262 30796
rect 26252 30784 26280 30815
rect 27246 30812 27252 30864
rect 27304 30852 27310 30864
rect 28902 30852 28908 30864
rect 27304 30824 28304 30852
rect 28863 30824 28908 30852
rect 27304 30812 27310 30824
rect 27430 30784 27436 30796
rect 23256 30756 25452 30784
rect 26252 30756 26832 30784
rect 23256 30744 23262 30756
rect 22649 30719 22707 30725
rect 22649 30685 22661 30719
rect 22695 30685 22707 30719
rect 22649 30679 22707 30685
rect 22738 30676 22744 30728
rect 22796 30716 22802 30728
rect 23293 30719 23351 30725
rect 23293 30716 23305 30719
rect 22796 30688 23305 30716
rect 22796 30676 22802 30688
rect 23293 30685 23305 30688
rect 23339 30685 23351 30719
rect 23293 30679 23351 30685
rect 23385 30719 23443 30725
rect 23385 30685 23397 30719
rect 23431 30716 23443 30719
rect 23474 30716 23480 30728
rect 23431 30688 23480 30716
rect 23431 30685 23443 30688
rect 23385 30679 23443 30685
rect 23474 30676 23480 30688
rect 23532 30676 23538 30728
rect 23566 30676 23572 30728
rect 23624 30716 23630 30728
rect 23750 30716 23756 30728
rect 23624 30688 23756 30716
rect 23624 30676 23630 30688
rect 23750 30676 23756 30688
rect 23808 30676 23814 30728
rect 24854 30676 24860 30728
rect 24912 30716 24918 30728
rect 24949 30719 25007 30725
rect 24949 30716 24961 30719
rect 24912 30688 24961 30716
rect 24912 30676 24918 30688
rect 24949 30685 24961 30688
rect 24995 30685 25007 30719
rect 25130 30716 25136 30728
rect 25091 30688 25136 30716
rect 24949 30679 25007 30685
rect 25130 30676 25136 30688
rect 25188 30676 25194 30728
rect 25424 30725 25452 30756
rect 25317 30719 25375 30725
rect 25317 30716 25329 30719
rect 25240 30688 25329 30716
rect 17644 30620 17689 30648
rect 17880 30620 18000 30648
rect 19429 30651 19487 30657
rect 17644 30608 17650 30620
rect 17880 30592 17908 30620
rect 19429 30617 19441 30651
rect 19475 30648 19487 30651
rect 22833 30651 22891 30657
rect 19475 30620 20392 30648
rect 19475 30617 19487 30620
rect 19429 30611 19487 30617
rect 9858 30580 9864 30592
rect 6564 30552 9864 30580
rect 9858 30540 9864 30552
rect 9916 30540 9922 30592
rect 11146 30540 11152 30592
rect 11204 30580 11210 30592
rect 11793 30583 11851 30589
rect 11793 30580 11805 30583
rect 11204 30552 11805 30580
rect 11204 30540 11210 30552
rect 11793 30549 11805 30552
rect 11839 30549 11851 30583
rect 11793 30543 11851 30549
rect 12526 30540 12532 30592
rect 12584 30580 12590 30592
rect 15010 30580 15016 30592
rect 12584 30552 15016 30580
rect 12584 30540 12590 30552
rect 15010 30540 15016 30552
rect 15068 30540 15074 30592
rect 15194 30540 15200 30592
rect 15252 30580 15258 30592
rect 15841 30583 15899 30589
rect 15841 30580 15853 30583
rect 15252 30552 15853 30580
rect 15252 30540 15258 30552
rect 15841 30549 15853 30552
rect 15887 30549 15899 30583
rect 15841 30543 15899 30549
rect 17862 30540 17868 30592
rect 17920 30540 17926 30592
rect 18046 30580 18052 30592
rect 18007 30552 18052 30580
rect 18046 30540 18052 30552
rect 18104 30540 18110 30592
rect 18138 30540 18144 30592
rect 18196 30580 18202 30592
rect 19889 30583 19947 30589
rect 19889 30580 19901 30583
rect 18196 30552 19901 30580
rect 18196 30540 18202 30552
rect 19889 30549 19901 30552
rect 19935 30549 19947 30583
rect 20364 30580 20392 30620
rect 22833 30617 22845 30651
rect 22879 30648 22891 30651
rect 22922 30648 22928 30660
rect 22879 30620 22928 30648
rect 22879 30617 22891 30620
rect 22833 30611 22891 30617
rect 22922 30608 22928 30620
rect 22980 30608 22986 30660
rect 20625 30583 20683 30589
rect 20625 30580 20637 30583
rect 20364 30552 20637 30580
rect 19889 30543 19947 30549
rect 20625 30549 20637 30552
rect 20671 30580 20683 30583
rect 20898 30580 20904 30592
rect 20671 30552 20904 30580
rect 20671 30549 20683 30552
rect 20625 30543 20683 30549
rect 20898 30540 20904 30552
rect 20956 30540 20962 30592
rect 23750 30580 23756 30592
rect 23711 30552 23756 30580
rect 23750 30540 23756 30552
rect 23808 30540 23814 30592
rect 25240 30580 25268 30688
rect 25317 30685 25329 30688
rect 25363 30685 25375 30719
rect 25317 30679 25375 30685
rect 25409 30719 25467 30725
rect 25409 30685 25421 30719
rect 25455 30685 25467 30719
rect 25409 30679 25467 30685
rect 25498 30676 25504 30728
rect 25556 30716 25562 30728
rect 25869 30719 25927 30725
rect 25869 30716 25881 30719
rect 25556 30688 25881 30716
rect 25556 30676 25562 30688
rect 25869 30685 25881 30688
rect 25915 30685 25927 30719
rect 25869 30679 25927 30685
rect 25958 30676 25964 30728
rect 26016 30716 26022 30728
rect 26697 30719 26755 30725
rect 26697 30716 26709 30719
rect 26016 30688 26709 30716
rect 26016 30676 26022 30688
rect 26697 30685 26709 30688
rect 26743 30685 26755 30719
rect 26697 30679 26755 30685
rect 25682 30608 25688 30660
rect 25740 30648 25746 30660
rect 26053 30651 26111 30657
rect 26053 30648 26065 30651
rect 25740 30620 26065 30648
rect 25740 30608 25746 30620
rect 26053 30617 26065 30620
rect 26099 30617 26111 30651
rect 26804 30648 26832 30756
rect 26896 30756 27436 30784
rect 26896 30725 26924 30756
rect 27430 30744 27436 30756
rect 27488 30744 27494 30796
rect 27890 30744 27896 30796
rect 27948 30784 27954 30796
rect 28169 30787 28227 30793
rect 28169 30784 28181 30787
rect 27948 30756 28181 30784
rect 27948 30744 27954 30756
rect 28169 30753 28181 30756
rect 28215 30753 28227 30787
rect 28276 30784 28304 30824
rect 28902 30812 28908 30824
rect 28960 30812 28966 30864
rect 31389 30855 31447 30861
rect 31389 30821 31401 30855
rect 31435 30852 31447 30855
rect 32490 30852 32496 30864
rect 31435 30824 32496 30852
rect 31435 30821 31447 30824
rect 31389 30815 31447 30821
rect 32416 30793 32444 30824
rect 32490 30812 32496 30824
rect 32548 30812 32554 30864
rect 32401 30787 32459 30793
rect 28276 30756 28948 30784
rect 28169 30747 28227 30753
rect 26881 30719 26939 30725
rect 26881 30685 26893 30719
rect 26927 30685 26939 30719
rect 26881 30679 26939 30685
rect 27341 30719 27399 30725
rect 27341 30685 27353 30719
rect 27387 30685 27399 30719
rect 27341 30679 27399 30685
rect 27525 30719 27583 30725
rect 27525 30685 27537 30719
rect 27571 30685 27583 30719
rect 27525 30679 27583 30685
rect 27356 30648 27384 30679
rect 26804 30620 27384 30648
rect 26053 30611 26111 30617
rect 26510 30580 26516 30592
rect 25240 30552 26516 30580
rect 26510 30540 26516 30552
rect 26568 30580 26574 30592
rect 26789 30583 26847 30589
rect 26789 30580 26801 30583
rect 26568 30552 26801 30580
rect 26568 30540 26574 30552
rect 26789 30549 26801 30552
rect 26835 30549 26847 30583
rect 27430 30580 27436 30592
rect 27391 30552 27436 30580
rect 26789 30543 26847 30549
rect 27430 30540 27436 30552
rect 27488 30540 27494 30592
rect 27540 30580 27568 30679
rect 27706 30676 27712 30728
rect 27764 30716 27770 30728
rect 28920 30725 28948 30756
rect 29748 30756 31064 30784
rect 28077 30719 28135 30725
rect 28077 30716 28089 30719
rect 27764 30688 28089 30716
rect 27764 30676 27770 30688
rect 28077 30685 28089 30688
rect 28123 30685 28135 30719
rect 28077 30679 28135 30685
rect 28905 30719 28963 30725
rect 28905 30685 28917 30719
rect 28951 30685 28963 30719
rect 28905 30679 28963 30685
rect 28994 30676 29000 30728
rect 29052 30716 29058 30728
rect 29748 30725 29776 30756
rect 29089 30719 29147 30725
rect 29089 30716 29101 30719
rect 29052 30688 29101 30716
rect 29052 30676 29058 30688
rect 29089 30685 29101 30688
rect 29135 30685 29147 30719
rect 29089 30679 29147 30685
rect 29733 30719 29791 30725
rect 29733 30685 29745 30719
rect 29779 30685 29791 30719
rect 30742 30716 30748 30728
rect 30703 30688 30748 30716
rect 29733 30679 29791 30685
rect 30742 30676 30748 30688
rect 30800 30676 30806 30728
rect 30834 30676 30840 30728
rect 30892 30716 30898 30728
rect 31036 30716 31064 30756
rect 32401 30753 32413 30787
rect 32447 30753 32459 30787
rect 32401 30747 32459 30753
rect 32677 30787 32735 30793
rect 32677 30753 32689 30787
rect 32723 30784 32735 30787
rect 34054 30784 34060 30796
rect 32723 30756 34060 30784
rect 32723 30753 32735 30756
rect 32677 30747 32735 30753
rect 34054 30744 34060 30756
rect 34112 30744 34118 30796
rect 34606 30744 34612 30796
rect 34664 30784 34670 30796
rect 35526 30784 35532 30796
rect 34664 30756 35532 30784
rect 34664 30744 34670 30756
rect 31251 30719 31309 30725
rect 31251 30716 31263 30719
rect 30892 30688 30937 30716
rect 31036 30688 31263 30716
rect 30892 30676 30898 30688
rect 31251 30685 31263 30688
rect 31297 30716 31309 30719
rect 31570 30716 31576 30728
rect 31297 30688 31576 30716
rect 31297 30685 31309 30688
rect 31251 30679 31309 30685
rect 31570 30676 31576 30688
rect 31628 30676 31634 30728
rect 32122 30676 32128 30728
rect 32180 30716 32186 30728
rect 32309 30719 32367 30725
rect 32309 30716 32321 30719
rect 32180 30688 32321 30716
rect 32180 30676 32186 30688
rect 32309 30685 32321 30688
rect 32355 30716 32367 30719
rect 32582 30716 32588 30728
rect 32355 30688 32588 30716
rect 32355 30685 32367 30688
rect 32309 30679 32367 30685
rect 32582 30676 32588 30688
rect 32640 30676 32646 30728
rect 35360 30725 35388 30756
rect 35526 30744 35532 30756
rect 35584 30744 35590 30796
rect 35069 30719 35127 30725
rect 35069 30716 35081 30719
rect 33152 30688 35081 30716
rect 27982 30608 27988 30660
rect 28040 30648 28046 30660
rect 29917 30651 29975 30657
rect 29917 30648 29929 30651
rect 28040 30620 29929 30648
rect 28040 30608 28046 30620
rect 29917 30617 29929 30620
rect 29963 30617 29975 30651
rect 29917 30611 29975 30617
rect 30101 30651 30159 30657
rect 30101 30617 30113 30651
rect 30147 30648 30159 30651
rect 30190 30648 30196 30660
rect 30147 30620 30196 30648
rect 30147 30617 30159 30620
rect 30101 30611 30159 30617
rect 30190 30608 30196 30620
rect 30248 30608 30254 30660
rect 30926 30608 30932 30660
rect 30984 30648 30990 30660
rect 31021 30651 31079 30657
rect 31021 30648 31033 30651
rect 30984 30620 31033 30648
rect 30984 30608 30990 30620
rect 31021 30617 31033 30620
rect 31067 30617 31079 30651
rect 31021 30611 31079 30617
rect 28166 30580 28172 30592
rect 27540 30552 28172 30580
rect 28166 30540 28172 30552
rect 28224 30540 28230 30592
rect 28445 30583 28503 30589
rect 28445 30549 28457 30583
rect 28491 30580 28503 30583
rect 28626 30580 28632 30592
rect 28491 30552 28632 30580
rect 28491 30549 28503 30552
rect 28445 30543 28503 30549
rect 28626 30540 28632 30552
rect 28684 30540 28690 30592
rect 31036 30580 31064 30611
rect 31110 30608 31116 30660
rect 31168 30648 31174 30660
rect 31168 30620 31754 30648
rect 31168 30608 31174 30620
rect 31386 30580 31392 30592
rect 31036 30552 31392 30580
rect 31386 30540 31392 30552
rect 31444 30540 31450 30592
rect 31726 30580 31754 30620
rect 31846 30608 31852 30660
rect 31904 30648 31910 30660
rect 33152 30648 33180 30688
rect 35069 30685 35081 30688
rect 35115 30685 35127 30719
rect 35069 30679 35127 30685
rect 35345 30719 35403 30725
rect 35345 30685 35357 30719
rect 35391 30685 35403 30719
rect 35345 30679 35403 30685
rect 35434 30676 35440 30728
rect 35492 30716 35498 30728
rect 36722 30716 36728 30728
rect 35492 30688 35537 30716
rect 36683 30688 36728 30716
rect 35492 30676 35498 30688
rect 36722 30676 36728 30688
rect 36780 30676 36786 30728
rect 31904 30620 33180 30648
rect 31904 30608 31910 30620
rect 34790 30608 34796 30660
rect 34848 30648 34854 30660
rect 35253 30651 35311 30657
rect 35253 30648 35265 30651
rect 34848 30620 35265 30648
rect 34848 30608 34854 30620
rect 35253 30617 35265 30620
rect 35299 30617 35311 30651
rect 36998 30648 37004 30660
rect 36959 30620 37004 30648
rect 35253 30611 35311 30617
rect 36998 30608 37004 30620
rect 37056 30608 37062 30660
rect 37274 30608 37280 30660
rect 37332 30648 37338 30660
rect 37737 30651 37795 30657
rect 37737 30648 37749 30651
rect 37332 30620 37749 30648
rect 37332 30608 37338 30620
rect 37737 30617 37749 30620
rect 37783 30617 37795 30651
rect 37737 30611 37795 30617
rect 35526 30580 35532 30592
rect 31726 30552 35532 30580
rect 35526 30540 35532 30552
rect 35584 30540 35590 30592
rect 35621 30583 35679 30589
rect 35621 30549 35633 30583
rect 35667 30580 35679 30583
rect 35802 30580 35808 30592
rect 35667 30552 35808 30580
rect 35667 30549 35679 30552
rect 35621 30543 35679 30549
rect 35802 30540 35808 30552
rect 35860 30540 35866 30592
rect 38010 30580 38016 30592
rect 37971 30552 38016 30580
rect 38010 30540 38016 30552
rect 38068 30540 38074 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 4890 30336 4896 30388
rect 4948 30376 4954 30388
rect 6546 30376 6552 30388
rect 4948 30348 6552 30376
rect 4948 30336 4954 30348
rect 6546 30336 6552 30348
rect 6604 30376 6610 30388
rect 7466 30376 7472 30388
rect 6604 30348 7472 30376
rect 6604 30336 6610 30348
rect 7466 30336 7472 30348
rect 7524 30376 7530 30388
rect 7926 30376 7932 30388
rect 7524 30348 7932 30376
rect 7524 30336 7530 30348
rect 7926 30336 7932 30348
rect 7984 30336 7990 30388
rect 9674 30336 9680 30388
rect 9732 30376 9738 30388
rect 10318 30376 10324 30388
rect 9732 30348 10324 30376
rect 9732 30336 9738 30348
rect 10318 30336 10324 30348
rect 10376 30336 10382 30388
rect 11790 30336 11796 30388
rect 11848 30376 11854 30388
rect 11848 30348 12480 30376
rect 11848 30336 11854 30348
rect 9582 30308 9588 30320
rect 2884 30280 9588 30308
rect 2774 30200 2780 30252
rect 2832 30240 2838 30252
rect 2884 30249 2912 30280
rect 9582 30268 9588 30280
rect 9640 30268 9646 30320
rect 10505 30311 10563 30317
rect 10505 30308 10517 30311
rect 9688 30280 10517 30308
rect 2869 30243 2927 30249
rect 2869 30240 2881 30243
rect 2832 30212 2881 30240
rect 2832 30200 2838 30212
rect 2869 30209 2881 30212
rect 2915 30209 2927 30243
rect 2869 30203 2927 30209
rect 3136 30243 3194 30249
rect 3136 30209 3148 30243
rect 3182 30240 3194 30243
rect 3970 30240 3976 30252
rect 3182 30212 3976 30240
rect 3182 30209 3194 30212
rect 3136 30203 3194 30209
rect 3970 30200 3976 30212
rect 4028 30200 4034 30252
rect 5169 30243 5227 30249
rect 5169 30209 5181 30243
rect 5215 30240 5227 30243
rect 5534 30240 5540 30252
rect 5215 30212 5540 30240
rect 5215 30209 5227 30212
rect 5169 30203 5227 30209
rect 5534 30200 5540 30212
rect 5592 30200 5598 30252
rect 6362 30200 6368 30252
rect 6420 30240 6426 30252
rect 6733 30243 6791 30249
rect 6733 30240 6745 30243
rect 6420 30212 6745 30240
rect 6420 30200 6426 30212
rect 6733 30209 6745 30212
rect 6779 30209 6791 30243
rect 6733 30203 6791 30209
rect 6914 30200 6920 30252
rect 6972 30240 6978 30252
rect 7009 30243 7067 30249
rect 7009 30240 7021 30243
rect 6972 30212 7021 30240
rect 6972 30200 6978 30212
rect 7009 30209 7021 30212
rect 7055 30209 7067 30243
rect 8662 30240 8668 30252
rect 8623 30212 8668 30240
rect 7009 30203 7067 30209
rect 8662 30200 8668 30212
rect 8720 30200 8726 30252
rect 9030 30240 9036 30252
rect 8991 30212 9036 30240
rect 9030 30200 9036 30212
rect 9088 30240 9094 30252
rect 9306 30240 9312 30252
rect 9088 30212 9312 30240
rect 9088 30200 9094 30212
rect 9306 30200 9312 30212
rect 9364 30200 9370 30252
rect 5353 30175 5411 30181
rect 5353 30141 5365 30175
rect 5399 30172 5411 30175
rect 6270 30172 6276 30184
rect 5399 30144 6276 30172
rect 5399 30141 5411 30144
rect 5353 30135 5411 30141
rect 6270 30132 6276 30144
rect 6328 30132 6334 30184
rect 6546 30172 6552 30184
rect 6507 30144 6552 30172
rect 6546 30132 6552 30144
rect 6604 30132 6610 30184
rect 6825 30175 6883 30181
rect 6825 30141 6837 30175
rect 6871 30172 6883 30175
rect 7098 30172 7104 30184
rect 6871 30144 7104 30172
rect 6871 30141 6883 30144
rect 6825 30135 6883 30141
rect 7098 30132 7104 30144
rect 7156 30132 7162 30184
rect 8110 30132 8116 30184
rect 8168 30172 8174 30184
rect 9688 30172 9716 30280
rect 10505 30277 10517 30280
rect 10551 30308 10563 30311
rect 11974 30308 11980 30320
rect 10551 30280 11980 30308
rect 10551 30277 10563 30280
rect 10505 30271 10563 30277
rect 11974 30268 11980 30280
rect 12032 30268 12038 30320
rect 12452 30317 12480 30348
rect 13832 30348 14412 30376
rect 13832 30317 13860 30348
rect 12437 30311 12495 30317
rect 12437 30277 12449 30311
rect 12483 30277 12495 30311
rect 12437 30271 12495 30277
rect 13817 30311 13875 30317
rect 13817 30277 13829 30311
rect 13863 30277 13875 30311
rect 14182 30308 14188 30320
rect 13817 30271 13875 30277
rect 14016 30280 14188 30308
rect 9953 30243 10011 30249
rect 9953 30209 9965 30243
rect 9999 30240 10011 30243
rect 10042 30240 10048 30252
rect 9999 30212 10048 30240
rect 9999 30209 10011 30212
rect 9953 30203 10011 30209
rect 10042 30200 10048 30212
rect 10100 30200 10106 30252
rect 10134 30200 10140 30252
rect 10192 30240 10198 30252
rect 12069 30243 12127 30249
rect 12069 30240 12081 30243
rect 10192 30212 12081 30240
rect 10192 30200 10198 30212
rect 12069 30209 12081 30212
rect 12115 30209 12127 30243
rect 12069 30203 12127 30209
rect 12253 30243 12311 30249
rect 12253 30209 12265 30243
rect 12299 30209 12311 30243
rect 12253 30203 12311 30209
rect 12897 30243 12955 30249
rect 12897 30209 12909 30243
rect 12943 30240 12955 30243
rect 13906 30240 13912 30252
rect 12943 30212 13912 30240
rect 12943 30209 12955 30212
rect 12897 30203 12955 30209
rect 8168 30144 9716 30172
rect 8168 30132 8174 30144
rect 11974 30132 11980 30184
rect 12032 30172 12038 30184
rect 12268 30172 12296 30203
rect 13906 30200 13912 30212
rect 13964 30200 13970 30252
rect 14016 30249 14044 30280
rect 14182 30268 14188 30280
rect 14240 30268 14246 30320
rect 14384 30308 14412 30348
rect 14458 30336 14464 30388
rect 14516 30376 14522 30388
rect 15105 30379 15163 30385
rect 15105 30376 15117 30379
rect 14516 30348 15117 30376
rect 14516 30336 14522 30348
rect 15105 30345 15117 30348
rect 15151 30376 15163 30379
rect 15746 30376 15752 30388
rect 15151 30348 15752 30376
rect 15151 30345 15163 30348
rect 15105 30339 15163 30345
rect 15746 30336 15752 30348
rect 15804 30336 15810 30388
rect 16574 30336 16580 30388
rect 16632 30376 16638 30388
rect 23198 30376 23204 30388
rect 16632 30348 23204 30376
rect 16632 30336 16638 30348
rect 23198 30336 23204 30348
rect 23256 30336 23262 30388
rect 23566 30336 23572 30388
rect 23624 30376 23630 30388
rect 26234 30376 26240 30388
rect 23624 30348 26240 30376
rect 23624 30336 23630 30348
rect 26234 30336 26240 30348
rect 26292 30336 26298 30388
rect 30377 30379 30435 30385
rect 30377 30345 30389 30379
rect 30423 30376 30435 30379
rect 30650 30376 30656 30388
rect 30423 30348 30656 30376
rect 30423 30345 30435 30348
rect 30377 30339 30435 30345
rect 30650 30336 30656 30348
rect 30708 30336 30714 30388
rect 30834 30336 30840 30388
rect 30892 30376 30898 30388
rect 35161 30379 35219 30385
rect 35161 30376 35173 30379
rect 30892 30348 35173 30376
rect 30892 30336 30898 30348
rect 35161 30345 35173 30348
rect 35207 30345 35219 30379
rect 35161 30339 35219 30345
rect 18138 30308 18144 30320
rect 14384 30280 18144 30308
rect 18138 30268 18144 30280
rect 18196 30268 18202 30320
rect 20254 30308 20260 30320
rect 20215 30280 20260 30308
rect 20254 30268 20260 30280
rect 20312 30308 20318 30320
rect 20312 30280 23428 30308
rect 20312 30268 20318 30280
rect 14001 30243 14059 30249
rect 14001 30209 14013 30243
rect 14047 30209 14059 30243
rect 14001 30203 14059 30209
rect 14093 30243 14151 30249
rect 14093 30209 14105 30243
rect 14139 30240 14151 30243
rect 14458 30240 14464 30252
rect 14139 30212 14464 30240
rect 14139 30209 14151 30212
rect 14093 30203 14151 30209
rect 14458 30200 14464 30212
rect 14516 30200 14522 30252
rect 14737 30243 14795 30249
rect 14737 30209 14749 30243
rect 14783 30209 14795 30243
rect 14737 30203 14795 30209
rect 13170 30172 13176 30184
rect 12032 30144 12296 30172
rect 13131 30144 13176 30172
rect 12032 30132 12038 30144
rect 13170 30132 13176 30144
rect 13228 30132 13234 30184
rect 13262 30132 13268 30184
rect 13320 30172 13326 30184
rect 14752 30172 14780 30203
rect 15194 30200 15200 30252
rect 15252 30240 15258 30252
rect 15657 30243 15715 30249
rect 15252 30212 15297 30240
rect 15252 30200 15258 30212
rect 15657 30209 15669 30243
rect 15703 30240 15715 30243
rect 16022 30240 16028 30252
rect 15703 30212 16028 30240
rect 15703 30209 15715 30212
rect 15657 30203 15715 30209
rect 16022 30200 16028 30212
rect 16080 30200 16086 30252
rect 17405 30243 17463 30249
rect 17405 30209 17417 30243
rect 17451 30240 17463 30243
rect 18046 30240 18052 30252
rect 17451 30212 18052 30240
rect 17451 30209 17463 30212
rect 17405 30203 17463 30209
rect 18046 30200 18052 30212
rect 18104 30200 18110 30252
rect 18233 30243 18291 30249
rect 18233 30209 18245 30243
rect 18279 30209 18291 30243
rect 18233 30203 18291 30209
rect 18417 30243 18475 30249
rect 18417 30209 18429 30243
rect 18463 30240 18475 30243
rect 18598 30240 18604 30252
rect 18463 30212 18604 30240
rect 18463 30209 18475 30212
rect 18417 30203 18475 30209
rect 15746 30172 15752 30184
rect 13320 30144 14780 30172
rect 15707 30144 15752 30172
rect 13320 30132 13326 30144
rect 5442 30064 5448 30116
rect 5500 30104 5506 30116
rect 6917 30107 6975 30113
rect 6917 30104 6929 30107
rect 5500 30076 6929 30104
rect 5500 30064 5506 30076
rect 6917 30073 6929 30076
rect 6963 30073 6975 30107
rect 12802 30104 12808 30116
rect 6917 30067 6975 30073
rect 7024 30076 12808 30104
rect 4249 30039 4307 30045
rect 4249 30005 4261 30039
rect 4295 30036 4307 30039
rect 4614 30036 4620 30048
rect 4295 30008 4620 30036
rect 4295 30005 4307 30008
rect 4249 29999 4307 30005
rect 4614 29996 4620 30008
rect 4672 30036 4678 30048
rect 7024 30036 7052 30076
rect 12802 30064 12808 30076
rect 12860 30064 12866 30116
rect 14277 30107 14335 30113
rect 13648 30076 14044 30104
rect 8202 30036 8208 30048
rect 4672 30008 7052 30036
rect 8163 30008 8208 30036
rect 4672 29996 4678 30008
rect 8202 29996 8208 30008
rect 8260 29996 8266 30048
rect 12820 30036 12848 30064
rect 13648 30036 13676 30076
rect 13814 30036 13820 30048
rect 12820 30008 13676 30036
rect 13775 30008 13820 30036
rect 13814 29996 13820 30008
rect 13872 29996 13878 30048
rect 14016 30036 14044 30076
rect 14277 30073 14289 30107
rect 14323 30104 14335 30107
rect 14642 30104 14648 30116
rect 14323 30076 14648 30104
rect 14323 30073 14335 30076
rect 14277 30067 14335 30073
rect 14642 30064 14648 30076
rect 14700 30064 14706 30116
rect 14752 30104 14780 30144
rect 15746 30132 15752 30144
rect 15804 30132 15810 30184
rect 17494 30172 17500 30184
rect 17455 30144 17500 30172
rect 17494 30132 17500 30144
rect 17552 30132 17558 30184
rect 17954 30172 17960 30184
rect 17604 30144 17960 30172
rect 16298 30104 16304 30116
rect 14752 30076 16304 30104
rect 16298 30064 16304 30076
rect 16356 30064 16362 30116
rect 16850 30064 16856 30116
rect 16908 30104 16914 30116
rect 17604 30104 17632 30144
rect 17954 30132 17960 30144
rect 18012 30132 18018 30184
rect 18248 30172 18276 30203
rect 18598 30200 18604 30212
rect 18656 30240 18662 30252
rect 19150 30240 19156 30252
rect 18656 30212 19156 30240
rect 18656 30200 18662 30212
rect 19150 30200 19156 30212
rect 19208 30200 19214 30252
rect 19978 30200 19984 30252
rect 20036 30240 20042 30252
rect 20438 30240 20444 30252
rect 20036 30212 20444 30240
rect 20036 30200 20042 30212
rect 20438 30200 20444 30212
rect 20496 30200 20502 30252
rect 22094 30200 22100 30252
rect 22152 30240 22158 30252
rect 22649 30243 22707 30249
rect 22152 30212 22232 30240
rect 22152 30200 22158 30212
rect 22204 30172 22232 30212
rect 22649 30209 22661 30243
rect 22695 30240 22707 30243
rect 22738 30240 22744 30252
rect 22695 30212 22744 30240
rect 22695 30209 22707 30212
rect 22649 30203 22707 30209
rect 22738 30200 22744 30212
rect 22796 30200 22802 30252
rect 22830 30200 22836 30252
rect 22888 30200 22894 30252
rect 22848 30172 22876 30200
rect 23014 30172 23020 30184
rect 18248 30144 19334 30172
rect 22204 30144 22876 30172
rect 22975 30144 23020 30172
rect 16908 30076 17632 30104
rect 16908 30064 16914 30076
rect 17678 30064 17684 30116
rect 17736 30104 17742 30116
rect 17773 30107 17831 30113
rect 17773 30104 17785 30107
rect 17736 30076 17785 30104
rect 17736 30064 17742 30076
rect 17773 30073 17785 30076
rect 17819 30073 17831 30107
rect 19306 30104 19334 30144
rect 23014 30132 23020 30144
rect 23072 30132 23078 30184
rect 23198 30172 23204 30184
rect 23159 30144 23204 30172
rect 23198 30132 23204 30144
rect 23256 30132 23262 30184
rect 23400 30172 23428 30280
rect 23658 30268 23664 30320
rect 23716 30308 23722 30320
rect 24305 30311 24363 30317
rect 24305 30308 24317 30311
rect 23716 30280 24317 30308
rect 23716 30268 23722 30280
rect 24305 30277 24317 30280
rect 24351 30277 24363 30311
rect 24305 30271 24363 30277
rect 24762 30268 24768 30320
rect 24820 30308 24826 30320
rect 24820 30280 27200 30308
rect 24820 30268 24826 30280
rect 24210 30200 24216 30252
rect 24268 30240 24274 30252
rect 24489 30243 24547 30249
rect 24489 30240 24501 30243
rect 24268 30212 24501 30240
rect 24268 30200 24274 30212
rect 24489 30209 24501 30212
rect 24535 30240 24547 30243
rect 24854 30240 24860 30252
rect 24535 30212 24860 30240
rect 24535 30209 24547 30212
rect 24489 30203 24547 30209
rect 24854 30200 24860 30212
rect 24912 30200 24918 30252
rect 25774 30200 25780 30252
rect 25832 30240 25838 30252
rect 26053 30243 26111 30249
rect 26053 30240 26065 30243
rect 25832 30212 26065 30240
rect 25832 30200 25838 30212
rect 26053 30209 26065 30212
rect 26099 30209 26111 30243
rect 26053 30203 26111 30209
rect 26234 30200 26240 30252
rect 26292 30240 26298 30252
rect 26421 30243 26479 30249
rect 26421 30240 26433 30243
rect 26292 30212 26433 30240
rect 26292 30200 26298 30212
rect 26421 30209 26433 30212
rect 26467 30209 26479 30243
rect 26421 30203 26479 30209
rect 26510 30200 26516 30252
rect 26568 30240 26574 30252
rect 27172 30249 27200 30280
rect 27540 30280 28120 30308
rect 27157 30243 27215 30249
rect 26568 30212 26613 30240
rect 26568 30200 26574 30212
rect 27157 30209 27169 30243
rect 27203 30209 27215 30243
rect 27157 30203 27215 30209
rect 24673 30175 24731 30181
rect 24673 30172 24685 30175
rect 23400 30144 24685 30172
rect 24673 30141 24685 30144
rect 24719 30172 24731 30175
rect 25222 30172 25228 30184
rect 24719 30144 25228 30172
rect 24719 30141 24731 30144
rect 24673 30135 24731 30141
rect 25222 30132 25228 30144
rect 25280 30132 25286 30184
rect 26145 30175 26203 30181
rect 26145 30141 26157 30175
rect 26191 30172 26203 30175
rect 27540 30172 27568 30280
rect 27617 30243 27675 30249
rect 27617 30209 27629 30243
rect 27663 30209 27675 30243
rect 27617 30203 27675 30209
rect 26191 30144 27568 30172
rect 26191 30141 26203 30144
rect 26145 30135 26203 30141
rect 19306 30076 22508 30104
rect 17773 30067 17831 30073
rect 14918 30045 14924 30048
rect 14875 30039 14924 30045
rect 14875 30036 14887 30039
rect 14016 30008 14887 30036
rect 14875 30005 14887 30008
rect 14921 30005 14924 30039
rect 14875 29999 14924 30005
rect 14918 29996 14924 29999
rect 14976 29996 14982 30048
rect 15013 30039 15071 30045
rect 15013 30005 15025 30039
rect 15059 30036 15071 30039
rect 15562 30036 15568 30048
rect 15059 30008 15568 30036
rect 15059 30005 15071 30008
rect 15013 29999 15071 30005
rect 15562 29996 15568 30008
rect 15620 29996 15626 30048
rect 15654 29996 15660 30048
rect 15712 30036 15718 30048
rect 15712 30008 15757 30036
rect 15712 29996 15718 30008
rect 15930 29996 15936 30048
rect 15988 30036 15994 30048
rect 16025 30039 16083 30045
rect 16025 30036 16037 30039
rect 15988 30008 16037 30036
rect 15988 29996 15994 30008
rect 16025 30005 16037 30008
rect 16071 30005 16083 30039
rect 17402 30036 17408 30048
rect 17363 30008 17408 30036
rect 16025 29999 16083 30005
rect 17402 29996 17408 30008
rect 17460 29996 17466 30048
rect 18230 30036 18236 30048
rect 18191 30008 18236 30036
rect 18230 29996 18236 30008
rect 18288 29996 18294 30048
rect 20622 30036 20628 30048
rect 20583 30008 20628 30036
rect 20622 29996 20628 30008
rect 20680 29996 20686 30048
rect 22480 30036 22508 30076
rect 22554 30064 22560 30116
rect 22612 30104 22618 30116
rect 22787 30107 22845 30113
rect 22787 30104 22799 30107
rect 22612 30076 22799 30104
rect 22612 30064 22618 30076
rect 22787 30073 22799 30076
rect 22833 30073 22845 30107
rect 22787 30067 22845 30073
rect 22922 30064 22928 30116
rect 22980 30104 22986 30116
rect 22980 30076 23025 30104
rect 22980 30064 22986 30076
rect 23290 30064 23296 30116
rect 23348 30104 23354 30116
rect 27632 30104 27660 30203
rect 27706 30132 27712 30184
rect 27764 30172 27770 30184
rect 27764 30144 27809 30172
rect 27764 30132 27770 30144
rect 23348 30076 27660 30104
rect 28092 30104 28120 30280
rect 28166 30268 28172 30320
rect 28224 30308 28230 30320
rect 31018 30308 31024 30320
rect 28224 30280 31024 30308
rect 28224 30268 28230 30280
rect 28350 30240 28356 30252
rect 28311 30212 28356 30240
rect 28350 30200 28356 30212
rect 28408 30200 28414 30252
rect 28500 30243 28558 30249
rect 28500 30209 28512 30243
rect 28546 30240 28558 30243
rect 28902 30240 28908 30252
rect 28546 30212 28908 30240
rect 28546 30209 28558 30212
rect 28500 30203 28558 30209
rect 28902 30200 28908 30212
rect 28960 30200 28966 30252
rect 29638 30200 29644 30252
rect 29696 30240 29702 30252
rect 29841 30249 29869 30280
rect 31018 30268 31024 30280
rect 31076 30268 31082 30320
rect 31386 30268 31392 30320
rect 31444 30308 31450 30320
rect 34054 30317 34060 30320
rect 34048 30308 34060 30317
rect 31444 30280 31489 30308
rect 34015 30280 34060 30308
rect 31444 30268 31450 30280
rect 34048 30271 34060 30280
rect 34054 30268 34060 30271
rect 34112 30268 34118 30320
rect 29733 30243 29791 30249
rect 29733 30240 29745 30243
rect 29696 30212 29745 30240
rect 29696 30200 29702 30212
rect 29733 30209 29745 30212
rect 29779 30209 29791 30243
rect 29733 30203 29791 30209
rect 29826 30243 29884 30249
rect 29826 30209 29838 30243
rect 29872 30209 29884 30243
rect 30006 30240 30012 30252
rect 29967 30212 30012 30240
rect 29826 30203 29884 30209
rect 30006 30200 30012 30212
rect 30064 30200 30070 30252
rect 30282 30249 30288 30252
rect 30101 30243 30159 30249
rect 30101 30209 30113 30243
rect 30147 30209 30159 30243
rect 30101 30203 30159 30209
rect 30239 30243 30288 30249
rect 30239 30209 30251 30243
rect 30285 30209 30288 30243
rect 30239 30203 30288 30209
rect 28718 30172 28724 30184
rect 28679 30144 28724 30172
rect 28718 30132 28724 30144
rect 28776 30132 28782 30184
rect 29362 30104 29368 30116
rect 28092 30076 29368 30104
rect 23348 30064 23354 30076
rect 24688 30048 24716 30076
rect 29362 30064 29368 30076
rect 29420 30064 29426 30116
rect 30116 30104 30144 30203
rect 30282 30200 30288 30203
rect 30340 30200 30346 30252
rect 30466 30200 30472 30252
rect 30524 30240 30530 30252
rect 30745 30243 30803 30249
rect 30745 30240 30757 30243
rect 30524 30212 30757 30240
rect 30524 30200 30530 30212
rect 30745 30209 30757 30212
rect 30791 30209 30803 30243
rect 31110 30240 31116 30252
rect 31071 30212 31116 30240
rect 30745 30203 30803 30209
rect 30760 30172 30788 30203
rect 31110 30200 31116 30212
rect 31168 30200 31174 30252
rect 31294 30249 31300 30252
rect 31261 30243 31300 30249
rect 31261 30209 31273 30243
rect 31261 30203 31300 30209
rect 31294 30200 31300 30203
rect 31352 30200 31358 30252
rect 31481 30243 31539 30249
rect 31481 30209 31493 30243
rect 31527 30209 31539 30243
rect 31481 30203 31539 30209
rect 31018 30172 31024 30184
rect 30760 30144 31024 30172
rect 31018 30132 31024 30144
rect 31076 30172 31082 30184
rect 31496 30172 31524 30203
rect 31570 30200 31576 30252
rect 31628 30249 31634 30252
rect 31628 30240 31636 30249
rect 31628 30212 31673 30240
rect 31628 30203 31636 30212
rect 31628 30200 31634 30203
rect 31076 30144 31524 30172
rect 31076 30132 31082 30144
rect 32214 30132 32220 30184
rect 32272 30172 32278 30184
rect 32766 30172 32772 30184
rect 32272 30144 32772 30172
rect 32272 30132 32278 30144
rect 32766 30132 32772 30144
rect 32824 30172 32830 30184
rect 33781 30175 33839 30181
rect 33781 30172 33793 30175
rect 32824 30144 33793 30172
rect 32824 30132 32830 30144
rect 33781 30141 33793 30144
rect 33827 30141 33839 30175
rect 33781 30135 33839 30141
rect 30374 30104 30380 30116
rect 30116 30076 30380 30104
rect 30374 30064 30380 30076
rect 30432 30104 30438 30116
rect 31846 30104 31852 30116
rect 30432 30076 31852 30104
rect 30432 30064 30438 30076
rect 31846 30064 31852 30076
rect 31904 30064 31910 30116
rect 35176 30104 35204 30339
rect 35894 30336 35900 30388
rect 35952 30376 35958 30388
rect 36449 30379 36507 30385
rect 35952 30348 36313 30376
rect 35952 30336 35958 30348
rect 36170 30308 36176 30320
rect 36131 30280 36176 30308
rect 36170 30268 36176 30280
rect 36228 30268 36234 30320
rect 36285 30252 36313 30348
rect 36449 30345 36461 30379
rect 36495 30345 36507 30379
rect 37826 30376 37832 30388
rect 37787 30348 37832 30376
rect 36449 30339 36507 30345
rect 36464 30308 36492 30339
rect 37826 30336 37832 30348
rect 37884 30336 37890 30388
rect 36722 30308 36728 30320
rect 36464 30280 36728 30308
rect 36722 30268 36728 30280
rect 36780 30308 36786 30320
rect 37921 30311 37979 30317
rect 37921 30308 37933 30311
rect 36780 30280 37933 30308
rect 36780 30268 36786 30280
rect 37921 30277 37933 30280
rect 37967 30277 37979 30311
rect 37921 30271 37979 30277
rect 35802 30240 35808 30252
rect 35763 30212 35808 30240
rect 35802 30200 35808 30212
rect 35860 30200 35866 30252
rect 35894 30200 35900 30252
rect 35952 30240 35958 30252
rect 35952 30212 35997 30240
rect 35952 30200 35958 30212
rect 36078 30200 36084 30252
rect 36136 30240 36142 30252
rect 36136 30212 36181 30240
rect 36136 30200 36142 30212
rect 36262 30200 36268 30252
rect 36320 30249 36326 30252
rect 36320 30240 36328 30249
rect 36320 30212 36413 30240
rect 36320 30203 36328 30212
rect 36320 30200 36326 30203
rect 38010 30172 38016 30184
rect 37971 30144 38016 30172
rect 38010 30132 38016 30144
rect 38068 30132 38074 30184
rect 36078 30104 36084 30116
rect 35176 30076 36084 30104
rect 36078 30064 36084 30076
rect 36136 30064 36142 30116
rect 24302 30036 24308 30048
rect 22480 30008 24308 30036
rect 24302 29996 24308 30008
rect 24360 29996 24366 30048
rect 24670 29996 24676 30048
rect 24728 29996 24734 30048
rect 25498 30036 25504 30048
rect 25459 30008 25504 30036
rect 25498 29996 25504 30008
rect 25556 29996 25562 30048
rect 28626 30036 28632 30048
rect 28587 30008 28632 30036
rect 28626 29996 28632 30008
rect 28684 29996 28690 30048
rect 28997 30039 29055 30045
rect 28997 30005 29009 30039
rect 29043 30036 29055 30039
rect 29454 30036 29460 30048
rect 29043 30008 29460 30036
rect 29043 30005 29055 30008
rect 28997 29999 29055 30005
rect 29454 29996 29460 30008
rect 29512 29996 29518 30048
rect 31386 29996 31392 30048
rect 31444 30036 31450 30048
rect 31570 30036 31576 30048
rect 31444 30008 31576 30036
rect 31444 29996 31450 30008
rect 31570 29996 31576 30008
rect 31628 29996 31634 30048
rect 31757 30039 31815 30045
rect 31757 30005 31769 30039
rect 31803 30036 31815 30039
rect 32398 30036 32404 30048
rect 31803 30008 32404 30036
rect 31803 30005 31815 30008
rect 31757 29999 31815 30005
rect 32398 29996 32404 30008
rect 32456 29996 32462 30048
rect 37458 30036 37464 30048
rect 37419 30008 37464 30036
rect 37458 29996 37464 30008
rect 37516 29996 37522 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 3970 29832 3976 29844
rect 3931 29804 3976 29832
rect 3970 29792 3976 29804
rect 4028 29792 4034 29844
rect 6362 29792 6368 29844
rect 6420 29832 6426 29844
rect 8754 29832 8760 29844
rect 6420 29804 8760 29832
rect 6420 29792 6426 29804
rect 8754 29792 8760 29804
rect 8812 29792 8818 29844
rect 9030 29792 9036 29844
rect 9088 29832 9094 29844
rect 10413 29835 10471 29841
rect 10413 29832 10425 29835
rect 9088 29804 10425 29832
rect 9088 29792 9094 29804
rect 10413 29801 10425 29804
rect 10459 29801 10471 29835
rect 10413 29795 10471 29801
rect 10502 29792 10508 29844
rect 10560 29832 10566 29844
rect 11790 29832 11796 29844
rect 10560 29804 11560 29832
rect 11751 29804 11796 29832
rect 10560 29792 10566 29804
rect 5258 29764 5264 29776
rect 3252 29736 5264 29764
rect 3252 29637 3280 29736
rect 5258 29724 5264 29736
rect 5316 29724 5322 29776
rect 6270 29764 6276 29776
rect 5368 29736 6276 29764
rect 4154 29656 4160 29708
rect 4212 29696 4218 29708
rect 4525 29699 4583 29705
rect 4525 29696 4537 29699
rect 4212 29668 4537 29696
rect 4212 29656 4218 29668
rect 4525 29665 4537 29668
rect 4571 29696 4583 29699
rect 5074 29696 5080 29708
rect 4571 29668 5080 29696
rect 4571 29665 4583 29668
rect 4525 29659 4583 29665
rect 5074 29656 5080 29668
rect 5132 29656 5138 29708
rect 5368 29696 5396 29736
rect 6270 29724 6276 29736
rect 6328 29724 6334 29776
rect 6546 29724 6552 29776
rect 6604 29764 6610 29776
rect 11425 29767 11483 29773
rect 11425 29764 11437 29767
rect 6604 29736 11437 29764
rect 6604 29724 6610 29736
rect 11425 29733 11437 29736
rect 11471 29733 11483 29767
rect 11532 29764 11560 29804
rect 11790 29792 11796 29804
rect 11848 29792 11854 29844
rect 11977 29835 12035 29841
rect 11977 29801 11989 29835
rect 12023 29832 12035 29835
rect 12250 29832 12256 29844
rect 12023 29804 12256 29832
rect 12023 29801 12035 29804
rect 11977 29795 12035 29801
rect 12250 29792 12256 29804
rect 12308 29792 12314 29844
rect 12437 29835 12495 29841
rect 12437 29801 12449 29835
rect 12483 29801 12495 29835
rect 12437 29795 12495 29801
rect 12728 29804 13216 29832
rect 12066 29764 12072 29776
rect 11532 29736 12072 29764
rect 11425 29727 11483 29733
rect 5626 29696 5632 29708
rect 5184 29668 5396 29696
rect 5587 29668 5632 29696
rect 3237 29631 3295 29637
rect 3237 29597 3249 29631
rect 3283 29597 3295 29631
rect 3237 29591 3295 29597
rect 3421 29631 3479 29637
rect 3421 29597 3433 29631
rect 3467 29597 3479 29631
rect 3421 29591 3479 29597
rect 4341 29631 4399 29637
rect 4341 29597 4353 29631
rect 4387 29628 4399 29631
rect 4614 29628 4620 29640
rect 4387 29600 4620 29628
rect 4387 29597 4399 29600
rect 4341 29591 4399 29597
rect 3436 29560 3464 29591
rect 4614 29588 4620 29600
rect 4672 29588 4678 29640
rect 5184 29560 5212 29668
rect 5626 29656 5632 29668
rect 5684 29696 5690 29708
rect 5994 29696 6000 29708
rect 5684 29668 6000 29696
rect 5684 29656 5690 29668
rect 5994 29656 6000 29668
rect 6052 29656 6058 29708
rect 6730 29696 6736 29708
rect 6104 29668 6736 29696
rect 5350 29628 5356 29640
rect 5311 29600 5356 29628
rect 5350 29588 5356 29600
rect 5408 29588 5414 29640
rect 5442 29588 5448 29640
rect 5500 29628 5506 29640
rect 6104 29637 6132 29668
rect 6730 29656 6736 29668
rect 6788 29656 6794 29708
rect 7650 29696 7656 29708
rect 7300 29668 7656 29696
rect 5537 29631 5595 29637
rect 5537 29628 5549 29631
rect 5500 29600 5549 29628
rect 5500 29588 5506 29600
rect 5537 29597 5549 29600
rect 5583 29597 5595 29631
rect 5537 29591 5595 29597
rect 6089 29631 6147 29637
rect 6089 29597 6101 29631
rect 6135 29597 6147 29631
rect 6089 29591 6147 29597
rect 6273 29631 6331 29637
rect 6273 29597 6285 29631
rect 6319 29628 6331 29631
rect 6638 29628 6644 29640
rect 6319 29600 6644 29628
rect 6319 29597 6331 29600
rect 6273 29591 6331 29597
rect 3436 29532 5212 29560
rect 5258 29520 5264 29572
rect 5316 29560 5322 29572
rect 6288 29560 6316 29591
rect 6638 29588 6644 29600
rect 6696 29588 6702 29640
rect 7006 29628 7012 29640
rect 6967 29600 7012 29628
rect 7006 29588 7012 29600
rect 7064 29588 7070 29640
rect 7098 29588 7104 29640
rect 7156 29628 7162 29640
rect 7300 29637 7328 29668
rect 7650 29656 7656 29668
rect 7708 29656 7714 29708
rect 11440 29696 11468 29727
rect 12066 29724 12072 29736
rect 12124 29764 12130 29776
rect 12452 29764 12480 29795
rect 12124 29736 12480 29764
rect 12124 29724 12130 29736
rect 12728 29696 12756 29804
rect 12805 29767 12863 29773
rect 12805 29733 12817 29767
rect 12851 29733 12863 29767
rect 13188 29764 13216 29804
rect 15470 29792 15476 29844
rect 15528 29832 15534 29844
rect 15933 29835 15991 29841
rect 15933 29832 15945 29835
rect 15528 29804 15945 29832
rect 15528 29792 15534 29804
rect 15933 29801 15945 29804
rect 15979 29801 15991 29835
rect 15933 29795 15991 29801
rect 17313 29835 17371 29841
rect 17313 29801 17325 29835
rect 17359 29801 17371 29835
rect 17770 29832 17776 29844
rect 17731 29804 17776 29832
rect 17313 29795 17371 29801
rect 14458 29764 14464 29776
rect 13188 29736 14464 29764
rect 12805 29727 12863 29733
rect 11440 29668 12756 29696
rect 7285 29631 7343 29637
rect 7285 29628 7297 29631
rect 7156 29600 7297 29628
rect 7156 29588 7162 29600
rect 7285 29597 7297 29600
rect 7331 29597 7343 29631
rect 7285 29591 7343 29597
rect 7561 29631 7619 29637
rect 7561 29597 7573 29631
rect 7607 29597 7619 29631
rect 7561 29591 7619 29597
rect 7745 29631 7803 29637
rect 7745 29597 7757 29631
rect 7791 29628 7803 29631
rect 8110 29628 8116 29640
rect 7791 29600 8116 29628
rect 7791 29597 7803 29600
rect 7745 29591 7803 29597
rect 5316 29532 6316 29560
rect 5316 29520 5322 29532
rect 6362 29520 6368 29572
rect 6420 29560 6426 29572
rect 7576 29560 7604 29591
rect 8110 29588 8116 29600
rect 8168 29588 8174 29640
rect 9214 29628 9220 29640
rect 8220 29600 9220 29628
rect 7834 29560 7840 29572
rect 6420 29532 7840 29560
rect 6420 29520 6426 29532
rect 7834 29520 7840 29532
rect 7892 29560 7898 29572
rect 8220 29560 8248 29600
rect 9214 29588 9220 29600
rect 9272 29588 9278 29640
rect 9950 29588 9956 29640
rect 10008 29628 10014 29640
rect 11974 29628 11980 29640
rect 10008 29600 11980 29628
rect 10008 29588 10014 29600
rect 11974 29588 11980 29600
rect 12032 29628 12038 29640
rect 12437 29631 12495 29637
rect 12437 29628 12449 29631
rect 12032 29600 12449 29628
rect 12032 29588 12038 29600
rect 12437 29597 12449 29600
rect 12483 29597 12495 29631
rect 12437 29591 12495 29597
rect 12526 29588 12532 29640
rect 12584 29628 12590 29640
rect 12820 29628 12848 29727
rect 14458 29724 14464 29736
rect 14516 29724 14522 29776
rect 15654 29724 15660 29776
rect 15712 29764 15718 29776
rect 17328 29764 17356 29795
rect 17770 29792 17776 29804
rect 17828 29792 17834 29844
rect 20257 29835 20315 29841
rect 20257 29801 20269 29835
rect 20303 29832 20315 29835
rect 22094 29832 22100 29844
rect 20303 29804 22100 29832
rect 20303 29801 20315 29804
rect 20257 29795 20315 29801
rect 22094 29792 22100 29804
rect 22152 29792 22158 29844
rect 22186 29792 22192 29844
rect 22244 29832 22250 29844
rect 22281 29835 22339 29841
rect 22281 29832 22293 29835
rect 22244 29804 22293 29832
rect 22244 29792 22250 29804
rect 22281 29801 22293 29804
rect 22327 29801 22339 29835
rect 23382 29832 23388 29844
rect 23343 29804 23388 29832
rect 22281 29795 22339 29801
rect 23382 29792 23388 29804
rect 23440 29792 23446 29844
rect 25961 29835 26019 29841
rect 25961 29801 25973 29835
rect 26007 29832 26019 29835
rect 26050 29832 26056 29844
rect 26007 29804 26056 29832
rect 26007 29801 26019 29804
rect 25961 29795 26019 29801
rect 26050 29792 26056 29804
rect 26108 29832 26114 29844
rect 26418 29832 26424 29844
rect 26108 29804 26424 29832
rect 26108 29792 26114 29804
rect 26418 29792 26424 29804
rect 26476 29792 26482 29844
rect 26510 29792 26516 29844
rect 26568 29832 26574 29844
rect 30469 29835 30527 29841
rect 26568 29804 28994 29832
rect 26568 29792 26574 29804
rect 15712 29736 17356 29764
rect 15712 29724 15718 29736
rect 20714 29724 20720 29776
rect 20772 29764 20778 29776
rect 21269 29767 21327 29773
rect 21269 29764 21281 29767
rect 20772 29736 21281 29764
rect 20772 29724 20778 29736
rect 21269 29733 21281 29736
rect 21315 29764 21327 29767
rect 22646 29764 22652 29776
rect 21315 29736 22652 29764
rect 21315 29733 21327 29736
rect 21269 29727 21327 29733
rect 22646 29724 22652 29736
rect 22704 29724 22710 29776
rect 22833 29767 22891 29773
rect 22833 29733 22845 29767
rect 22879 29764 22891 29767
rect 28350 29764 28356 29776
rect 22879 29736 28356 29764
rect 22879 29733 22891 29736
rect 22833 29727 22891 29733
rect 28350 29724 28356 29736
rect 28408 29724 28414 29776
rect 28966 29764 28994 29804
rect 30469 29801 30481 29835
rect 30515 29832 30527 29835
rect 30742 29832 30748 29844
rect 30515 29804 30748 29832
rect 30515 29801 30527 29804
rect 30469 29795 30527 29801
rect 30742 29792 30748 29804
rect 30800 29792 30806 29844
rect 31726 29804 35296 29832
rect 30650 29764 30656 29776
rect 28966 29736 30656 29764
rect 30650 29724 30656 29736
rect 30708 29724 30714 29776
rect 14274 29656 14280 29708
rect 14332 29696 14338 29708
rect 15013 29699 15071 29705
rect 15013 29696 15025 29699
rect 14332 29668 15025 29696
rect 14332 29656 14338 29668
rect 15013 29665 15025 29668
rect 15059 29665 15071 29699
rect 15013 29659 15071 29665
rect 15378 29656 15384 29708
rect 15436 29696 15442 29708
rect 17405 29699 17463 29705
rect 17405 29696 17417 29699
rect 15436 29668 17417 29696
rect 15436 29656 15442 29668
rect 17405 29665 17417 29668
rect 17451 29696 17463 29699
rect 18230 29696 18236 29708
rect 17451 29668 18236 29696
rect 17451 29665 17463 29668
rect 17405 29659 17463 29665
rect 18230 29656 18236 29668
rect 18288 29656 18294 29708
rect 19978 29656 19984 29708
rect 20036 29696 20042 29708
rect 20036 29668 20760 29696
rect 20036 29656 20042 29668
rect 13265 29631 13323 29637
rect 13265 29628 13277 29631
rect 12584 29600 12629 29628
rect 12820 29600 13277 29628
rect 12584 29588 12590 29600
rect 7892 29532 8248 29560
rect 9125 29563 9183 29569
rect 7892 29520 7898 29532
rect 9125 29529 9137 29563
rect 9171 29560 9183 29563
rect 11698 29560 11704 29572
rect 9171 29532 11704 29560
rect 9171 29529 9183 29532
rect 9125 29523 9183 29529
rect 11698 29520 11704 29532
rect 11756 29520 11762 29572
rect 11793 29563 11851 29569
rect 11793 29529 11805 29563
rect 11839 29560 11851 29563
rect 12820 29560 12848 29600
rect 13265 29597 13277 29600
rect 13311 29597 13323 29631
rect 13265 29591 13323 29597
rect 13354 29588 13360 29640
rect 13412 29628 13418 29640
rect 13449 29631 13507 29637
rect 13449 29628 13461 29631
rect 13412 29600 13461 29628
rect 13412 29588 13418 29600
rect 13449 29597 13461 29600
rect 13495 29597 13507 29631
rect 13449 29591 13507 29597
rect 13906 29588 13912 29640
rect 13964 29628 13970 29640
rect 15746 29628 15752 29640
rect 13964 29600 15752 29628
rect 13964 29588 13970 29600
rect 15746 29588 15752 29600
rect 15804 29588 15810 29640
rect 15841 29631 15899 29637
rect 15841 29597 15853 29631
rect 15887 29628 15899 29631
rect 16482 29628 16488 29640
rect 15887 29600 16488 29628
rect 15887 29597 15899 29600
rect 15841 29591 15899 29597
rect 16482 29588 16488 29600
rect 16540 29588 16546 29640
rect 16577 29631 16635 29637
rect 16577 29597 16589 29631
rect 16623 29597 16635 29631
rect 16577 29591 16635 29597
rect 16761 29631 16819 29637
rect 16761 29597 16773 29631
rect 16807 29628 16819 29631
rect 16850 29628 16856 29640
rect 16807 29600 16856 29628
rect 16807 29597 16819 29600
rect 16761 29591 16819 29597
rect 11839 29532 12848 29560
rect 11839 29529 11851 29532
rect 11793 29523 11851 29529
rect 13170 29520 13176 29572
rect 13228 29560 13234 29572
rect 14277 29563 14335 29569
rect 14277 29560 14289 29563
rect 13228 29532 14289 29560
rect 13228 29520 13234 29532
rect 14277 29529 14289 29532
rect 14323 29560 14335 29563
rect 16022 29560 16028 29572
rect 14323 29532 16028 29560
rect 14323 29529 14335 29532
rect 14277 29523 14335 29529
rect 16022 29520 16028 29532
rect 16080 29520 16086 29572
rect 16592 29560 16620 29591
rect 16850 29588 16856 29600
rect 16908 29588 16914 29640
rect 17589 29631 17647 29637
rect 17589 29597 17601 29631
rect 17635 29628 17647 29631
rect 17770 29628 17776 29640
rect 17635 29600 17776 29628
rect 17635 29597 17647 29600
rect 17589 29591 17647 29597
rect 17770 29588 17776 29600
rect 17828 29588 17834 29640
rect 20254 29588 20260 29640
rect 20312 29628 20318 29640
rect 20441 29631 20499 29637
rect 20441 29628 20453 29631
rect 20312 29600 20453 29628
rect 20312 29588 20318 29600
rect 20441 29597 20453 29600
rect 20487 29597 20499 29631
rect 20622 29628 20628 29640
rect 20583 29600 20628 29628
rect 20441 29591 20499 29597
rect 20622 29588 20628 29600
rect 20680 29588 20686 29640
rect 20732 29637 20760 29668
rect 21358 29656 21364 29708
rect 21416 29696 21422 29708
rect 21453 29699 21511 29705
rect 21453 29696 21465 29699
rect 21416 29668 21465 29696
rect 21416 29656 21422 29668
rect 21453 29665 21465 29668
rect 21499 29696 21511 29699
rect 22002 29696 22008 29708
rect 21499 29668 22008 29696
rect 21499 29665 21511 29668
rect 21453 29659 21511 29665
rect 22002 29656 22008 29668
rect 22060 29696 22066 29708
rect 22465 29699 22523 29705
rect 22060 29668 22232 29696
rect 22060 29656 22066 29668
rect 20717 29631 20775 29637
rect 20717 29597 20729 29631
rect 20763 29597 20775 29631
rect 21174 29628 21180 29640
rect 21135 29600 21180 29628
rect 20717 29591 20775 29597
rect 21174 29588 21180 29600
rect 21232 29588 21238 29640
rect 22204 29637 22232 29668
rect 22465 29665 22477 29699
rect 22511 29696 22523 29699
rect 24118 29696 24124 29708
rect 22511 29668 24124 29696
rect 22511 29665 22523 29668
rect 22465 29659 22523 29665
rect 24118 29656 24124 29668
rect 24176 29656 24182 29708
rect 27341 29699 27399 29705
rect 27341 29696 27353 29699
rect 24688 29668 27353 29696
rect 22194 29631 22252 29637
rect 22194 29597 22206 29631
rect 22240 29597 22252 29631
rect 22194 29591 22252 29597
rect 22554 29588 22560 29640
rect 22612 29628 22618 29640
rect 22649 29631 22707 29637
rect 22649 29628 22661 29631
rect 22612 29600 22661 29628
rect 22612 29588 22618 29600
rect 22649 29597 22661 29600
rect 22695 29597 22707 29631
rect 22649 29591 22707 29597
rect 23014 29588 23020 29640
rect 23072 29628 23078 29640
rect 23293 29631 23351 29637
rect 23293 29628 23305 29631
rect 23072 29600 23305 29628
rect 23072 29588 23078 29600
rect 23293 29597 23305 29600
rect 23339 29597 23351 29631
rect 23293 29591 23351 29597
rect 23382 29588 23388 29640
rect 23440 29628 23446 29640
rect 23477 29631 23535 29637
rect 23477 29628 23489 29631
rect 23440 29600 23489 29628
rect 23440 29588 23446 29600
rect 23477 29597 23489 29600
rect 23523 29597 23535 29631
rect 23477 29591 23535 29597
rect 23658 29588 23664 29640
rect 23716 29628 23722 29640
rect 24581 29631 24639 29637
rect 24581 29628 24593 29631
rect 23716 29600 24593 29628
rect 23716 29588 23722 29600
rect 24581 29597 24593 29600
rect 24627 29597 24639 29631
rect 24581 29591 24639 29597
rect 17310 29560 17316 29572
rect 16592 29532 16804 29560
rect 17271 29532 17316 29560
rect 16776 29504 16804 29532
rect 17310 29520 17316 29532
rect 17368 29520 17374 29572
rect 18322 29520 18328 29572
rect 18380 29560 18386 29572
rect 19242 29560 19248 29572
rect 18380 29532 19248 29560
rect 18380 29520 18386 29532
rect 19242 29520 19248 29532
rect 19300 29520 19306 29572
rect 20530 29520 20536 29572
rect 20588 29560 20594 29572
rect 24688 29560 24716 29668
rect 27341 29665 27353 29668
rect 27387 29696 27399 29699
rect 27706 29696 27712 29708
rect 27387 29668 27712 29696
rect 27387 29665 27399 29668
rect 27341 29659 27399 29665
rect 27706 29656 27712 29668
rect 27764 29656 27770 29708
rect 24765 29631 24823 29637
rect 24765 29597 24777 29631
rect 24811 29628 24823 29631
rect 25038 29628 25044 29640
rect 24811 29600 25044 29628
rect 24811 29597 24823 29600
rect 24765 29591 24823 29597
rect 25038 29588 25044 29600
rect 25096 29628 25102 29640
rect 25498 29628 25504 29640
rect 25096 29600 25504 29628
rect 25096 29588 25102 29600
rect 25498 29588 25504 29600
rect 25556 29628 25562 29640
rect 26878 29628 26884 29640
rect 25556 29600 26740 29628
rect 26839 29600 26884 29628
rect 25556 29588 25562 29600
rect 20588 29532 24716 29560
rect 25777 29563 25835 29569
rect 20588 29520 20594 29532
rect 25777 29529 25789 29563
rect 25823 29529 25835 29563
rect 26712 29560 26740 29600
rect 26878 29588 26884 29600
rect 26936 29588 26942 29640
rect 27065 29631 27123 29637
rect 27065 29597 27077 29631
rect 27111 29597 27123 29631
rect 27065 29591 27123 29597
rect 27080 29560 27108 29591
rect 27522 29588 27528 29640
rect 27580 29628 27586 29640
rect 28261 29631 28319 29637
rect 28261 29628 28273 29631
rect 27580 29600 28273 29628
rect 27580 29588 27586 29600
rect 28261 29597 28273 29600
rect 28307 29597 28319 29631
rect 28261 29591 28319 29597
rect 29638 29588 29644 29640
rect 29696 29628 29702 29640
rect 30006 29637 30012 29640
rect 29825 29631 29883 29637
rect 29825 29628 29837 29631
rect 29696 29600 29837 29628
rect 29696 29588 29702 29600
rect 29825 29597 29837 29600
rect 29871 29597 29883 29631
rect 29825 29591 29883 29597
rect 29973 29631 30012 29637
rect 29973 29597 29985 29631
rect 29973 29591 30012 29597
rect 30006 29588 30012 29591
rect 30064 29588 30070 29640
rect 30098 29588 30104 29640
rect 30156 29628 30162 29640
rect 30374 29637 30380 29640
rect 30331 29631 30380 29637
rect 30156 29600 30201 29628
rect 30156 29588 30162 29600
rect 30331 29597 30343 29631
rect 30377 29597 30380 29631
rect 30331 29591 30380 29597
rect 30374 29588 30380 29591
rect 30432 29588 30438 29640
rect 31726 29628 31754 29804
rect 32401 29767 32459 29773
rect 32401 29733 32413 29767
rect 32447 29733 32459 29767
rect 32401 29727 32459 29733
rect 31849 29699 31907 29705
rect 31849 29665 31861 29699
rect 31895 29696 31907 29699
rect 32214 29696 32220 29708
rect 31895 29668 32220 29696
rect 31895 29665 31907 29668
rect 31849 29659 31907 29665
rect 32214 29656 32220 29668
rect 32272 29656 32278 29708
rect 32416 29696 32444 29727
rect 32582 29724 32588 29776
rect 32640 29764 32646 29776
rect 32640 29736 33364 29764
rect 32640 29724 32646 29736
rect 32416 29668 33180 29696
rect 32398 29628 32404 29640
rect 30484 29600 31754 29628
rect 32359 29600 32404 29628
rect 26712 29532 27108 29560
rect 25777 29523 25835 29529
rect 3326 29492 3332 29504
rect 3287 29464 3332 29492
rect 3326 29452 3332 29464
rect 3384 29452 3390 29504
rect 4433 29495 4491 29501
rect 4433 29461 4445 29495
rect 4479 29492 4491 29495
rect 5169 29495 5227 29501
rect 5169 29492 5181 29495
rect 4479 29464 5181 29492
rect 4479 29461 4491 29464
rect 4433 29455 4491 29461
rect 5169 29461 5181 29464
rect 5215 29461 5227 29495
rect 6178 29492 6184 29504
rect 6139 29464 6184 29492
rect 5169 29455 5227 29461
rect 6178 29452 6184 29464
rect 6236 29492 6242 29504
rect 6822 29492 6828 29504
rect 6236 29464 6828 29492
rect 6236 29452 6242 29464
rect 6822 29452 6828 29464
rect 6880 29452 6886 29504
rect 7282 29492 7288 29504
rect 7243 29464 7288 29492
rect 7282 29452 7288 29464
rect 7340 29452 7346 29504
rect 8662 29452 8668 29504
rect 8720 29492 8726 29504
rect 11974 29492 11980 29504
rect 8720 29464 11980 29492
rect 8720 29452 8726 29464
rect 11974 29452 11980 29464
rect 12032 29452 12038 29504
rect 13357 29495 13415 29501
rect 13357 29461 13369 29495
rect 13403 29492 13415 29495
rect 15930 29492 15936 29504
rect 13403 29464 15936 29492
rect 13403 29461 13415 29464
rect 13357 29455 13415 29461
rect 15930 29452 15936 29464
rect 15988 29452 15994 29504
rect 16206 29452 16212 29504
rect 16264 29492 16270 29504
rect 16669 29495 16727 29501
rect 16669 29492 16681 29495
rect 16264 29464 16681 29492
rect 16264 29452 16270 29464
rect 16669 29461 16681 29464
rect 16715 29461 16727 29495
rect 16669 29455 16727 29461
rect 16758 29452 16764 29504
rect 16816 29492 16822 29504
rect 18966 29492 18972 29504
rect 16816 29464 18972 29492
rect 16816 29452 16822 29464
rect 18966 29452 18972 29464
rect 19024 29452 19030 29504
rect 19150 29452 19156 29504
rect 19208 29492 19214 29504
rect 19426 29492 19432 29504
rect 19208 29464 19432 29492
rect 19208 29452 19214 29464
rect 19426 29452 19432 29464
rect 19484 29452 19490 29504
rect 20714 29452 20720 29504
rect 20772 29492 20778 29504
rect 21453 29495 21511 29501
rect 21453 29492 21465 29495
rect 20772 29464 21465 29492
rect 20772 29452 20778 29464
rect 21453 29461 21465 29464
rect 21499 29461 21511 29495
rect 24670 29492 24676 29504
rect 24631 29464 24676 29492
rect 21453 29455 21511 29461
rect 24670 29452 24676 29464
rect 24728 29452 24734 29504
rect 24762 29452 24768 29504
rect 24820 29492 24826 29504
rect 25792 29492 25820 29523
rect 27890 29520 27896 29572
rect 27948 29560 27954 29572
rect 28537 29563 28595 29569
rect 28537 29560 28549 29563
rect 27948 29532 28549 29560
rect 27948 29520 27954 29532
rect 28537 29529 28549 29532
rect 28583 29529 28595 29563
rect 28537 29523 28595 29529
rect 29546 29520 29552 29572
rect 29604 29560 29610 29572
rect 30193 29563 30251 29569
rect 30193 29560 30205 29563
rect 29604 29532 30205 29560
rect 29604 29520 29610 29532
rect 30193 29529 30205 29532
rect 30239 29560 30251 29563
rect 30484 29560 30512 29600
rect 32398 29588 32404 29600
rect 32456 29588 32462 29640
rect 32490 29588 32496 29640
rect 32548 29628 32554 29640
rect 33152 29637 33180 29668
rect 33336 29637 33364 29736
rect 32677 29631 32735 29637
rect 32677 29628 32689 29631
rect 32548 29600 32689 29628
rect 32548 29588 32554 29600
rect 32677 29597 32689 29600
rect 32723 29597 32735 29631
rect 32677 29591 32735 29597
rect 33137 29631 33195 29637
rect 33137 29597 33149 29631
rect 33183 29597 33195 29631
rect 33137 29591 33195 29597
rect 33321 29631 33379 29637
rect 33321 29597 33333 29631
rect 33367 29597 33379 29631
rect 33321 29591 33379 29597
rect 34790 29588 34796 29640
rect 34848 29588 34854 29640
rect 35268 29637 35296 29804
rect 37826 29792 37832 29844
rect 37884 29832 37890 29844
rect 38197 29835 38255 29841
rect 38197 29832 38209 29835
rect 37884 29804 38209 29832
rect 37884 29792 37890 29804
rect 38197 29801 38209 29804
rect 38243 29801 38255 29835
rect 38197 29795 38255 29801
rect 35434 29656 35440 29708
rect 35492 29696 35498 29708
rect 35492 29668 35664 29696
rect 35492 29656 35498 29668
rect 35253 29631 35311 29637
rect 35253 29597 35265 29631
rect 35299 29597 35311 29631
rect 35526 29628 35532 29640
rect 35487 29600 35532 29628
rect 35253 29591 35311 29597
rect 35526 29588 35532 29600
rect 35584 29588 35590 29640
rect 35636 29637 35664 29668
rect 36354 29656 36360 29708
rect 36412 29696 36418 29708
rect 36814 29696 36820 29708
rect 36412 29668 36820 29696
rect 36412 29656 36418 29668
rect 36814 29656 36820 29668
rect 36872 29656 36878 29708
rect 35621 29631 35679 29637
rect 35621 29597 35633 29631
rect 35667 29597 35679 29631
rect 35621 29591 35679 29597
rect 37084 29631 37142 29637
rect 37084 29597 37096 29631
rect 37130 29628 37142 29631
rect 37458 29628 37464 29640
rect 37130 29600 37464 29628
rect 37130 29597 37142 29600
rect 37084 29591 37142 29597
rect 37458 29588 37464 29600
rect 37516 29588 37522 29640
rect 31018 29560 31024 29572
rect 30239 29532 30512 29560
rect 30979 29532 31024 29560
rect 30239 29529 30251 29532
rect 30193 29523 30251 29529
rect 31018 29520 31024 29532
rect 31076 29520 31082 29572
rect 34808 29560 34836 29588
rect 35434 29560 35440 29572
rect 34808 29532 35440 29560
rect 35434 29520 35440 29532
rect 35492 29520 35498 29572
rect 24820 29464 25820 29492
rect 24820 29452 24826 29464
rect 25958 29452 25964 29504
rect 26016 29501 26022 29504
rect 26016 29495 26035 29501
rect 26023 29461 26035 29495
rect 26016 29455 26035 29461
rect 26145 29495 26203 29501
rect 26145 29461 26157 29495
rect 26191 29492 26203 29495
rect 26602 29492 26608 29504
rect 26191 29464 26608 29492
rect 26191 29461 26203 29464
rect 26145 29455 26203 29461
rect 26016 29452 26022 29455
rect 26602 29452 26608 29464
rect 26660 29452 26666 29504
rect 30650 29452 30656 29504
rect 30708 29492 30714 29504
rect 31754 29492 31760 29504
rect 30708 29464 31760 29492
rect 30708 29452 30714 29464
rect 31754 29452 31760 29464
rect 31812 29452 31818 29504
rect 32585 29495 32643 29501
rect 32585 29461 32597 29495
rect 32631 29492 32643 29495
rect 32766 29492 32772 29504
rect 32631 29464 32772 29492
rect 32631 29461 32643 29464
rect 32585 29455 32643 29461
rect 32766 29452 32772 29464
rect 32824 29452 32830 29504
rect 33226 29492 33232 29504
rect 33187 29464 33232 29492
rect 33226 29452 33232 29464
rect 33284 29452 33290 29504
rect 35710 29452 35716 29504
rect 35768 29492 35774 29504
rect 35805 29495 35863 29501
rect 35805 29492 35817 29495
rect 35768 29464 35817 29492
rect 35768 29452 35774 29464
rect 35805 29461 35817 29464
rect 35851 29461 35863 29495
rect 35805 29455 35863 29461
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 5166 29248 5172 29300
rect 5224 29288 5230 29300
rect 10134 29288 10140 29300
rect 5224 29260 10140 29288
rect 5224 29248 5230 29260
rect 3326 29180 3332 29232
rect 3384 29220 3390 29232
rect 4249 29223 4307 29229
rect 4249 29220 4261 29223
rect 3384 29192 4261 29220
rect 3384 29180 3390 29192
rect 4249 29189 4261 29192
rect 4295 29189 4307 29223
rect 4249 29183 4307 29189
rect 4341 29223 4399 29229
rect 4341 29189 4353 29223
rect 4387 29220 4399 29223
rect 4798 29220 4804 29232
rect 4387 29192 4804 29220
rect 4387 29189 4399 29192
rect 4341 29183 4399 29189
rect 4798 29180 4804 29192
rect 4856 29220 4862 29232
rect 5442 29220 5448 29232
rect 4856 29192 5448 29220
rect 4856 29180 4862 29192
rect 5442 29180 5448 29192
rect 5500 29180 5506 29232
rect 7006 29180 7012 29232
rect 7064 29220 7070 29232
rect 7466 29220 7472 29232
rect 7064 29192 7472 29220
rect 7064 29180 7070 29192
rect 7466 29180 7472 29192
rect 7524 29220 7530 29232
rect 8864 29229 8892 29260
rect 10134 29248 10140 29260
rect 10192 29248 10198 29300
rect 10505 29291 10563 29297
rect 10505 29257 10517 29291
rect 10551 29257 10563 29291
rect 11790 29288 11796 29300
rect 11751 29260 11796 29288
rect 10505 29251 10563 29257
rect 7653 29223 7711 29229
rect 7653 29220 7665 29223
rect 7524 29192 7665 29220
rect 7524 29180 7530 29192
rect 7653 29189 7665 29192
rect 7699 29189 7711 29223
rect 7653 29183 7711 29189
rect 8849 29223 8907 29229
rect 8849 29189 8861 29223
rect 8895 29189 8907 29223
rect 10520 29220 10548 29251
rect 11790 29248 11796 29260
rect 11848 29248 11854 29300
rect 15654 29248 15660 29300
rect 15712 29288 15718 29300
rect 15841 29291 15899 29297
rect 15841 29288 15853 29291
rect 15712 29260 15853 29288
rect 15712 29248 15718 29260
rect 15841 29257 15853 29260
rect 15887 29257 15899 29291
rect 17862 29288 17868 29300
rect 15841 29251 15899 29257
rect 16132 29260 17868 29288
rect 16132 29220 16160 29260
rect 17862 29248 17868 29260
rect 17920 29248 17926 29300
rect 19168 29260 19334 29288
rect 10520 29192 16160 29220
rect 8849 29183 8907 29189
rect 16206 29180 16212 29232
rect 16264 29220 16270 29232
rect 19168 29220 19196 29260
rect 16264 29192 17080 29220
rect 16264 29180 16270 29192
rect 4062 29152 4068 29164
rect 4023 29124 4068 29152
rect 4062 29112 4068 29124
rect 4120 29112 4126 29164
rect 4433 29155 4491 29161
rect 4433 29121 4445 29155
rect 4479 29121 4491 29155
rect 4433 29115 4491 29121
rect 4448 29084 4476 29115
rect 4890 29112 4896 29164
rect 4948 29152 4954 29164
rect 5077 29155 5135 29161
rect 5077 29152 5089 29155
rect 4948 29124 5089 29152
rect 4948 29112 4954 29124
rect 5077 29121 5089 29124
rect 5123 29121 5135 29155
rect 5258 29152 5264 29164
rect 5219 29124 5264 29152
rect 5077 29115 5135 29121
rect 5258 29112 5264 29124
rect 5316 29112 5322 29164
rect 7285 29155 7343 29161
rect 7285 29121 7297 29155
rect 7331 29152 7343 29155
rect 7558 29152 7564 29164
rect 7331 29124 7564 29152
rect 7331 29121 7343 29124
rect 7285 29115 7343 29121
rect 7558 29112 7564 29124
rect 7616 29112 7622 29164
rect 8754 29112 8760 29164
rect 8812 29152 8818 29164
rect 9125 29155 9183 29161
rect 9125 29152 9137 29155
rect 8812 29124 9137 29152
rect 8812 29112 8818 29124
rect 9125 29121 9137 29124
rect 9171 29152 9183 29155
rect 9582 29152 9588 29164
rect 9171 29124 9588 29152
rect 9171 29121 9183 29124
rect 9125 29115 9183 29121
rect 9582 29112 9588 29124
rect 9640 29112 9646 29164
rect 9858 29112 9864 29164
rect 9916 29152 9922 29164
rect 10045 29155 10103 29161
rect 10045 29152 10057 29155
rect 9916 29124 10057 29152
rect 9916 29112 9922 29124
rect 10045 29121 10057 29124
rect 10091 29121 10103 29155
rect 10045 29115 10103 29121
rect 10226 29112 10232 29164
rect 10284 29152 10290 29164
rect 10321 29155 10379 29161
rect 10321 29152 10333 29155
rect 10284 29124 10333 29152
rect 10284 29112 10290 29124
rect 10321 29121 10333 29124
rect 10367 29152 10379 29155
rect 11514 29152 11520 29164
rect 10367 29124 11520 29152
rect 10367 29121 10379 29124
rect 10321 29115 10379 29121
rect 11514 29112 11520 29124
rect 11572 29112 11578 29164
rect 11606 29112 11612 29164
rect 11664 29152 11670 29164
rect 11701 29155 11759 29161
rect 11701 29152 11713 29155
rect 11664 29124 11713 29152
rect 11664 29112 11670 29124
rect 11701 29121 11713 29124
rect 11747 29121 11759 29155
rect 11882 29152 11888 29164
rect 11843 29124 11888 29152
rect 11701 29115 11759 29121
rect 11882 29112 11888 29124
rect 11940 29112 11946 29164
rect 12802 29152 12808 29164
rect 12763 29124 12808 29152
rect 12802 29112 12808 29124
rect 12860 29112 12866 29164
rect 13630 29152 13636 29164
rect 13591 29124 13636 29152
rect 13630 29112 13636 29124
rect 13688 29112 13694 29164
rect 16025 29155 16083 29161
rect 16025 29121 16037 29155
rect 16071 29152 16083 29155
rect 16853 29155 16911 29161
rect 16853 29152 16865 29155
rect 16071 29124 16865 29152
rect 16071 29121 16083 29124
rect 16025 29115 16083 29121
rect 16853 29121 16865 29124
rect 16899 29152 16911 29155
rect 16942 29152 16948 29164
rect 16899 29124 16948 29152
rect 16899 29121 16911 29124
rect 16853 29115 16911 29121
rect 16942 29112 16948 29124
rect 17000 29112 17006 29164
rect 17052 29161 17080 29192
rect 17144 29192 19196 29220
rect 19306 29220 19334 29260
rect 19426 29248 19432 29300
rect 19484 29288 19490 29300
rect 19484 29260 19564 29288
rect 19484 29248 19490 29260
rect 19536 29229 19564 29260
rect 22278 29248 22284 29300
rect 22336 29288 22342 29300
rect 22922 29288 22928 29300
rect 22336 29260 22928 29288
rect 22336 29248 22342 29260
rect 22922 29248 22928 29260
rect 22980 29248 22986 29300
rect 23382 29288 23388 29300
rect 23343 29260 23388 29288
rect 23382 29248 23388 29260
rect 23440 29248 23446 29300
rect 23566 29248 23572 29300
rect 23624 29288 23630 29300
rect 24026 29288 24032 29300
rect 23624 29260 24032 29288
rect 23624 29248 23630 29260
rect 24026 29248 24032 29260
rect 24084 29248 24090 29300
rect 24946 29288 24952 29300
rect 24907 29260 24952 29288
rect 24946 29248 24952 29260
rect 25004 29248 25010 29300
rect 25958 29288 25964 29300
rect 25148 29260 25964 29288
rect 19521 29223 19579 29229
rect 19306 29192 19472 29220
rect 17037 29155 17095 29161
rect 17037 29121 17049 29155
rect 17083 29121 17095 29155
rect 17037 29115 17095 29121
rect 5350 29084 5356 29096
rect 4448 29056 5356 29084
rect 5350 29044 5356 29056
rect 5408 29044 5414 29096
rect 9033 29087 9091 29093
rect 9033 29053 9045 29087
rect 9079 29084 9091 29087
rect 9214 29084 9220 29096
rect 9079 29056 9220 29084
rect 9079 29053 9091 29056
rect 9033 29047 9091 29053
rect 9214 29044 9220 29056
rect 9272 29044 9278 29096
rect 9766 29044 9772 29096
rect 9824 29084 9830 29096
rect 10134 29084 10140 29096
rect 9824 29056 10140 29084
rect 9824 29044 9830 29056
rect 10134 29044 10140 29056
rect 10192 29044 10198 29096
rect 12897 29087 12955 29093
rect 12897 29053 12909 29087
rect 12943 29053 12955 29087
rect 12897 29047 12955 29053
rect 4614 29016 4620 29028
rect 4575 28988 4620 29016
rect 4614 28976 4620 28988
rect 4672 28976 4678 29028
rect 4890 28976 4896 29028
rect 4948 29016 4954 29028
rect 7098 29016 7104 29028
rect 4948 28988 7104 29016
rect 4948 28976 4954 28988
rect 7098 28976 7104 28988
rect 7156 28976 7162 29028
rect 9309 29019 9367 29025
rect 9309 28985 9321 29019
rect 9355 29016 9367 29019
rect 11146 29016 11152 29028
rect 9355 28988 11152 29016
rect 9355 28985 9367 28988
rect 9309 28979 9367 28985
rect 11146 28976 11152 28988
rect 11204 28976 11210 29028
rect 12912 29016 12940 29047
rect 14182 29044 14188 29096
rect 14240 29084 14246 29096
rect 14369 29087 14427 29093
rect 14369 29084 14381 29087
rect 14240 29056 14381 29084
rect 14240 29044 14246 29056
rect 14369 29053 14381 29056
rect 14415 29053 14427 29087
rect 14369 29047 14427 29053
rect 14918 29044 14924 29096
rect 14976 29084 14982 29096
rect 16209 29087 16267 29093
rect 16209 29084 16221 29087
rect 14976 29056 16221 29084
rect 14976 29044 14982 29056
rect 16209 29053 16221 29056
rect 16255 29053 16267 29087
rect 16209 29047 16267 29053
rect 13078 29016 13084 29028
rect 12912 28988 13084 29016
rect 13078 28976 13084 28988
rect 13136 28976 13142 29028
rect 13173 29019 13231 29025
rect 13173 28985 13185 29019
rect 13219 29016 13231 29019
rect 14642 29016 14648 29028
rect 13219 28988 14648 29016
rect 13219 28985 13231 28988
rect 13173 28979 13231 28985
rect 14642 28976 14648 28988
rect 14700 28976 14706 29028
rect 16224 29016 16252 29047
rect 16298 29044 16304 29096
rect 16356 29084 16362 29096
rect 16482 29084 16488 29096
rect 16356 29056 16488 29084
rect 16356 29044 16362 29056
rect 16482 29044 16488 29056
rect 16540 29044 16546 29096
rect 17144 29016 17172 29192
rect 19444 29164 19472 29192
rect 19521 29189 19533 29223
rect 19567 29220 19579 29223
rect 21910 29220 21916 29232
rect 19567 29192 21916 29220
rect 19567 29189 19579 29192
rect 19521 29183 19579 29189
rect 21910 29180 21916 29192
rect 21968 29180 21974 29232
rect 17957 29155 18015 29161
rect 17957 29121 17969 29155
rect 18003 29152 18015 29155
rect 18138 29152 18144 29164
rect 18003 29124 18144 29152
rect 18003 29121 18015 29124
rect 17957 29115 18015 29121
rect 18138 29112 18144 29124
rect 18196 29152 18202 29164
rect 18196 29124 19196 29152
rect 18196 29112 18202 29124
rect 17402 29084 17408 29096
rect 17363 29056 17408 29084
rect 17402 29044 17408 29056
rect 17460 29044 17466 29096
rect 18506 29084 18512 29096
rect 18467 29056 18512 29084
rect 18506 29044 18512 29056
rect 18564 29044 18570 29096
rect 18782 29084 18788 29096
rect 18743 29056 18788 29084
rect 18782 29044 18788 29056
rect 18840 29044 18846 29096
rect 19168 29084 19196 29124
rect 19242 29112 19248 29164
rect 19300 29152 19306 29164
rect 19337 29155 19395 29161
rect 19337 29152 19349 29155
rect 19300 29124 19349 29152
rect 19300 29112 19306 29124
rect 19337 29121 19349 29124
rect 19383 29121 19395 29155
rect 19337 29115 19395 29121
rect 19426 29112 19432 29164
rect 19484 29112 19490 29164
rect 19705 29155 19763 29161
rect 19705 29121 19717 29155
rect 19751 29152 19763 29155
rect 20254 29152 20260 29164
rect 19751 29124 20260 29152
rect 19751 29121 19763 29124
rect 19705 29115 19763 29121
rect 20254 29112 20260 29124
rect 20312 29112 20318 29164
rect 20349 29155 20407 29161
rect 20349 29121 20361 29155
rect 20395 29121 20407 29155
rect 20714 29152 20720 29164
rect 20675 29124 20720 29152
rect 20349 29115 20407 29121
rect 19610 29084 19616 29096
rect 19168 29056 19616 29084
rect 19610 29044 19616 29056
rect 19668 29084 19674 29096
rect 19978 29084 19984 29096
rect 19668 29056 19984 29084
rect 19668 29044 19674 29056
rect 19978 29044 19984 29056
rect 20036 29044 20042 29096
rect 20364 29084 20392 29115
rect 20714 29112 20720 29124
rect 20772 29112 20778 29164
rect 22002 29112 22008 29164
rect 22060 29152 22066 29164
rect 22557 29155 22615 29161
rect 22557 29152 22569 29155
rect 22060 29124 22569 29152
rect 22060 29112 22066 29124
rect 22557 29121 22569 29124
rect 22603 29121 22615 29155
rect 22557 29115 22615 29121
rect 22741 29155 22799 29161
rect 22741 29121 22753 29155
rect 22787 29152 22799 29155
rect 23382 29152 23388 29164
rect 22787 29124 23388 29152
rect 22787 29121 22799 29124
rect 22741 29115 22799 29121
rect 23382 29112 23388 29124
rect 23440 29112 23446 29164
rect 23566 29152 23572 29164
rect 23527 29124 23572 29152
rect 23566 29112 23572 29124
rect 23624 29112 23630 29164
rect 23750 29152 23756 29164
rect 23711 29124 23756 29152
rect 23750 29112 23756 29124
rect 23808 29152 23814 29164
rect 24762 29152 24768 29164
rect 23808 29124 24768 29152
rect 23808 29112 23814 29124
rect 24762 29112 24768 29124
rect 24820 29112 24826 29164
rect 25148 29161 25176 29260
rect 25958 29248 25964 29260
rect 26016 29288 26022 29300
rect 26329 29291 26387 29297
rect 26329 29288 26341 29291
rect 26016 29260 26341 29288
rect 26016 29248 26022 29260
rect 26329 29257 26341 29260
rect 26375 29257 26387 29291
rect 30558 29288 30564 29300
rect 26329 29251 26387 29257
rect 28460 29260 30564 29288
rect 25222 29180 25228 29232
rect 25280 29220 25286 29232
rect 26878 29220 26884 29232
rect 25280 29192 26884 29220
rect 25280 29180 25286 29192
rect 26878 29180 26884 29192
rect 26936 29180 26942 29232
rect 27706 29220 27712 29232
rect 27667 29192 27712 29220
rect 27706 29180 27712 29192
rect 27764 29180 27770 29232
rect 25133 29155 25191 29161
rect 25133 29121 25145 29155
rect 25179 29121 25191 29155
rect 25240 29152 25268 29180
rect 25317 29155 25375 29161
rect 25317 29152 25329 29155
rect 25240 29124 25329 29152
rect 25133 29115 25191 29121
rect 25317 29121 25329 29124
rect 25363 29121 25375 29155
rect 25317 29115 25375 29121
rect 25406 29112 25412 29164
rect 25464 29152 25470 29164
rect 25958 29152 25964 29164
rect 25464 29124 25509 29152
rect 25919 29124 25964 29152
rect 25464 29112 25470 29124
rect 25958 29112 25964 29124
rect 26016 29112 26022 29164
rect 27341 29155 27399 29161
rect 27341 29152 27353 29155
rect 26160 29124 27353 29152
rect 21450 29084 21456 29096
rect 20272 29056 21456 29084
rect 20272 29028 20300 29056
rect 21450 29044 21456 29056
rect 21508 29044 21514 29096
rect 22646 29044 22652 29096
rect 22704 29084 22710 29096
rect 23658 29084 23664 29096
rect 22704 29056 23664 29084
rect 22704 29044 22710 29056
rect 23658 29044 23664 29056
rect 23716 29044 23722 29096
rect 23845 29087 23903 29093
rect 23845 29053 23857 29087
rect 23891 29053 23903 29087
rect 23845 29047 23903 29053
rect 16224 28988 17172 29016
rect 18417 29019 18475 29025
rect 18417 28985 18429 29019
rect 18463 29016 18475 29019
rect 19058 29016 19064 29028
rect 18463 28988 19064 29016
rect 18463 28985 18475 28988
rect 18417 28979 18475 28985
rect 19058 28976 19064 28988
rect 19116 28976 19122 29028
rect 20254 28976 20260 29028
rect 20312 28976 20318 29028
rect 20901 29019 20959 29025
rect 20901 28985 20913 29019
rect 20947 29016 20959 29019
rect 22554 29016 22560 29028
rect 20947 28988 22560 29016
rect 20947 28985 20959 28988
rect 20901 28979 20959 28985
rect 22554 28976 22560 28988
rect 22612 28976 22618 29028
rect 22925 29019 22983 29025
rect 22925 28985 22937 29019
rect 22971 29016 22983 29019
rect 23198 29016 23204 29028
rect 22971 28988 23204 29016
rect 22971 28985 22983 28988
rect 22925 28979 22983 28985
rect 23198 28976 23204 28988
rect 23256 28976 23262 29028
rect 3970 28908 3976 28960
rect 4028 28948 4034 28960
rect 4154 28948 4160 28960
rect 4028 28920 4160 28948
rect 4028 28908 4034 28920
rect 4154 28908 4160 28920
rect 4212 28908 4218 28960
rect 4706 28908 4712 28960
rect 4764 28948 4770 28960
rect 5445 28951 5503 28957
rect 5445 28948 5457 28951
rect 4764 28920 5457 28948
rect 4764 28908 4770 28920
rect 5445 28917 5457 28920
rect 5491 28917 5503 28951
rect 5445 28911 5503 28917
rect 6730 28908 6736 28960
rect 6788 28948 6794 28960
rect 8849 28951 8907 28957
rect 8849 28948 8861 28951
rect 6788 28920 8861 28948
rect 6788 28908 6794 28920
rect 8849 28917 8861 28920
rect 8895 28948 8907 28951
rect 9122 28948 9128 28960
rect 8895 28920 9128 28948
rect 8895 28917 8907 28920
rect 8849 28911 8907 28917
rect 9122 28908 9128 28920
rect 9180 28908 9186 28960
rect 9214 28908 9220 28960
rect 9272 28948 9278 28960
rect 10045 28951 10103 28957
rect 10045 28948 10057 28951
rect 9272 28920 10057 28948
rect 9272 28908 9278 28920
rect 10045 28917 10057 28920
rect 10091 28917 10103 28951
rect 10045 28911 10103 28917
rect 12434 28908 12440 28960
rect 12492 28948 12498 28960
rect 12805 28951 12863 28957
rect 12805 28948 12817 28951
rect 12492 28920 12817 28948
rect 12492 28908 12498 28920
rect 12805 28917 12817 28920
rect 12851 28948 12863 28951
rect 15838 28948 15844 28960
rect 12851 28920 15844 28948
rect 12851 28917 12863 28920
rect 12805 28911 12863 28917
rect 15838 28908 15844 28920
rect 15896 28948 15902 28960
rect 16298 28948 16304 28960
rect 15896 28920 16304 28948
rect 15896 28908 15902 28920
rect 16298 28908 16304 28920
rect 16356 28908 16362 28960
rect 18325 28951 18383 28957
rect 18325 28917 18337 28951
rect 18371 28948 18383 28951
rect 19334 28948 19340 28960
rect 18371 28920 19340 28948
rect 18371 28917 18383 28920
rect 18325 28911 18383 28917
rect 19334 28908 19340 28920
rect 19392 28908 19398 28960
rect 20717 28951 20775 28957
rect 20717 28917 20729 28951
rect 20763 28948 20775 28951
rect 20806 28948 20812 28960
rect 20763 28920 20812 28948
rect 20763 28917 20775 28920
rect 20717 28911 20775 28917
rect 20806 28908 20812 28920
rect 20864 28908 20870 28960
rect 21726 28908 21732 28960
rect 21784 28948 21790 28960
rect 22278 28948 22284 28960
rect 21784 28920 22284 28948
rect 21784 28908 21790 28920
rect 22278 28908 22284 28920
rect 22336 28908 22342 28960
rect 23290 28908 23296 28960
rect 23348 28948 23354 28960
rect 23860 28948 23888 29047
rect 24780 29016 24808 29112
rect 25222 29084 25228 29096
rect 25183 29056 25228 29084
rect 25222 29044 25228 29056
rect 25280 29044 25286 29096
rect 25866 29044 25872 29096
rect 25924 29084 25930 29096
rect 26053 29087 26111 29093
rect 26053 29084 26065 29087
rect 25924 29056 26065 29084
rect 25924 29044 25930 29056
rect 26053 29053 26065 29056
rect 26099 29053 26111 29087
rect 26053 29047 26111 29053
rect 26160 29016 26188 29124
rect 27341 29121 27353 29124
rect 27387 29121 27399 29155
rect 27341 29115 27399 29121
rect 27525 29155 27583 29161
rect 27525 29121 27537 29155
rect 27571 29152 27583 29155
rect 27614 29152 27620 29164
rect 27571 29124 27620 29152
rect 27571 29121 27583 29124
rect 27525 29115 27583 29121
rect 27614 29112 27620 29124
rect 27672 29112 27678 29164
rect 28166 29152 28172 29164
rect 28127 29124 28172 29152
rect 28166 29112 28172 29124
rect 28224 29112 28230 29164
rect 28460 29161 28488 29260
rect 30558 29248 30564 29260
rect 30616 29248 30622 29300
rect 32398 29248 32404 29300
rect 32456 29288 32462 29300
rect 32493 29291 32551 29297
rect 32493 29288 32505 29291
rect 32456 29260 32505 29288
rect 32456 29248 32462 29260
rect 32493 29257 32505 29260
rect 32539 29257 32551 29291
rect 32493 29251 32551 29257
rect 32582 29248 32588 29300
rect 32640 29288 32646 29300
rect 32677 29291 32735 29297
rect 32677 29288 32689 29291
rect 32640 29260 32689 29288
rect 32640 29248 32646 29260
rect 32677 29257 32689 29260
rect 32723 29257 32735 29291
rect 32677 29251 32735 29257
rect 36357 29291 36415 29297
rect 36357 29257 36369 29291
rect 36403 29257 36415 29291
rect 36357 29251 36415 29257
rect 29362 29220 29368 29232
rect 29323 29192 29368 29220
rect 29362 29180 29368 29192
rect 29420 29180 29426 29232
rect 30466 29220 30472 29232
rect 30300 29192 30472 29220
rect 28353 29155 28411 29161
rect 28353 29121 28365 29155
rect 28399 29121 28411 29155
rect 28353 29115 28411 29121
rect 28445 29155 28503 29161
rect 28445 29121 28457 29155
rect 28491 29121 28503 29155
rect 28445 29115 28503 29121
rect 28537 29155 28595 29161
rect 28537 29121 28549 29155
rect 28583 29121 28595 29155
rect 29638 29152 29644 29164
rect 29599 29124 29644 29152
rect 28537 29115 28595 29121
rect 27982 29044 27988 29096
rect 28040 29084 28046 29096
rect 28368 29084 28396 29115
rect 28040 29056 28396 29084
rect 28040 29044 28046 29056
rect 24780 28988 26188 29016
rect 27062 28976 27068 29028
rect 27120 29016 27126 29028
rect 27341 29019 27399 29025
rect 27341 29016 27353 29019
rect 27120 28988 27353 29016
rect 27120 28976 27126 28988
rect 27341 28985 27353 28988
rect 27387 29016 27399 29019
rect 27522 29016 27528 29028
rect 27387 28988 27528 29016
rect 27387 28985 27399 28988
rect 27341 28979 27399 28985
rect 27522 28976 27528 28988
rect 27580 28976 27586 29028
rect 28350 28976 28356 29028
rect 28408 29016 28414 29028
rect 28552 29016 28580 29115
rect 29638 29112 29644 29124
rect 29696 29112 29702 29164
rect 29549 29087 29607 29093
rect 29549 29053 29561 29087
rect 29595 29084 29607 29087
rect 30300 29084 30328 29192
rect 30466 29180 30472 29192
rect 30524 29180 30530 29232
rect 30742 29180 30748 29232
rect 30800 29220 30806 29232
rect 32309 29223 32367 29229
rect 30800 29192 30972 29220
rect 30800 29180 30806 29192
rect 30944 29161 30972 29192
rect 32309 29189 32321 29223
rect 32355 29220 32367 29223
rect 32766 29220 32772 29232
rect 32355 29192 32772 29220
rect 32355 29189 32367 29192
rect 32309 29183 32367 29189
rect 32766 29180 32772 29192
rect 32824 29180 32830 29232
rect 33226 29180 33232 29232
rect 33284 29220 33290 29232
rect 33566 29223 33624 29229
rect 33566 29220 33578 29223
rect 33284 29192 33578 29220
rect 33284 29180 33290 29192
rect 33566 29189 33578 29192
rect 33612 29189 33624 29223
rect 36078 29220 36084 29232
rect 36039 29192 36084 29220
rect 33566 29183 33624 29189
rect 36078 29180 36084 29192
rect 36136 29180 36142 29232
rect 30377 29155 30435 29161
rect 30377 29121 30389 29155
rect 30423 29121 30435 29155
rect 30377 29115 30435 29121
rect 30929 29155 30987 29161
rect 30929 29121 30941 29155
rect 30975 29121 30987 29155
rect 30929 29115 30987 29121
rect 29595 29056 30328 29084
rect 29595 29053 29607 29056
rect 29549 29047 29607 29053
rect 28718 29016 28724 29028
rect 28408 28988 28580 29016
rect 28679 28988 28724 29016
rect 28408 28976 28414 28988
rect 28718 28976 28724 28988
rect 28776 28976 28782 29028
rect 29825 29019 29883 29025
rect 29825 28985 29837 29019
rect 29871 29016 29883 29019
rect 30392 29016 30420 29115
rect 31294 29112 31300 29164
rect 31352 29152 31358 29164
rect 31754 29152 31760 29164
rect 31352 29124 31760 29152
rect 31352 29112 31358 29124
rect 31754 29112 31760 29124
rect 31812 29152 31818 29164
rect 35710 29152 35716 29164
rect 31812 29124 34744 29152
rect 35671 29124 35716 29152
rect 31812 29112 31818 29124
rect 30745 29087 30803 29093
rect 30745 29053 30757 29087
rect 30791 29084 30803 29087
rect 31570 29084 31576 29096
rect 30791 29056 31576 29084
rect 30791 29053 30803 29056
rect 30745 29047 30803 29053
rect 31570 29044 31576 29056
rect 31628 29044 31634 29096
rect 33042 29044 33048 29096
rect 33100 29084 33106 29096
rect 33321 29087 33379 29093
rect 33321 29084 33333 29087
rect 33100 29056 33333 29084
rect 33100 29044 33106 29056
rect 33321 29053 33333 29056
rect 33367 29053 33379 29087
rect 33321 29047 33379 29053
rect 34716 29025 34744 29124
rect 35710 29112 35716 29124
rect 35768 29112 35774 29164
rect 35802 29112 35808 29164
rect 35860 29152 35866 29164
rect 35860 29124 35905 29152
rect 35860 29112 35866 29124
rect 35986 29112 35992 29164
rect 36044 29152 36050 29164
rect 36262 29161 36268 29164
rect 36219 29155 36268 29161
rect 36044 29124 36089 29152
rect 36044 29112 36050 29124
rect 36219 29121 36231 29155
rect 36265 29121 36268 29155
rect 36219 29115 36268 29121
rect 36262 29112 36268 29115
rect 36320 29112 36326 29164
rect 36372 29152 36400 29251
rect 37461 29155 37519 29161
rect 37461 29152 37473 29155
rect 36372 29124 37473 29152
rect 37461 29121 37473 29124
rect 37507 29152 37519 29155
rect 37918 29152 37924 29164
rect 37507 29124 37924 29152
rect 37507 29121 37519 29124
rect 37461 29115 37519 29121
rect 37918 29112 37924 29124
rect 37976 29112 37982 29164
rect 37734 29084 37740 29096
rect 37695 29056 37740 29084
rect 37734 29044 37740 29056
rect 37792 29044 37798 29096
rect 29871 28988 30420 29016
rect 34701 29019 34759 29025
rect 29871 28985 29883 28988
rect 29825 28979 29883 28985
rect 34701 28985 34713 29019
rect 34747 29016 34759 29019
rect 36630 29016 36636 29028
rect 34747 28988 36636 29016
rect 34747 28985 34759 28988
rect 34701 28979 34759 28985
rect 36630 28976 36636 28988
rect 36688 28976 36694 29028
rect 25314 28948 25320 28960
rect 23348 28920 25320 28948
rect 23348 28908 23354 28920
rect 25314 28908 25320 28920
rect 25372 28908 25378 28960
rect 26145 28951 26203 28957
rect 26145 28917 26157 28951
rect 26191 28948 26203 28951
rect 26234 28948 26240 28960
rect 26191 28920 26240 28948
rect 26191 28917 26203 28920
rect 26145 28911 26203 28917
rect 26234 28908 26240 28920
rect 26292 28908 26298 28960
rect 29362 28948 29368 28960
rect 29323 28920 29368 28948
rect 29362 28908 29368 28920
rect 29420 28908 29426 28960
rect 32490 28948 32496 28960
rect 32451 28920 32496 28948
rect 32490 28908 32496 28920
rect 32548 28908 32554 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 4617 28747 4675 28753
rect 4617 28713 4629 28747
rect 4663 28744 4675 28747
rect 4798 28744 4804 28756
rect 4663 28716 4804 28744
rect 4663 28713 4675 28716
rect 4617 28707 4675 28713
rect 4798 28704 4804 28716
rect 4856 28704 4862 28756
rect 6178 28744 6184 28756
rect 5184 28716 6184 28744
rect 4525 28543 4583 28549
rect 4525 28509 4537 28543
rect 4571 28540 4583 28543
rect 4706 28540 4712 28552
rect 4571 28512 4712 28540
rect 4571 28509 4583 28512
rect 4525 28503 4583 28509
rect 4706 28500 4712 28512
rect 4764 28500 4770 28552
rect 5184 28549 5212 28716
rect 6178 28704 6184 28716
rect 6236 28704 6242 28756
rect 7374 28704 7380 28756
rect 7432 28744 7438 28756
rect 9214 28744 9220 28756
rect 7432 28716 9220 28744
rect 7432 28704 7438 28716
rect 9214 28704 9220 28716
rect 9272 28704 9278 28756
rect 11054 28744 11060 28756
rect 10967 28716 11060 28744
rect 11054 28704 11060 28716
rect 11112 28744 11118 28756
rect 11882 28744 11888 28756
rect 11112 28716 11888 28744
rect 11112 28704 11118 28716
rect 11882 28704 11888 28716
rect 11940 28704 11946 28756
rect 11974 28704 11980 28756
rect 12032 28744 12038 28756
rect 13998 28744 14004 28756
rect 12032 28716 14004 28744
rect 12032 28704 12038 28716
rect 13998 28704 14004 28716
rect 14056 28704 14062 28756
rect 14826 28744 14832 28756
rect 14787 28716 14832 28744
rect 14826 28704 14832 28716
rect 14884 28704 14890 28756
rect 15562 28704 15568 28756
rect 15620 28744 15626 28756
rect 16117 28747 16175 28753
rect 16117 28744 16129 28747
rect 15620 28716 16129 28744
rect 15620 28704 15626 28716
rect 16117 28713 16129 28716
rect 16163 28713 16175 28747
rect 16850 28744 16856 28756
rect 16117 28707 16175 28713
rect 16408 28716 16856 28744
rect 5534 28636 5540 28688
rect 5592 28676 5598 28688
rect 11241 28679 11299 28685
rect 5592 28648 9628 28676
rect 5592 28636 5598 28648
rect 8570 28608 8576 28620
rect 5368 28580 7052 28608
rect 5368 28552 5396 28580
rect 5169 28543 5227 28549
rect 5169 28509 5181 28543
rect 5215 28509 5227 28543
rect 5350 28540 5356 28552
rect 5311 28512 5356 28540
rect 5169 28503 5227 28509
rect 5350 28500 5356 28512
rect 5408 28500 5414 28552
rect 5537 28543 5595 28549
rect 5537 28509 5549 28543
rect 5583 28540 5595 28543
rect 6914 28540 6920 28552
rect 5583 28512 6920 28540
rect 5583 28509 5595 28512
rect 5537 28503 5595 28509
rect 6914 28500 6920 28512
rect 6972 28500 6978 28552
rect 7024 28540 7052 28580
rect 8312 28580 8576 28608
rect 8312 28552 8340 28580
rect 8570 28568 8576 28580
rect 8628 28568 8634 28620
rect 8294 28540 8300 28552
rect 7024 28512 7144 28540
rect 8207 28512 8300 28540
rect 5442 28432 5448 28484
rect 5500 28472 5506 28484
rect 5500 28444 5545 28472
rect 5500 28432 5506 28444
rect 6454 28432 6460 28484
rect 6512 28472 6518 28484
rect 6641 28475 6699 28481
rect 6641 28472 6653 28475
rect 6512 28444 6653 28472
rect 6512 28432 6518 28444
rect 6641 28441 6653 28444
rect 6687 28441 6699 28475
rect 6641 28435 6699 28441
rect 6730 28432 6736 28484
rect 6788 28472 6794 28484
rect 6825 28475 6883 28481
rect 6825 28472 6837 28475
rect 6788 28444 6837 28472
rect 6788 28432 6794 28444
rect 6825 28441 6837 28444
rect 6871 28441 6883 28475
rect 7006 28472 7012 28484
rect 6967 28444 7012 28472
rect 6825 28435 6883 28441
rect 7006 28432 7012 28444
rect 7064 28432 7070 28484
rect 5718 28404 5724 28416
rect 5679 28376 5724 28404
rect 5718 28364 5724 28376
rect 5776 28364 5782 28416
rect 7116 28404 7144 28512
rect 8294 28500 8300 28512
rect 8352 28500 8358 28552
rect 8389 28543 8447 28549
rect 8389 28509 8401 28543
rect 8435 28509 8447 28543
rect 9122 28540 9128 28552
rect 9083 28512 9128 28540
rect 8389 28503 8447 28509
rect 8110 28432 8116 28484
rect 8168 28472 8174 28484
rect 8404 28472 8432 28503
rect 9122 28500 9128 28512
rect 9180 28500 9186 28552
rect 9600 28549 9628 28648
rect 11241 28645 11253 28679
rect 11287 28676 11299 28679
rect 13538 28676 13544 28688
rect 11287 28648 13544 28676
rect 11287 28645 11299 28648
rect 11241 28639 11299 28645
rect 13538 28636 13544 28648
rect 13596 28676 13602 28688
rect 15194 28676 15200 28688
rect 13596 28648 15200 28676
rect 13596 28636 13602 28648
rect 15194 28636 15200 28648
rect 15252 28636 15258 28688
rect 16408 28685 16436 28716
rect 16850 28704 16856 28716
rect 16908 28704 16914 28756
rect 17310 28704 17316 28756
rect 17368 28744 17374 28756
rect 17865 28747 17923 28753
rect 17865 28744 17877 28747
rect 17368 28716 17877 28744
rect 17368 28704 17374 28716
rect 17865 28713 17877 28716
rect 17911 28713 17923 28747
rect 17865 28707 17923 28713
rect 18506 28704 18512 28756
rect 18564 28744 18570 28756
rect 18564 28716 21404 28744
rect 18564 28704 18570 28716
rect 16393 28679 16451 28685
rect 16393 28645 16405 28679
rect 16439 28645 16451 28679
rect 16758 28676 16764 28688
rect 16393 28639 16451 28645
rect 16500 28648 16764 28676
rect 11146 28568 11152 28620
rect 11204 28608 11210 28620
rect 13354 28608 13360 28620
rect 11204 28580 12434 28608
rect 11204 28568 11210 28580
rect 9585 28543 9643 28549
rect 9585 28509 9597 28543
rect 9631 28509 9643 28543
rect 12406 28540 12434 28580
rect 12912 28580 13360 28608
rect 12912 28549 12940 28580
rect 13354 28568 13360 28580
rect 13412 28608 13418 28620
rect 14366 28608 14372 28620
rect 13412 28580 14372 28608
rect 13412 28568 13418 28580
rect 14366 28568 14372 28580
rect 14424 28568 14430 28620
rect 16500 28617 16528 28648
rect 16758 28636 16764 28648
rect 16816 28636 16822 28688
rect 16868 28676 16896 28704
rect 17678 28676 17684 28688
rect 16868 28648 17684 28676
rect 17678 28636 17684 28648
rect 17736 28636 17742 28688
rect 19334 28676 19340 28688
rect 17788 28648 19340 28676
rect 16485 28611 16543 28617
rect 16485 28577 16497 28611
rect 16531 28577 16543 28611
rect 16485 28571 16543 28577
rect 12713 28543 12771 28549
rect 12713 28540 12725 28543
rect 9585 28503 9643 28509
rect 9688 28512 11744 28540
rect 12406 28512 12725 28540
rect 8168 28444 8432 28472
rect 8168 28432 8174 28444
rect 8478 28432 8484 28484
rect 8536 28472 8542 28484
rect 9688 28472 9716 28512
rect 8536 28444 9716 28472
rect 8536 28432 8542 28444
rect 10410 28432 10416 28484
rect 10468 28472 10474 28484
rect 10873 28475 10931 28481
rect 10873 28472 10885 28475
rect 10468 28444 10885 28472
rect 10468 28432 10474 28444
rect 10873 28441 10885 28444
rect 10919 28472 10931 28475
rect 10962 28472 10968 28484
rect 10919 28444 10968 28472
rect 10919 28441 10931 28444
rect 10873 28435 10931 28441
rect 10962 28432 10968 28444
rect 11020 28432 11026 28484
rect 8018 28404 8024 28416
rect 7116 28376 8024 28404
rect 8018 28364 8024 28376
rect 8076 28404 8082 28416
rect 8297 28407 8355 28413
rect 8297 28404 8309 28407
rect 8076 28376 8309 28404
rect 8076 28364 8082 28376
rect 8297 28373 8309 28376
rect 8343 28373 8355 28407
rect 8297 28367 8355 28373
rect 9122 28364 9128 28416
rect 9180 28404 9186 28416
rect 9217 28407 9275 28413
rect 9217 28404 9229 28407
rect 9180 28376 9229 28404
rect 9180 28364 9186 28376
rect 9217 28373 9229 28376
rect 9263 28404 9275 28407
rect 11057 28407 11115 28413
rect 11057 28404 11069 28407
rect 9263 28376 11069 28404
rect 9263 28373 9275 28376
rect 9217 28367 9275 28373
rect 11057 28373 11069 28376
rect 11103 28404 11115 28407
rect 11606 28404 11612 28416
rect 11103 28376 11612 28404
rect 11103 28373 11115 28376
rect 11057 28367 11115 28373
rect 11606 28364 11612 28376
rect 11664 28364 11670 28416
rect 11716 28404 11744 28512
rect 12713 28509 12725 28512
rect 12759 28509 12771 28543
rect 12713 28503 12771 28509
rect 12897 28543 12955 28549
rect 12897 28509 12909 28543
rect 12943 28509 12955 28543
rect 14274 28540 14280 28552
rect 14235 28512 14280 28540
rect 12897 28503 12955 28509
rect 14274 28500 14280 28512
rect 14332 28500 14338 28552
rect 14458 28540 14464 28552
rect 14419 28512 14464 28540
rect 14458 28500 14464 28512
rect 14516 28500 14522 28552
rect 14642 28540 14648 28552
rect 14603 28512 14648 28540
rect 14642 28500 14648 28512
rect 14700 28500 14706 28552
rect 16298 28540 16304 28552
rect 16259 28512 16304 28540
rect 16298 28500 16304 28512
rect 16356 28500 16362 28552
rect 16577 28543 16635 28549
rect 16577 28509 16589 28543
rect 16623 28509 16635 28543
rect 16758 28540 16764 28552
rect 16719 28512 16764 28540
rect 16577 28503 16635 28509
rect 11790 28432 11796 28484
rect 11848 28472 11854 28484
rect 11977 28475 12035 28481
rect 11848 28444 11893 28472
rect 11848 28432 11854 28444
rect 11977 28441 11989 28475
rect 12023 28472 12035 28475
rect 14553 28475 14611 28481
rect 12023 28444 12296 28472
rect 12023 28441 12035 28444
rect 11977 28435 12035 28441
rect 12161 28407 12219 28413
rect 12161 28404 12173 28407
rect 11716 28376 12173 28404
rect 12161 28373 12173 28376
rect 12207 28373 12219 28407
rect 12268 28404 12296 28444
rect 14553 28441 14565 28475
rect 14599 28472 14611 28475
rect 16206 28472 16212 28484
rect 14599 28444 16212 28472
rect 14599 28441 14611 28444
rect 14553 28435 14611 28441
rect 16206 28432 16212 28444
rect 16264 28432 16270 28484
rect 16592 28472 16620 28503
rect 16758 28500 16764 28512
rect 16816 28500 16822 28552
rect 17788 28549 17816 28648
rect 19334 28636 19340 28648
rect 19392 28636 19398 28688
rect 20438 28676 20444 28688
rect 19444 28648 20444 28676
rect 19444 28552 19472 28648
rect 20438 28636 20444 28648
rect 20496 28636 20502 28688
rect 20622 28608 20628 28620
rect 19812 28580 20628 28608
rect 17773 28543 17831 28549
rect 17773 28509 17785 28543
rect 17819 28509 17831 28543
rect 17773 28503 17831 28509
rect 17862 28500 17868 28552
rect 17920 28540 17926 28552
rect 17957 28543 18015 28549
rect 17957 28540 17969 28543
rect 17920 28512 17969 28540
rect 17920 28500 17926 28512
rect 17957 28509 17969 28512
rect 18003 28509 18015 28543
rect 17957 28503 18015 28509
rect 17034 28472 17040 28484
rect 16592 28444 17040 28472
rect 17034 28432 17040 28444
rect 17092 28432 17098 28484
rect 17972 28472 18000 28503
rect 18874 28500 18880 28552
rect 18932 28540 18938 28552
rect 19426 28540 19432 28552
rect 18932 28512 19432 28540
rect 18932 28500 18938 28512
rect 19426 28500 19432 28512
rect 19484 28500 19490 28552
rect 19610 28500 19616 28552
rect 19668 28540 19674 28552
rect 19812 28549 19840 28580
rect 20622 28568 20628 28580
rect 20680 28608 20686 28620
rect 21269 28611 21327 28617
rect 21269 28608 21281 28611
rect 20680 28580 21281 28608
rect 20680 28568 20686 28580
rect 21269 28577 21281 28580
rect 21315 28577 21327 28611
rect 21376 28608 21404 28716
rect 21542 28704 21548 28756
rect 21600 28744 21606 28756
rect 23293 28747 23351 28753
rect 23293 28744 23305 28747
rect 21600 28716 23305 28744
rect 21600 28704 21606 28716
rect 23293 28713 23305 28716
rect 23339 28744 23351 28747
rect 23474 28744 23480 28756
rect 23339 28716 23480 28744
rect 23339 28713 23351 28716
rect 23293 28707 23351 28713
rect 23474 28704 23480 28716
rect 23532 28704 23538 28756
rect 24854 28704 24860 28756
rect 24912 28744 24918 28756
rect 24949 28747 25007 28753
rect 24949 28744 24961 28747
rect 24912 28716 24961 28744
rect 24912 28704 24918 28716
rect 24949 28713 24961 28716
rect 24995 28744 25007 28747
rect 25958 28744 25964 28756
rect 24995 28716 25964 28744
rect 24995 28713 25007 28716
rect 24949 28707 25007 28713
rect 25958 28704 25964 28716
rect 26016 28704 26022 28756
rect 27246 28704 27252 28756
rect 27304 28744 27310 28756
rect 27982 28744 27988 28756
rect 27304 28716 27988 28744
rect 27304 28704 27310 28716
rect 27982 28704 27988 28716
rect 28040 28704 28046 28756
rect 30190 28744 30196 28756
rect 30103 28716 30196 28744
rect 30190 28704 30196 28716
rect 30248 28744 30254 28756
rect 32582 28744 32588 28756
rect 30248 28716 32588 28744
rect 30248 28704 30254 28716
rect 32582 28704 32588 28716
rect 32640 28704 32646 28756
rect 35342 28704 35348 28756
rect 35400 28744 35406 28756
rect 35710 28744 35716 28756
rect 35400 28716 35716 28744
rect 35400 28704 35406 28716
rect 35710 28704 35716 28716
rect 35768 28704 35774 28756
rect 23385 28679 23443 28685
rect 23385 28645 23397 28679
rect 23431 28676 23443 28679
rect 25041 28679 25099 28685
rect 23431 28648 24992 28676
rect 23431 28645 23443 28648
rect 23385 28639 23443 28645
rect 24964 28608 24992 28648
rect 25041 28645 25053 28679
rect 25087 28676 25099 28679
rect 26234 28676 26240 28688
rect 25087 28648 26240 28676
rect 25087 28645 25099 28648
rect 25041 28639 25099 28645
rect 26234 28636 26240 28648
rect 26292 28636 26298 28688
rect 28442 28636 28448 28688
rect 28500 28676 28506 28688
rect 28902 28676 28908 28688
rect 28500 28648 28908 28676
rect 28500 28636 28506 28648
rect 28902 28636 28908 28648
rect 28960 28636 28966 28688
rect 25133 28611 25191 28617
rect 25133 28608 25145 28611
rect 21376 28580 23612 28608
rect 24964 28580 25145 28608
rect 21269 28571 21327 28577
rect 19705 28543 19763 28549
rect 19705 28540 19717 28543
rect 19668 28512 19717 28540
rect 19668 28500 19674 28512
rect 19705 28509 19717 28512
rect 19751 28509 19763 28543
rect 19705 28503 19763 28509
rect 19797 28543 19855 28549
rect 19797 28509 19809 28543
rect 19843 28509 19855 28543
rect 19797 28503 19855 28509
rect 19889 28543 19947 28549
rect 19889 28509 19901 28543
rect 19935 28509 19947 28543
rect 19889 28503 19947 28509
rect 20073 28543 20131 28549
rect 20073 28509 20085 28543
rect 20119 28540 20131 28543
rect 20530 28540 20536 28552
rect 20119 28512 20536 28540
rect 20119 28509 20131 28512
rect 20073 28503 20131 28509
rect 19904 28472 19932 28503
rect 20530 28500 20536 28512
rect 20588 28500 20594 28552
rect 20993 28543 21051 28549
rect 20993 28509 21005 28543
rect 21039 28540 21051 28543
rect 21358 28540 21364 28552
rect 21039 28512 21364 28540
rect 21039 28509 21051 28512
rect 20993 28503 21051 28509
rect 21358 28500 21364 28512
rect 21416 28500 21422 28552
rect 21634 28500 21640 28552
rect 21692 28540 21698 28552
rect 21818 28540 21824 28552
rect 21692 28512 21824 28540
rect 21692 28500 21698 28512
rect 21818 28500 21824 28512
rect 21876 28540 21882 28552
rect 23584 28549 23612 28580
rect 25133 28577 25145 28580
rect 25179 28608 25191 28611
rect 25866 28608 25872 28620
rect 25179 28580 25872 28608
rect 25179 28577 25191 28580
rect 25133 28571 25191 28577
rect 25866 28568 25872 28580
rect 25924 28568 25930 28620
rect 30006 28608 30012 28620
rect 28000 28580 30012 28608
rect 23109 28543 23167 28549
rect 23109 28540 23121 28543
rect 21876 28512 23121 28540
rect 21876 28500 21882 28512
rect 23109 28509 23121 28512
rect 23155 28509 23167 28543
rect 23109 28503 23167 28509
rect 23201 28543 23259 28549
rect 23201 28509 23213 28543
rect 23247 28509 23259 28543
rect 23201 28503 23259 28509
rect 23569 28543 23627 28549
rect 23569 28509 23581 28543
rect 23615 28540 23627 28543
rect 24581 28543 24639 28549
rect 24581 28540 24593 28543
rect 23615 28512 24593 28540
rect 23615 28509 23627 28512
rect 23569 28503 23627 28509
rect 24581 28509 24593 28512
rect 24627 28509 24639 28543
rect 24581 28503 24639 28509
rect 17972 28444 19932 28472
rect 12710 28404 12716 28416
rect 12268 28376 12716 28404
rect 12161 28367 12219 28373
rect 12710 28364 12716 28376
rect 12768 28364 12774 28416
rect 12805 28407 12863 28413
rect 12805 28373 12817 28407
rect 12851 28404 12863 28407
rect 13262 28404 13268 28416
rect 12851 28376 13268 28404
rect 12851 28373 12863 28376
rect 12805 28367 12863 28373
rect 13262 28364 13268 28376
rect 13320 28364 13326 28416
rect 15010 28364 15016 28416
rect 15068 28404 15074 28416
rect 19429 28407 19487 28413
rect 19429 28404 19441 28407
rect 15068 28376 19441 28404
rect 15068 28364 15074 28376
rect 19429 28373 19441 28376
rect 19475 28373 19487 28407
rect 20548 28404 20576 28500
rect 21478 28475 21536 28481
rect 21478 28441 21490 28475
rect 21524 28472 21536 28475
rect 22646 28472 22652 28484
rect 21524 28444 22652 28472
rect 21524 28441 21536 28444
rect 21478 28435 21536 28441
rect 22646 28432 22652 28444
rect 22704 28432 22710 28484
rect 21361 28407 21419 28413
rect 21361 28404 21373 28407
rect 20548 28376 21373 28404
rect 19429 28367 19487 28373
rect 21361 28373 21373 28376
rect 21407 28373 21419 28407
rect 21361 28367 21419 28373
rect 21637 28407 21695 28413
rect 21637 28373 21649 28407
rect 21683 28404 21695 28407
rect 22094 28404 22100 28416
rect 21683 28376 22100 28404
rect 21683 28373 21695 28376
rect 21637 28367 21695 28373
rect 22094 28364 22100 28376
rect 22152 28364 22158 28416
rect 22833 28407 22891 28413
rect 22833 28373 22845 28407
rect 22879 28404 22891 28407
rect 22922 28404 22928 28416
rect 22879 28376 22928 28404
rect 22879 28373 22891 28376
rect 22833 28367 22891 28373
rect 22922 28364 22928 28376
rect 22980 28364 22986 28416
rect 23216 28404 23244 28503
rect 24670 28500 24676 28552
rect 24728 28540 24734 28552
rect 28000 28549 28028 28580
rect 30006 28568 30012 28580
rect 30064 28568 30070 28620
rect 27249 28543 27307 28549
rect 27249 28540 27261 28543
rect 24728 28512 27261 28540
rect 24728 28500 24734 28512
rect 27249 28509 27261 28512
rect 27295 28509 27307 28543
rect 27249 28503 27307 28509
rect 27985 28543 28043 28549
rect 27985 28509 27997 28543
rect 28031 28509 28043 28543
rect 28350 28540 28356 28552
rect 28311 28512 28356 28540
rect 27985 28503 28043 28509
rect 28350 28500 28356 28512
rect 28408 28540 28414 28552
rect 28810 28540 28816 28552
rect 28408 28512 28816 28540
rect 28408 28500 28414 28512
rect 28810 28500 28816 28512
rect 28868 28500 28874 28552
rect 30208 28549 30236 28704
rect 31662 28636 31668 28688
rect 31720 28676 31726 28688
rect 31941 28679 31999 28685
rect 31720 28648 31800 28676
rect 31720 28636 31726 28648
rect 30466 28608 30472 28620
rect 30427 28580 30472 28608
rect 30466 28568 30472 28580
rect 30524 28568 30530 28620
rect 30193 28543 30251 28549
rect 30193 28509 30205 28543
rect 30239 28509 30251 28543
rect 30193 28503 30251 28509
rect 30374 28500 30380 28552
rect 30432 28540 30438 28552
rect 30558 28540 30564 28552
rect 30432 28512 30564 28540
rect 30432 28500 30438 28512
rect 30558 28500 30564 28512
rect 30616 28500 30622 28552
rect 31294 28540 31300 28552
rect 31255 28512 31300 28540
rect 31294 28500 31300 28512
rect 31352 28500 31358 28552
rect 31386 28500 31392 28552
rect 31444 28540 31450 28552
rect 31444 28512 31489 28540
rect 31444 28500 31450 28512
rect 31570 28500 31576 28552
rect 31628 28540 31634 28552
rect 31772 28549 31800 28648
rect 31941 28645 31953 28679
rect 31987 28676 31999 28679
rect 32490 28676 32496 28688
rect 31987 28648 32496 28676
rect 31987 28645 31999 28648
rect 31941 28639 31999 28645
rect 32490 28636 32496 28648
rect 32548 28676 32554 28688
rect 32548 28648 32720 28676
rect 32548 28636 32554 28648
rect 32692 28617 32720 28648
rect 32677 28611 32735 28617
rect 32677 28577 32689 28611
rect 32723 28577 32735 28611
rect 33134 28608 33140 28620
rect 33095 28580 33140 28608
rect 32677 28571 32735 28577
rect 33134 28568 33140 28580
rect 33192 28568 33198 28620
rect 35713 28611 35771 28617
rect 35713 28577 35725 28611
rect 35759 28608 35771 28611
rect 36814 28608 36820 28620
rect 35759 28580 36820 28608
rect 35759 28577 35771 28580
rect 35713 28571 35771 28577
rect 36814 28568 36820 28580
rect 36872 28568 36878 28620
rect 31762 28543 31820 28549
rect 31628 28512 31673 28540
rect 31628 28500 31634 28512
rect 31762 28509 31774 28543
rect 31808 28509 31820 28543
rect 32766 28540 32772 28552
rect 32727 28512 32772 28540
rect 31762 28503 31820 28509
rect 32766 28500 32772 28512
rect 32824 28500 32830 28552
rect 24118 28432 24124 28484
rect 24176 28472 24182 28484
rect 28169 28475 28227 28481
rect 28169 28472 28181 28475
rect 24176 28444 28181 28472
rect 24176 28432 24182 28444
rect 28169 28441 28181 28444
rect 28215 28441 28227 28475
rect 28169 28435 28227 28441
rect 28258 28432 28264 28484
rect 28316 28472 28322 28484
rect 30926 28472 30932 28484
rect 28316 28444 30932 28472
rect 28316 28432 28322 28444
rect 30926 28432 30932 28444
rect 30984 28432 30990 28484
rect 31665 28475 31723 28481
rect 31665 28441 31677 28475
rect 31711 28472 31723 28475
rect 32214 28472 32220 28484
rect 31711 28444 32220 28472
rect 31711 28441 31723 28444
rect 31665 28435 31723 28441
rect 32214 28432 32220 28444
rect 32272 28432 32278 28484
rect 34885 28475 34943 28481
rect 34885 28441 34897 28475
rect 34931 28472 34943 28475
rect 35342 28472 35348 28484
rect 34931 28444 35348 28472
rect 34931 28441 34943 28444
rect 34885 28435 34943 28441
rect 35342 28432 35348 28444
rect 35400 28432 35406 28484
rect 37084 28475 37142 28481
rect 37084 28441 37096 28475
rect 37130 28472 37142 28475
rect 37458 28472 37464 28484
rect 37130 28444 37464 28472
rect 37130 28441 37142 28444
rect 37084 28435 37142 28441
rect 37458 28432 37464 28444
rect 37516 28432 37522 28484
rect 23290 28404 23296 28416
rect 23216 28376 23296 28404
rect 23290 28364 23296 28376
rect 23348 28364 23354 28416
rect 24946 28364 24952 28416
rect 25004 28404 25010 28416
rect 25409 28407 25467 28413
rect 25409 28404 25421 28407
rect 25004 28376 25421 28404
rect 25004 28364 25010 28376
rect 25409 28373 25421 28376
rect 25455 28373 25467 28407
rect 25409 28367 25467 28373
rect 27246 28364 27252 28416
rect 27304 28404 27310 28416
rect 27433 28407 27491 28413
rect 27433 28404 27445 28407
rect 27304 28376 27445 28404
rect 27304 28364 27310 28376
rect 27433 28373 27445 28376
rect 27479 28373 27491 28407
rect 27433 28367 27491 28373
rect 27614 28364 27620 28416
rect 27672 28404 27678 28416
rect 28537 28407 28595 28413
rect 28537 28404 28549 28407
rect 27672 28376 28549 28404
rect 27672 28364 27678 28376
rect 28537 28373 28549 28376
rect 28583 28373 28595 28407
rect 28537 28367 28595 28373
rect 30006 28364 30012 28416
rect 30064 28404 30070 28416
rect 35802 28404 35808 28416
rect 30064 28376 35808 28404
rect 30064 28364 30070 28376
rect 35802 28364 35808 28376
rect 35860 28364 35866 28416
rect 38194 28404 38200 28416
rect 38155 28376 38200 28404
rect 38194 28364 38200 28376
rect 38252 28364 38258 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 5184 28172 7052 28200
rect 4798 28024 4804 28076
rect 4856 28064 4862 28076
rect 5184 28073 5212 28172
rect 4893 28067 4951 28073
rect 4893 28064 4905 28067
rect 4856 28036 4905 28064
rect 4856 28024 4862 28036
rect 4893 28033 4905 28036
rect 4939 28033 4951 28067
rect 4893 28027 4951 28033
rect 5169 28067 5227 28073
rect 5169 28033 5181 28067
rect 5215 28033 5227 28067
rect 7024 28064 7052 28172
rect 7098 28160 7104 28212
rect 7156 28200 7162 28212
rect 8478 28200 8484 28212
rect 7156 28172 8484 28200
rect 7156 28160 7162 28172
rect 8478 28160 8484 28172
rect 8536 28200 8542 28212
rect 11054 28200 11060 28212
rect 8536 28172 9076 28200
rect 11015 28172 11060 28200
rect 8536 28160 8542 28172
rect 7285 28135 7343 28141
rect 7285 28101 7297 28135
rect 7331 28132 7343 28135
rect 7374 28132 7380 28144
rect 7331 28104 7380 28132
rect 7331 28101 7343 28104
rect 7285 28095 7343 28101
rect 7374 28092 7380 28104
rect 7432 28092 7438 28144
rect 9048 28132 9076 28172
rect 11054 28160 11060 28172
rect 11112 28160 11118 28212
rect 11790 28160 11796 28212
rect 11848 28200 11854 28212
rect 16942 28200 16948 28212
rect 11848 28172 14587 28200
rect 16903 28172 16948 28200
rect 11848 28160 11854 28172
rect 9048 28104 9168 28132
rect 7558 28064 7564 28076
rect 7024 28036 7564 28064
rect 5169 28027 5227 28033
rect 7558 28024 7564 28036
rect 7616 28024 7622 28076
rect 8294 28064 8300 28076
rect 8255 28036 8300 28064
rect 8294 28024 8300 28036
rect 8352 28024 8358 28076
rect 8573 28067 8631 28073
rect 8573 28033 8585 28067
rect 8619 28064 8631 28067
rect 9030 28064 9036 28076
rect 8619 28036 9036 28064
rect 8619 28033 8631 28036
rect 8573 28027 8631 28033
rect 9030 28024 9036 28036
rect 9088 28024 9094 28076
rect 9140 28073 9168 28104
rect 9306 28092 9312 28144
rect 9364 28132 9370 28144
rect 9582 28132 9588 28144
rect 9364 28104 9588 28132
rect 9364 28092 9370 28104
rect 9582 28092 9588 28104
rect 9640 28132 9646 28144
rect 9640 28104 11192 28132
rect 9640 28092 9646 28104
rect 9125 28067 9183 28073
rect 9125 28033 9137 28067
rect 9171 28033 9183 28067
rect 9398 28064 9404 28076
rect 9359 28036 9404 28064
rect 9125 28027 9183 28033
rect 9398 28024 9404 28036
rect 9456 28024 9462 28076
rect 9953 28067 10011 28073
rect 9953 28033 9965 28067
rect 9999 28033 10011 28067
rect 10226 28064 10232 28076
rect 10187 28036 10232 28064
rect 9953 28027 10011 28033
rect 5077 27999 5135 28005
rect 5077 27965 5089 27999
rect 5123 27996 5135 27999
rect 5258 27996 5264 28008
rect 5123 27968 5264 27996
rect 5123 27965 5135 27968
rect 5077 27959 5135 27965
rect 5258 27956 5264 27968
rect 5316 27956 5322 28008
rect 6362 27956 6368 28008
rect 6420 27996 6426 28008
rect 6917 27999 6975 28005
rect 6917 27996 6929 27999
rect 6420 27968 6929 27996
rect 6420 27956 6426 27968
rect 6917 27965 6929 27968
rect 6963 27996 6975 27999
rect 7834 27996 7840 28008
rect 6963 27968 7840 27996
rect 6963 27965 6975 27968
rect 6917 27959 6975 27965
rect 7834 27956 7840 27968
rect 7892 27956 7898 28008
rect 9858 27996 9864 28008
rect 9232 27968 9864 27996
rect 7098 27888 7104 27940
rect 7156 27928 7162 27940
rect 7469 27931 7527 27937
rect 7469 27928 7481 27931
rect 7156 27900 7481 27928
rect 7156 27888 7162 27900
rect 7469 27897 7481 27900
rect 7515 27897 7527 27931
rect 7469 27891 7527 27897
rect 7558 27888 7564 27940
rect 7616 27928 7622 27940
rect 8389 27931 8447 27937
rect 8389 27928 8401 27931
rect 7616 27900 8401 27928
rect 7616 27888 7622 27900
rect 8389 27897 8401 27900
rect 8435 27897 8447 27931
rect 8389 27891 8447 27897
rect 4982 27860 4988 27872
rect 4943 27832 4988 27860
rect 4982 27820 4988 27832
rect 5040 27820 5046 27872
rect 5074 27820 5080 27872
rect 5132 27860 5138 27872
rect 5353 27863 5411 27869
rect 5353 27860 5365 27863
rect 5132 27832 5365 27860
rect 5132 27820 5138 27832
rect 5353 27829 5365 27832
rect 5399 27829 5411 27863
rect 5353 27823 5411 27829
rect 6730 27820 6736 27872
rect 6788 27860 6794 27872
rect 7285 27863 7343 27869
rect 7285 27860 7297 27863
rect 6788 27832 7297 27860
rect 6788 27820 6794 27832
rect 7285 27829 7297 27832
rect 7331 27829 7343 27863
rect 7285 27823 7343 27829
rect 8294 27820 8300 27872
rect 8352 27860 8358 27872
rect 9232 27869 9260 27968
rect 9858 27956 9864 27968
rect 9916 27996 9922 28008
rect 9968 27996 9996 28027
rect 10226 28024 10232 28036
rect 10284 28024 10290 28076
rect 11164 28073 11192 28104
rect 10965 28067 11023 28073
rect 10965 28033 10977 28067
rect 11011 28033 11023 28067
rect 10965 28027 11023 28033
rect 11149 28067 11207 28073
rect 11149 28033 11161 28067
rect 11195 28033 11207 28067
rect 12710 28064 12716 28076
rect 12671 28036 12716 28064
rect 11149 28027 11207 28033
rect 10134 27996 10140 28008
rect 9916 27968 9996 27996
rect 10095 27968 10140 27996
rect 9916 27956 9922 27968
rect 10134 27956 10140 27968
rect 10192 27956 10198 28008
rect 10980 27996 11008 28027
rect 12710 28024 12716 28036
rect 12768 28024 12774 28076
rect 13188 28073 13216 28172
rect 13262 28092 13268 28144
rect 13320 28132 13326 28144
rect 14185 28135 14243 28141
rect 14185 28132 14197 28135
rect 13320 28104 14197 28132
rect 13320 28092 13326 28104
rect 14185 28101 14197 28104
rect 14231 28101 14243 28135
rect 14185 28095 14243 28101
rect 13173 28067 13231 28073
rect 13173 28033 13185 28067
rect 13219 28033 13231 28067
rect 13173 28027 13231 28033
rect 13449 28067 13507 28073
rect 13449 28033 13461 28067
rect 13495 28064 13507 28067
rect 13722 28064 13728 28076
rect 13495 28036 13728 28064
rect 13495 28033 13507 28036
rect 13449 28027 13507 28033
rect 13722 28024 13728 28036
rect 13780 28064 13786 28076
rect 14001 28067 14059 28073
rect 14001 28064 14013 28067
rect 13780 28036 14013 28064
rect 13780 28024 13786 28036
rect 14001 28033 14013 28036
rect 14047 28033 14059 28067
rect 14001 28027 14059 28033
rect 14277 28067 14335 28073
rect 14277 28033 14289 28067
rect 14323 28033 14335 28067
rect 14277 28027 14335 28033
rect 12066 27996 12072 28008
rect 10980 27968 12072 27996
rect 12066 27956 12072 27968
rect 12124 27956 12130 28008
rect 10413 27931 10471 27937
rect 10413 27897 10425 27931
rect 10459 27928 10471 27931
rect 11422 27928 11428 27940
rect 10459 27900 11428 27928
rect 10459 27897 10471 27900
rect 10413 27891 10471 27897
rect 11422 27888 11428 27900
rect 11480 27888 11486 27940
rect 14292 27928 14320 28027
rect 14366 28024 14372 28076
rect 14424 28064 14430 28076
rect 14424 28036 14469 28064
rect 14424 28024 14430 28036
rect 14559 27996 14587 28172
rect 16942 28160 16948 28172
rect 17000 28160 17006 28212
rect 17586 28160 17592 28212
rect 17644 28200 17650 28212
rect 24121 28203 24179 28209
rect 24121 28200 24133 28203
rect 17644 28172 24133 28200
rect 17644 28160 17650 28172
rect 24121 28169 24133 28172
rect 24167 28169 24179 28203
rect 25593 28203 25651 28209
rect 25593 28200 25605 28203
rect 24121 28163 24179 28169
rect 24412 28172 25605 28200
rect 16758 28092 16764 28144
rect 16816 28132 16822 28144
rect 18782 28132 18788 28144
rect 16816 28104 18788 28132
rect 16816 28092 16822 28104
rect 16868 28073 16896 28104
rect 18782 28092 18788 28104
rect 18840 28092 18846 28144
rect 20438 28092 20444 28144
rect 20496 28132 20502 28144
rect 21542 28132 21548 28144
rect 20496 28104 21548 28132
rect 20496 28092 20502 28104
rect 21542 28092 21548 28104
rect 21600 28092 21606 28144
rect 22554 28132 22560 28144
rect 22515 28104 22560 28132
rect 22554 28092 22560 28104
rect 22612 28092 22618 28144
rect 23661 28135 23719 28141
rect 23661 28101 23673 28135
rect 23707 28132 23719 28135
rect 24302 28132 24308 28144
rect 23707 28104 24308 28132
rect 23707 28101 23719 28104
rect 23661 28095 23719 28101
rect 24302 28092 24308 28104
rect 24360 28092 24366 28144
rect 16853 28067 16911 28073
rect 16853 28033 16865 28067
rect 16899 28033 16911 28067
rect 16853 28027 16911 28033
rect 17034 28024 17040 28076
rect 17092 28064 17098 28076
rect 18598 28064 18604 28076
rect 17092 28036 18604 28064
rect 17092 28024 17098 28036
rect 18598 28024 18604 28036
rect 18656 28024 18662 28076
rect 18874 28064 18880 28076
rect 18835 28036 18880 28064
rect 18874 28024 18880 28036
rect 18932 28024 18938 28076
rect 18966 28024 18972 28076
rect 19024 28064 19030 28076
rect 19061 28067 19119 28073
rect 19061 28064 19073 28067
rect 19024 28036 19073 28064
rect 19024 28024 19030 28036
rect 19061 28033 19073 28036
rect 19107 28033 19119 28067
rect 19061 28027 19119 28033
rect 19978 28024 19984 28076
rect 20036 28064 20042 28076
rect 20073 28067 20131 28073
rect 20073 28064 20085 28067
rect 20036 28036 20085 28064
rect 20036 28024 20042 28036
rect 20073 28033 20085 28036
rect 20119 28033 20131 28067
rect 20073 28027 20131 28033
rect 22094 28024 22100 28076
rect 22152 28064 22158 28076
rect 22152 28036 22197 28064
rect 22152 28024 22158 28036
rect 23106 28024 23112 28076
rect 23164 28064 23170 28076
rect 24412 28064 24440 28172
rect 25593 28169 25605 28172
rect 25639 28200 25651 28203
rect 25774 28200 25780 28212
rect 25639 28172 25780 28200
rect 25639 28169 25651 28172
rect 25593 28163 25651 28169
rect 25774 28160 25780 28172
rect 25832 28160 25838 28212
rect 26510 28160 26516 28212
rect 26568 28200 26574 28212
rect 28902 28200 28908 28212
rect 26568 28172 28908 28200
rect 26568 28160 26574 28172
rect 24854 28092 24860 28144
rect 24912 28132 24918 28144
rect 25222 28132 25228 28144
rect 24912 28104 25228 28132
rect 24912 28092 24918 28104
rect 25222 28092 25228 28104
rect 25280 28132 25286 28144
rect 27154 28132 27160 28144
rect 25280 28104 25728 28132
rect 27115 28104 27160 28132
rect 25280 28092 25286 28104
rect 23164 28036 24440 28064
rect 24581 28067 24639 28073
rect 23164 28024 23170 28036
rect 24581 28033 24593 28067
rect 24627 28064 24639 28067
rect 24670 28064 24676 28076
rect 24627 28036 24676 28064
rect 24627 28033 24639 28036
rect 24581 28027 24639 28033
rect 24670 28024 24676 28036
rect 24728 28024 24734 28076
rect 25498 28064 25504 28076
rect 25459 28036 25504 28064
rect 25498 28024 25504 28036
rect 25556 28024 25562 28076
rect 25700 28073 25728 28104
rect 27154 28092 27160 28104
rect 27212 28092 27218 28144
rect 27982 28092 27988 28144
rect 28040 28132 28046 28144
rect 28442 28132 28448 28144
rect 28040 28104 28448 28132
rect 28040 28092 28046 28104
rect 28442 28092 28448 28104
rect 28500 28092 28506 28144
rect 28552 28141 28580 28172
rect 28902 28160 28908 28172
rect 28960 28160 28966 28212
rect 30098 28160 30104 28212
rect 30156 28160 30162 28212
rect 30745 28203 30803 28209
rect 30745 28169 30757 28203
rect 30791 28200 30803 28203
rect 31110 28200 31116 28212
rect 30791 28172 31116 28200
rect 30791 28169 30803 28172
rect 30745 28163 30803 28169
rect 31110 28160 31116 28172
rect 31168 28160 31174 28212
rect 36262 28200 36268 28212
rect 36223 28172 36268 28200
rect 36262 28160 36268 28172
rect 36320 28160 36326 28212
rect 37458 28200 37464 28212
rect 37419 28172 37464 28200
rect 37458 28160 37464 28172
rect 37516 28160 37522 28212
rect 37918 28200 37924 28212
rect 37879 28172 37924 28200
rect 37918 28160 37924 28172
rect 37976 28160 37982 28212
rect 28537 28135 28595 28141
rect 28537 28101 28549 28135
rect 28583 28101 28595 28135
rect 29914 28132 29920 28144
rect 28537 28095 28595 28101
rect 28966 28104 29920 28132
rect 25685 28067 25743 28073
rect 25685 28033 25697 28067
rect 25731 28033 25743 28067
rect 25685 28027 25743 28033
rect 26694 28024 26700 28076
rect 26752 28064 26758 28076
rect 27617 28067 27675 28073
rect 27617 28064 27629 28067
rect 26752 28036 27629 28064
rect 26752 28024 26758 28036
rect 27617 28033 27629 28036
rect 27663 28033 27675 28067
rect 27617 28027 27675 28033
rect 28261 28067 28319 28073
rect 28261 28033 28273 28067
rect 28307 28064 28319 28067
rect 28681 28067 28739 28073
rect 28307 28036 28396 28064
rect 28307 28033 28319 28036
rect 28261 28027 28319 28033
rect 20162 27996 20168 28008
rect 14559 27968 19288 27996
rect 20123 27968 20168 27996
rect 15654 27928 15660 27940
rect 14292 27900 15660 27928
rect 15654 27888 15660 27900
rect 15712 27888 15718 27940
rect 18414 27888 18420 27940
rect 18472 27928 18478 27940
rect 19153 27931 19211 27937
rect 19153 27928 19165 27931
rect 18472 27900 19165 27928
rect 18472 27888 18478 27900
rect 19153 27897 19165 27900
rect 19199 27897 19211 27931
rect 19260 27928 19288 27968
rect 20162 27956 20168 27968
rect 20220 27956 20226 28008
rect 20714 27956 20720 28008
rect 20772 27996 20778 28008
rect 20990 27996 20996 28008
rect 20772 27968 20996 27996
rect 20772 27956 20778 27968
rect 20990 27956 20996 27968
rect 21048 27956 21054 28008
rect 22278 27956 22284 28008
rect 22336 27996 22342 28008
rect 22465 27999 22523 28005
rect 22465 27996 22477 27999
rect 22336 27968 22477 27996
rect 22336 27956 22342 27968
rect 22465 27965 22477 27968
rect 22511 27965 22523 27999
rect 24765 27999 24823 28005
rect 24765 27996 24777 27999
rect 22465 27959 22523 27965
rect 24044 27968 24777 27996
rect 24044 27940 24072 27968
rect 24765 27965 24777 27968
rect 24811 27965 24823 27999
rect 27433 27999 27491 28005
rect 27433 27996 27445 27999
rect 24765 27959 24823 27965
rect 24872 27968 27445 27996
rect 19260 27900 23980 27928
rect 19153 27891 19211 27897
rect 9217 27863 9275 27869
rect 9217 27860 9229 27863
rect 8352 27832 9229 27860
rect 8352 27820 8358 27832
rect 9217 27829 9229 27832
rect 9263 27829 9275 27863
rect 9217 27823 9275 27829
rect 10229 27863 10287 27869
rect 10229 27829 10241 27863
rect 10275 27860 10287 27863
rect 10318 27860 10324 27872
rect 10275 27832 10324 27860
rect 10275 27829 10287 27832
rect 10229 27823 10287 27829
rect 10318 27820 10324 27832
rect 10376 27820 10382 27872
rect 14550 27860 14556 27872
rect 14511 27832 14556 27860
rect 14550 27820 14556 27832
rect 14608 27820 14614 27872
rect 20070 27860 20076 27872
rect 20031 27832 20076 27860
rect 20070 27820 20076 27832
rect 20128 27820 20134 27872
rect 20441 27863 20499 27869
rect 20441 27829 20453 27863
rect 20487 27860 20499 27863
rect 22002 27860 22008 27872
rect 20487 27832 22008 27860
rect 20487 27829 20499 27832
rect 20441 27823 20499 27829
rect 22002 27820 22008 27832
rect 22060 27820 22066 27872
rect 23952 27860 23980 27900
rect 24026 27888 24032 27940
rect 24084 27928 24090 27940
rect 24084 27900 24129 27928
rect 24084 27888 24090 27900
rect 24670 27888 24676 27940
rect 24728 27928 24734 27940
rect 24872 27928 24900 27968
rect 27433 27965 27445 27968
rect 27479 27965 27491 27999
rect 28368 27996 28396 28036
rect 28681 28033 28693 28067
rect 28727 28064 28739 28067
rect 28810 28064 28816 28076
rect 28727 28036 28816 28064
rect 28727 28033 28739 28036
rect 28681 28027 28739 28033
rect 28810 28024 28816 28036
rect 28868 28024 28874 28076
rect 28966 27996 28994 28104
rect 29914 28092 29920 28104
rect 29972 28092 29978 28144
rect 30116 28132 30144 28160
rect 30377 28135 30435 28141
rect 30377 28132 30389 28135
rect 30116 28104 30389 28132
rect 30377 28101 30389 28104
rect 30423 28101 30435 28135
rect 30377 28095 30435 28101
rect 33134 28092 33140 28144
rect 33192 28132 33198 28144
rect 34118 28135 34176 28141
rect 34118 28132 34130 28135
rect 33192 28104 34130 28132
rect 33192 28092 33198 28104
rect 34118 28101 34130 28104
rect 34164 28101 34176 28135
rect 34118 28095 34176 28101
rect 35802 28092 35808 28144
rect 35860 28132 35866 28144
rect 37829 28135 37887 28141
rect 37829 28132 37841 28135
rect 35860 28104 37841 28132
rect 35860 28092 35866 28104
rect 37829 28101 37841 28104
rect 37875 28132 37887 28135
rect 38194 28132 38200 28144
rect 37875 28104 38200 28132
rect 37875 28101 37887 28104
rect 37829 28095 37887 28101
rect 38194 28092 38200 28104
rect 38252 28092 38258 28144
rect 29638 28024 29644 28076
rect 29696 28064 29702 28076
rect 30006 28064 30012 28076
rect 29696 28036 30012 28064
rect 29696 28024 29702 28036
rect 30006 28024 30012 28036
rect 30064 28064 30070 28076
rect 30101 28067 30159 28073
rect 30101 28064 30113 28067
rect 30064 28036 30113 28064
rect 30064 28024 30070 28036
rect 30101 28033 30113 28036
rect 30147 28033 30159 28067
rect 30101 28027 30159 28033
rect 30190 28024 30196 28076
rect 30248 28064 30254 28076
rect 30469 28067 30527 28073
rect 30469 28064 30481 28067
rect 30248 28036 30293 28064
rect 30392 28036 30481 28064
rect 30248 28024 30254 28036
rect 30392 28008 30420 28036
rect 30469 28033 30481 28036
rect 30515 28033 30527 28067
rect 30469 28027 30527 28033
rect 30558 28024 30564 28076
rect 30616 28073 30622 28076
rect 30616 28064 30624 28073
rect 31202 28064 31208 28076
rect 30616 28036 31208 28064
rect 30616 28027 30624 28036
rect 30616 28024 30622 28027
rect 31202 28024 31208 28036
rect 31260 28024 31266 28076
rect 32674 28024 32680 28076
rect 32732 28064 32738 28076
rect 33042 28064 33048 28076
rect 32732 28036 33048 28064
rect 32732 28024 32738 28036
rect 33042 28024 33048 28036
rect 33100 28064 33106 28076
rect 33873 28067 33931 28073
rect 33873 28064 33885 28067
rect 33100 28036 33885 28064
rect 33100 28024 33106 28036
rect 33873 28033 33885 28036
rect 33919 28033 33931 28067
rect 36078 28064 36084 28076
rect 36039 28036 36084 28064
rect 33873 28027 33931 28033
rect 36078 28024 36084 28036
rect 36136 28024 36142 28076
rect 28368 27968 28994 27996
rect 27433 27959 27491 27965
rect 30374 27956 30380 28008
rect 30432 27956 30438 28008
rect 38010 27996 38016 28008
rect 37971 27968 38016 27996
rect 38010 27956 38016 27968
rect 38068 27956 38074 28008
rect 24728 27900 24900 27928
rect 24728 27888 24734 27900
rect 25958 27888 25964 27940
rect 26016 27928 26022 27940
rect 27338 27928 27344 27940
rect 26016 27900 27344 27928
rect 26016 27888 26022 27900
rect 27338 27888 27344 27900
rect 27396 27888 27402 27940
rect 27522 27888 27528 27940
rect 27580 27928 27586 27940
rect 31386 27928 31392 27940
rect 27580 27900 31392 27928
rect 27580 27888 27586 27900
rect 31386 27888 31392 27900
rect 31444 27928 31450 27940
rect 31444 27900 33272 27928
rect 31444 27888 31450 27900
rect 33244 27872 33272 27900
rect 26142 27860 26148 27872
rect 23952 27832 26148 27860
rect 26142 27820 26148 27832
rect 26200 27820 26206 27872
rect 27430 27860 27436 27872
rect 27391 27832 27436 27860
rect 27430 27820 27436 27832
rect 27488 27820 27494 27872
rect 27798 27860 27804 27872
rect 27759 27832 27804 27860
rect 27798 27820 27804 27832
rect 27856 27820 27862 27872
rect 28810 27860 28816 27872
rect 28771 27832 28816 27860
rect 28810 27820 28816 27832
rect 28868 27820 28874 27872
rect 28902 27820 28908 27872
rect 28960 27860 28966 27872
rect 31938 27860 31944 27872
rect 28960 27832 31944 27860
rect 28960 27820 28966 27832
rect 31938 27820 31944 27832
rect 31996 27820 32002 27872
rect 33226 27820 33232 27872
rect 33284 27860 33290 27872
rect 35253 27863 35311 27869
rect 35253 27860 35265 27863
rect 33284 27832 35265 27860
rect 33284 27820 33290 27832
rect 35253 27829 35265 27832
rect 35299 27829 35311 27863
rect 35253 27823 35311 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 3970 27616 3976 27668
rect 4028 27656 4034 27668
rect 4430 27656 4436 27668
rect 4028 27628 4436 27656
rect 4028 27616 4034 27628
rect 4430 27616 4436 27628
rect 4488 27616 4494 27668
rect 4540 27628 4752 27656
rect 4249 27591 4307 27597
rect 4249 27557 4261 27591
rect 4295 27588 4307 27591
rect 4540 27588 4568 27628
rect 4295 27560 4568 27588
rect 4295 27557 4307 27560
rect 4249 27551 4307 27557
rect 4614 27548 4620 27600
rect 4672 27548 4678 27600
rect 4724 27588 4752 27628
rect 4798 27616 4804 27668
rect 4856 27656 4862 27668
rect 8110 27656 8116 27668
rect 4856 27628 8116 27656
rect 4856 27616 4862 27628
rect 8110 27616 8116 27628
rect 8168 27616 8174 27668
rect 13262 27656 13268 27668
rect 8220 27628 11008 27656
rect 13223 27628 13268 27656
rect 5626 27588 5632 27600
rect 4724 27560 5632 27588
rect 5626 27548 5632 27560
rect 5684 27548 5690 27600
rect 6914 27548 6920 27600
rect 6972 27588 6978 27600
rect 7009 27591 7067 27597
rect 7009 27588 7021 27591
rect 6972 27560 7021 27588
rect 6972 27548 6978 27560
rect 7009 27557 7021 27560
rect 7055 27557 7067 27591
rect 7009 27551 7067 27557
rect 7374 27548 7380 27600
rect 7432 27588 7438 27600
rect 8220 27588 8248 27628
rect 9950 27588 9956 27600
rect 7432 27560 8248 27588
rect 9911 27560 9956 27588
rect 7432 27548 7438 27560
rect 4341 27523 4399 27529
rect 4341 27489 4353 27523
rect 4387 27520 4399 27523
rect 4632 27520 4660 27548
rect 4387 27492 4660 27520
rect 4387 27489 4399 27492
rect 4341 27483 4399 27489
rect 4706 27480 4712 27532
rect 4764 27520 4770 27532
rect 5353 27523 5411 27529
rect 5353 27520 5365 27523
rect 4764 27492 5365 27520
rect 4764 27480 4770 27492
rect 5353 27489 5365 27492
rect 5399 27489 5411 27523
rect 8018 27520 8024 27532
rect 7979 27492 8024 27520
rect 5353 27483 5411 27489
rect 8018 27480 8024 27492
rect 8076 27480 8082 27532
rect 8220 27529 8248 27560
rect 9950 27548 9956 27560
rect 10008 27548 10014 27600
rect 10980 27588 11008 27628
rect 13262 27616 13268 27628
rect 13320 27616 13326 27668
rect 13998 27616 14004 27668
rect 14056 27656 14062 27668
rect 20714 27656 20720 27668
rect 14056 27628 20720 27656
rect 14056 27616 14062 27628
rect 20714 27616 20720 27628
rect 20772 27616 20778 27668
rect 21634 27656 21640 27668
rect 21008 27628 21640 27656
rect 13725 27591 13783 27597
rect 10980 27560 11376 27588
rect 8113 27523 8171 27529
rect 8113 27489 8125 27523
rect 8159 27489 8171 27523
rect 8113 27483 8171 27489
rect 8205 27523 8263 27529
rect 8205 27489 8217 27523
rect 8251 27489 8263 27523
rect 8205 27483 8263 27489
rect 4157 27455 4215 27461
rect 4157 27421 4169 27455
rect 4203 27421 4215 27455
rect 4430 27452 4436 27464
rect 4391 27424 4436 27452
rect 4157 27415 4215 27421
rect 4172 27384 4200 27415
rect 4430 27412 4436 27424
rect 4488 27412 4494 27464
rect 4614 27452 4620 27464
rect 4575 27424 4620 27452
rect 4614 27412 4620 27424
rect 4672 27412 4678 27464
rect 5074 27452 5080 27464
rect 5035 27424 5080 27452
rect 5074 27412 5080 27424
rect 5132 27412 5138 27464
rect 5258 27452 5264 27464
rect 5219 27424 5264 27452
rect 5258 27412 5264 27424
rect 5316 27412 5322 27464
rect 5442 27452 5448 27464
rect 5403 27424 5448 27452
rect 5442 27412 5448 27424
rect 5500 27412 5506 27464
rect 5629 27455 5687 27461
rect 5629 27421 5641 27455
rect 5675 27452 5687 27455
rect 5675 27424 6040 27452
rect 5675 27421 5687 27424
rect 5629 27415 5687 27421
rect 5718 27384 5724 27396
rect 4172 27356 5724 27384
rect 5718 27344 5724 27356
rect 5776 27344 5782 27396
rect 6012 27384 6040 27424
rect 6086 27412 6092 27464
rect 6144 27452 6150 27464
rect 6733 27455 6791 27461
rect 6733 27452 6745 27455
rect 6144 27424 6745 27452
rect 6144 27412 6150 27424
rect 6733 27421 6745 27424
rect 6779 27421 6791 27455
rect 7006 27452 7012 27464
rect 6967 27424 7012 27452
rect 6733 27415 6791 27421
rect 7006 27412 7012 27424
rect 7064 27412 7070 27464
rect 8128 27396 8156 27483
rect 9398 27480 9404 27532
rect 9456 27520 9462 27532
rect 9456 27492 11192 27520
rect 9456 27480 9462 27492
rect 8297 27455 8355 27461
rect 8297 27421 8309 27455
rect 8343 27450 8355 27455
rect 9214 27452 9220 27464
rect 8404 27450 9220 27452
rect 8343 27424 9220 27450
rect 8343 27422 8432 27424
rect 8343 27421 8355 27422
rect 8297 27415 8355 27421
rect 9214 27412 9220 27424
rect 9272 27412 9278 27464
rect 11164 27461 11192 27492
rect 11348 27461 11376 27560
rect 13725 27557 13737 27591
rect 13771 27588 13783 27591
rect 13814 27588 13820 27600
rect 13771 27560 13820 27588
rect 13771 27557 13783 27560
rect 13725 27551 13783 27557
rect 13814 27548 13820 27560
rect 13872 27548 13878 27600
rect 15654 27588 15660 27600
rect 15615 27560 15660 27588
rect 15654 27548 15660 27560
rect 15712 27548 15718 27600
rect 17034 27548 17040 27600
rect 17092 27588 17098 27600
rect 17313 27591 17371 27597
rect 17313 27588 17325 27591
rect 17092 27560 17325 27588
rect 17092 27548 17098 27560
rect 17313 27557 17325 27560
rect 17359 27557 17371 27591
rect 21008 27588 21036 27628
rect 21634 27616 21640 27628
rect 21692 27616 21698 27668
rect 23290 27616 23296 27668
rect 23348 27656 23354 27668
rect 26786 27656 26792 27668
rect 23348 27628 26792 27656
rect 23348 27616 23354 27628
rect 26786 27616 26792 27628
rect 26844 27616 26850 27668
rect 27154 27616 27160 27668
rect 27212 27656 27218 27668
rect 27212 27628 27844 27656
rect 27212 27616 27218 27628
rect 17313 27551 17371 27557
rect 19904 27560 21036 27588
rect 18233 27523 18291 27529
rect 18233 27489 18245 27523
rect 18279 27520 18291 27523
rect 18966 27520 18972 27532
rect 18279 27492 18972 27520
rect 18279 27489 18291 27492
rect 18233 27483 18291 27489
rect 18966 27480 18972 27492
rect 19024 27480 19030 27532
rect 10413 27455 10471 27461
rect 10413 27421 10425 27455
rect 10459 27421 10471 27455
rect 10413 27415 10471 27421
rect 11149 27455 11207 27461
rect 11149 27421 11161 27455
rect 11195 27421 11207 27455
rect 11149 27415 11207 27421
rect 11333 27455 11391 27461
rect 11333 27421 11345 27455
rect 11379 27421 11391 27455
rect 11333 27415 11391 27421
rect 6012 27356 8064 27384
rect 3970 27316 3976 27328
rect 3931 27288 3976 27316
rect 3970 27276 3976 27288
rect 4028 27276 4034 27328
rect 4522 27276 4528 27328
rect 4580 27316 4586 27328
rect 5813 27319 5871 27325
rect 5813 27316 5825 27319
rect 4580 27288 5825 27316
rect 4580 27276 4586 27288
rect 5813 27285 5825 27288
rect 5859 27285 5871 27319
rect 7834 27316 7840 27328
rect 7795 27288 7840 27316
rect 5813 27279 5871 27285
rect 7834 27276 7840 27288
rect 7892 27276 7898 27328
rect 8036 27316 8064 27356
rect 8110 27344 8116 27396
rect 8168 27384 8174 27396
rect 9030 27384 9036 27396
rect 8168 27356 9036 27384
rect 8168 27344 8174 27356
rect 9030 27344 9036 27356
rect 9088 27344 9094 27396
rect 9582 27384 9588 27396
rect 9543 27356 9588 27384
rect 9582 27344 9588 27356
rect 9640 27344 9646 27396
rect 9769 27387 9827 27393
rect 9769 27353 9781 27387
rect 9815 27384 9827 27387
rect 9858 27384 9864 27396
rect 9815 27356 9864 27384
rect 9815 27353 9827 27356
rect 9769 27347 9827 27353
rect 9858 27344 9864 27356
rect 9916 27344 9922 27396
rect 10428 27384 10456 27415
rect 11422 27412 11428 27464
rect 11480 27452 11486 27464
rect 13173 27455 13231 27461
rect 13173 27452 13185 27455
rect 11480 27424 13185 27452
rect 11480 27412 11486 27424
rect 13173 27421 13185 27424
rect 13219 27421 13231 27455
rect 13173 27415 13231 27421
rect 13541 27455 13599 27461
rect 13541 27421 13553 27455
rect 13587 27421 13599 27455
rect 13541 27415 13599 27421
rect 11790 27384 11796 27396
rect 10428 27356 11796 27384
rect 11790 27344 11796 27356
rect 11848 27344 11854 27396
rect 13556 27384 13584 27415
rect 14182 27412 14188 27464
rect 14240 27452 14246 27464
rect 14550 27461 14556 27464
rect 14277 27455 14335 27461
rect 14277 27452 14289 27455
rect 14240 27424 14289 27452
rect 14240 27412 14246 27424
rect 14277 27421 14289 27424
rect 14323 27421 14335 27455
rect 14544 27452 14556 27461
rect 14511 27424 14556 27452
rect 14277 27415 14335 27421
rect 14544 27415 14556 27424
rect 14550 27412 14556 27415
rect 14608 27412 14614 27464
rect 17497 27455 17555 27461
rect 17497 27421 17509 27455
rect 17543 27421 17555 27455
rect 17497 27415 17555 27421
rect 17589 27455 17647 27461
rect 17589 27421 17601 27455
rect 17635 27452 17647 27455
rect 17678 27452 17684 27464
rect 17635 27424 17684 27452
rect 17635 27421 17647 27424
rect 17589 27415 17647 27421
rect 17512 27384 17540 27415
rect 17678 27412 17684 27424
rect 17736 27412 17742 27464
rect 18141 27455 18199 27461
rect 18141 27421 18153 27455
rect 18187 27452 18199 27455
rect 18874 27452 18880 27464
rect 18187 27424 18880 27452
rect 18187 27421 18199 27424
rect 18141 27415 18199 27421
rect 18874 27412 18880 27424
rect 18932 27412 18938 27464
rect 19058 27412 19064 27464
rect 19116 27452 19122 27464
rect 19429 27455 19487 27461
rect 19429 27452 19441 27455
rect 19116 27424 19441 27452
rect 19116 27412 19122 27424
rect 19429 27421 19441 27424
rect 19475 27421 19487 27455
rect 19429 27415 19487 27421
rect 18322 27384 18328 27396
rect 13556 27356 17448 27384
rect 17512 27356 18328 27384
rect 10134 27316 10140 27328
rect 8036 27288 10140 27316
rect 10134 27276 10140 27288
rect 10192 27276 10198 27328
rect 10594 27316 10600 27328
rect 10555 27288 10600 27316
rect 10594 27276 10600 27288
rect 10652 27276 10658 27328
rect 11238 27316 11244 27328
rect 11199 27288 11244 27316
rect 11238 27276 11244 27288
rect 11296 27276 11302 27328
rect 17420 27316 17448 27356
rect 18322 27344 18328 27356
rect 18380 27384 18386 27396
rect 19150 27384 19156 27396
rect 18380 27356 19156 27384
rect 18380 27344 18386 27356
rect 19150 27344 19156 27356
rect 19208 27344 19214 27396
rect 19904 27384 19932 27560
rect 21910 27548 21916 27600
rect 21968 27588 21974 27600
rect 24029 27591 24087 27597
rect 24029 27588 24041 27591
rect 21968 27560 24041 27588
rect 21968 27548 21974 27560
rect 24029 27557 24041 27560
rect 24075 27557 24087 27591
rect 24029 27551 24087 27557
rect 25866 27548 25872 27600
rect 25924 27588 25930 27600
rect 25924 27560 27752 27588
rect 25924 27548 25930 27560
rect 22112 27492 22304 27520
rect 20070 27412 20076 27464
rect 20128 27452 20134 27464
rect 20165 27455 20223 27461
rect 20165 27452 20177 27455
rect 20128 27424 20177 27452
rect 20128 27412 20134 27424
rect 20165 27421 20177 27424
rect 20211 27421 20223 27455
rect 20165 27415 20223 27421
rect 21085 27455 21143 27461
rect 21085 27421 21097 27455
rect 21131 27451 21143 27455
rect 22112 27452 22140 27492
rect 21192 27451 22140 27452
rect 21131 27424 22140 27451
rect 21131 27423 21220 27424
rect 21131 27421 21143 27423
rect 21085 27415 21143 27421
rect 19981 27387 20039 27393
rect 19981 27384 19993 27387
rect 19904 27356 19993 27384
rect 19981 27353 19993 27356
rect 20027 27353 20039 27387
rect 19981 27347 20039 27353
rect 21637 27387 21695 27393
rect 21637 27353 21649 27387
rect 21683 27384 21695 27387
rect 21910 27384 21916 27396
rect 21683 27356 21916 27384
rect 21683 27353 21695 27356
rect 21637 27347 21695 27353
rect 21910 27344 21916 27356
rect 21968 27344 21974 27396
rect 22276 27384 22304 27492
rect 24118 27480 24124 27532
rect 24176 27520 24182 27532
rect 25590 27520 25596 27532
rect 24176 27492 25596 27520
rect 24176 27480 24182 27492
rect 25590 27480 25596 27492
rect 25648 27480 25654 27532
rect 26237 27523 26295 27529
rect 26237 27489 26249 27523
rect 26283 27520 26295 27523
rect 26283 27492 27476 27520
rect 26283 27489 26295 27492
rect 26237 27483 26295 27489
rect 22738 27452 22744 27464
rect 22699 27424 22744 27452
rect 22738 27412 22744 27424
rect 22796 27412 22802 27464
rect 23474 27452 23480 27464
rect 23435 27424 23480 27452
rect 23474 27412 23480 27424
rect 23532 27412 23538 27464
rect 25498 27412 25504 27464
rect 25556 27452 25562 27464
rect 26418 27452 26424 27464
rect 25556 27424 26424 27452
rect 25556 27412 25562 27424
rect 26418 27412 26424 27424
rect 26476 27452 26482 27464
rect 26513 27455 26571 27461
rect 26513 27452 26525 27455
rect 26476 27424 26525 27452
rect 26476 27412 26482 27424
rect 26513 27421 26525 27424
rect 26559 27421 26571 27455
rect 26513 27415 26571 27421
rect 26602 27449 26660 27455
rect 26602 27430 26614 27449
rect 26648 27430 26660 27449
rect 23201 27387 23259 27393
rect 23201 27384 23213 27387
rect 22276 27356 23213 27384
rect 23201 27353 23213 27356
rect 23247 27384 23259 27387
rect 24486 27384 24492 27396
rect 23247 27356 24492 27384
rect 23247 27353 23259 27356
rect 23201 27347 23259 27353
rect 24486 27344 24492 27356
rect 24544 27344 24550 27396
rect 26602 27378 26608 27430
rect 26660 27378 26666 27430
rect 26694 27412 26700 27464
rect 26752 27452 26758 27464
rect 26752 27424 26797 27452
rect 26752 27412 26758 27424
rect 26878 27412 26884 27464
rect 26936 27452 26942 27464
rect 26936 27424 26981 27452
rect 26936 27412 26942 27424
rect 18414 27316 18420 27328
rect 17420 27288 18420 27316
rect 18414 27276 18420 27288
rect 18472 27276 18478 27328
rect 18506 27276 18512 27328
rect 18564 27316 18570 27328
rect 19613 27319 19671 27325
rect 19613 27316 19625 27319
rect 18564 27288 19625 27316
rect 18564 27276 18570 27288
rect 19613 27285 19625 27288
rect 19659 27285 19671 27319
rect 19613 27279 19671 27285
rect 20073 27319 20131 27325
rect 20073 27285 20085 27319
rect 20119 27316 20131 27319
rect 25774 27316 25780 27328
rect 20119 27288 25780 27316
rect 20119 27285 20131 27288
rect 20073 27279 20131 27285
rect 25774 27276 25780 27288
rect 25832 27276 25838 27328
rect 27246 27276 27252 27328
rect 27304 27316 27310 27328
rect 27341 27319 27399 27325
rect 27341 27316 27353 27319
rect 27304 27288 27353 27316
rect 27304 27276 27310 27288
rect 27341 27285 27353 27288
rect 27387 27285 27399 27319
rect 27448 27316 27476 27492
rect 27614 27452 27620 27464
rect 27575 27424 27620 27452
rect 27614 27412 27620 27424
rect 27672 27412 27678 27464
rect 27724 27461 27752 27560
rect 27816 27461 27844 27628
rect 31294 27616 31300 27668
rect 31352 27656 31358 27668
rect 31481 27659 31539 27665
rect 31481 27656 31493 27659
rect 31352 27628 31493 27656
rect 31352 27616 31358 27628
rect 31481 27625 31493 27628
rect 31527 27625 31539 27659
rect 31481 27619 31539 27625
rect 30374 27548 30380 27600
rect 30432 27588 30438 27600
rect 35526 27588 35532 27600
rect 30432 27560 35532 27588
rect 30432 27548 30438 27560
rect 35526 27548 35532 27560
rect 35584 27548 35590 27600
rect 29270 27480 29276 27532
rect 29328 27520 29334 27532
rect 29917 27523 29975 27529
rect 29917 27520 29929 27523
rect 29328 27492 29929 27520
rect 29328 27480 29334 27492
rect 29917 27489 29929 27492
rect 29963 27489 29975 27523
rect 29917 27483 29975 27489
rect 30098 27480 30104 27532
rect 30156 27520 30162 27532
rect 30156 27492 31156 27520
rect 30156 27480 30162 27492
rect 27709 27455 27767 27461
rect 27709 27421 27721 27455
rect 27755 27421 27767 27455
rect 27709 27415 27767 27421
rect 27801 27455 27859 27461
rect 27801 27421 27813 27455
rect 27847 27421 27859 27455
rect 27801 27415 27859 27421
rect 27985 27455 28043 27461
rect 27985 27421 27997 27455
rect 28031 27421 28043 27455
rect 27985 27415 28043 27421
rect 28000 27316 28028 27415
rect 28442 27412 28448 27464
rect 28500 27452 28506 27464
rect 28813 27455 28871 27461
rect 28813 27452 28825 27455
rect 28500 27424 28825 27452
rect 28500 27412 28506 27424
rect 28813 27421 28825 27424
rect 28859 27421 28871 27455
rect 28813 27415 28871 27421
rect 28902 27412 28908 27464
rect 28960 27452 28966 27464
rect 30009 27455 30067 27461
rect 30009 27452 30021 27455
rect 28960 27424 30021 27452
rect 28960 27412 28966 27424
rect 30009 27421 30021 27424
rect 30055 27421 30067 27455
rect 30009 27415 30067 27421
rect 28629 27387 28687 27393
rect 28629 27353 28641 27387
rect 28675 27384 28687 27387
rect 29086 27384 29092 27396
rect 28675 27356 29092 27384
rect 28675 27353 28687 27356
rect 28629 27347 28687 27353
rect 29086 27344 29092 27356
rect 29144 27344 29150 27396
rect 29181 27387 29239 27393
rect 29181 27353 29193 27387
rect 29227 27384 29239 27387
rect 30116 27384 30144 27480
rect 30377 27455 30435 27461
rect 30377 27421 30389 27455
rect 30423 27452 30435 27455
rect 30466 27452 30472 27464
rect 30423 27424 30472 27452
rect 30423 27421 30435 27424
rect 30377 27415 30435 27421
rect 30466 27412 30472 27424
rect 30524 27412 30530 27464
rect 30837 27455 30895 27461
rect 30837 27421 30849 27455
rect 30883 27421 30895 27455
rect 30837 27415 30895 27421
rect 30282 27384 30288 27396
rect 29227 27356 30144 27384
rect 30243 27356 30288 27384
rect 29227 27353 29239 27356
rect 29181 27347 29239 27353
rect 30282 27344 30288 27356
rect 30340 27344 30346 27396
rect 27448 27288 28028 27316
rect 27341 27279 27399 27285
rect 28442 27276 28448 27328
rect 28500 27316 28506 27328
rect 29362 27316 29368 27328
rect 28500 27288 29368 27316
rect 28500 27276 28506 27288
rect 29362 27276 29368 27288
rect 29420 27276 29426 27328
rect 29730 27316 29736 27328
rect 29691 27288 29736 27316
rect 29730 27276 29736 27288
rect 29788 27276 29794 27328
rect 30006 27276 30012 27328
rect 30064 27316 30070 27328
rect 30852 27316 30880 27415
rect 30926 27412 30932 27464
rect 30984 27452 30990 27464
rect 31128 27461 31156 27492
rect 31202 27480 31208 27532
rect 31260 27480 31266 27532
rect 34790 27520 34796 27532
rect 32324 27492 34796 27520
rect 31113 27455 31171 27461
rect 30984 27424 31029 27452
rect 30984 27412 30990 27424
rect 31113 27421 31125 27455
rect 31159 27421 31171 27455
rect 31220 27452 31248 27480
rect 32324 27461 32352 27492
rect 34790 27480 34796 27492
rect 34848 27520 34854 27532
rect 35802 27520 35808 27532
rect 34848 27492 35808 27520
rect 34848 27480 34854 27492
rect 35802 27480 35808 27492
rect 35860 27480 35866 27532
rect 31302 27455 31360 27461
rect 31302 27452 31314 27455
rect 31220 27424 31314 27452
rect 31113 27415 31171 27421
rect 31302 27421 31314 27424
rect 31348 27421 31360 27455
rect 31941 27455 31999 27461
rect 31941 27452 31953 27455
rect 31302 27415 31360 27421
rect 31726 27424 31953 27452
rect 31202 27344 31208 27396
rect 31260 27384 31266 27396
rect 31260 27356 31305 27384
rect 31260 27344 31266 27356
rect 30064 27288 30880 27316
rect 30064 27276 30070 27288
rect 30926 27276 30932 27328
rect 30984 27316 30990 27328
rect 31726 27316 31754 27424
rect 31941 27421 31953 27424
rect 31987 27421 31999 27455
rect 31941 27415 31999 27421
rect 32309 27455 32367 27461
rect 32309 27421 32321 27455
rect 32355 27421 32367 27455
rect 32309 27415 32367 27421
rect 32858 27412 32864 27464
rect 32916 27452 32922 27464
rect 32953 27455 33011 27461
rect 32953 27452 32965 27455
rect 32916 27424 32965 27452
rect 32916 27412 32922 27424
rect 32953 27421 32965 27424
rect 32999 27421 33011 27455
rect 32953 27415 33011 27421
rect 33137 27455 33195 27461
rect 33137 27421 33149 27455
rect 33183 27421 33195 27455
rect 36906 27452 36912 27464
rect 36867 27424 36912 27452
rect 33137 27415 33195 27421
rect 32030 27344 32036 27396
rect 32088 27384 32094 27396
rect 32125 27387 32183 27393
rect 32125 27384 32137 27387
rect 32088 27356 32137 27384
rect 32088 27344 32094 27356
rect 32125 27353 32137 27356
rect 32171 27353 32183 27387
rect 32125 27347 32183 27353
rect 32214 27344 32220 27396
rect 32272 27384 32278 27396
rect 32272 27356 32317 27384
rect 32272 27344 32278 27356
rect 32766 27344 32772 27396
rect 32824 27384 32830 27396
rect 33152 27384 33180 27415
rect 36906 27412 36912 27424
rect 36964 27412 36970 27464
rect 37090 27412 37096 27464
rect 37148 27452 37154 27464
rect 37829 27455 37887 27461
rect 37829 27452 37841 27455
rect 37148 27424 37841 27452
rect 37148 27412 37154 27424
rect 37829 27421 37841 27424
rect 37875 27421 37887 27455
rect 37829 27415 37887 27421
rect 37182 27384 37188 27396
rect 32824 27356 33180 27384
rect 37143 27356 37188 27384
rect 32824 27344 32830 27356
rect 37182 27344 37188 27356
rect 37240 27344 37246 27396
rect 38102 27384 38108 27396
rect 38063 27356 38108 27384
rect 38102 27344 38108 27356
rect 38160 27344 38166 27396
rect 32490 27316 32496 27328
rect 30984 27288 31754 27316
rect 32451 27288 32496 27316
rect 30984 27276 30990 27288
rect 32490 27276 32496 27288
rect 32548 27276 32554 27328
rect 32950 27276 32956 27328
rect 33008 27316 33014 27328
rect 33045 27319 33103 27325
rect 33045 27316 33057 27319
rect 33008 27288 33057 27316
rect 33008 27276 33014 27288
rect 33045 27285 33057 27288
rect 33091 27285 33103 27319
rect 33045 27279 33103 27285
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 4157 27115 4215 27121
rect 4157 27081 4169 27115
rect 4203 27112 4215 27115
rect 4430 27112 4436 27124
rect 4203 27084 4436 27112
rect 4203 27081 4215 27084
rect 4157 27075 4215 27081
rect 4430 27072 4436 27084
rect 4488 27112 4494 27124
rect 16574 27112 16580 27124
rect 4488 27084 16580 27112
rect 4488 27072 4494 27084
rect 16574 27072 16580 27084
rect 16632 27072 16638 27124
rect 20073 27115 20131 27121
rect 20073 27081 20085 27115
rect 20119 27112 20131 27115
rect 20162 27112 20168 27124
rect 20119 27084 20168 27112
rect 20119 27081 20131 27084
rect 20073 27075 20131 27081
rect 20162 27072 20168 27084
rect 20220 27072 20226 27124
rect 22465 27115 22523 27121
rect 22465 27081 22477 27115
rect 22511 27112 22523 27115
rect 24670 27112 24676 27124
rect 22511 27084 24676 27112
rect 22511 27081 22523 27084
rect 22465 27075 22523 27081
rect 24670 27072 24676 27084
rect 24728 27072 24734 27124
rect 24765 27115 24823 27121
rect 24765 27081 24777 27115
rect 24811 27112 24823 27115
rect 24811 27084 25452 27112
rect 24811 27081 24823 27084
rect 24765 27075 24823 27081
rect 3044 27047 3102 27053
rect 3044 27013 3056 27047
rect 3090 27044 3102 27047
rect 3970 27044 3976 27056
rect 3090 27016 3976 27044
rect 3090 27013 3102 27016
rect 3044 27007 3102 27013
rect 3970 27004 3976 27016
rect 4028 27004 4034 27056
rect 4522 27004 4528 27056
rect 4580 27044 4586 27056
rect 5077 27047 5135 27053
rect 5077 27044 5089 27047
rect 4580 27016 5089 27044
rect 4580 27004 4586 27016
rect 5077 27013 5089 27016
rect 5123 27013 5135 27047
rect 5077 27007 5135 27013
rect 5166 27004 5172 27056
rect 5224 27044 5230 27056
rect 20990 27044 20996 27056
rect 5224 27016 13676 27044
rect 5224 27004 5230 27016
rect 2774 26976 2780 26988
rect 2735 26948 2780 26976
rect 2774 26936 2780 26948
rect 2832 26936 2838 26988
rect 5537 26979 5595 26985
rect 5537 26945 5549 26979
rect 5583 26976 5595 26979
rect 5718 26976 5724 26988
rect 5583 26948 5724 26976
rect 5583 26945 5595 26948
rect 5537 26939 5595 26945
rect 5718 26936 5724 26948
rect 5776 26936 5782 26988
rect 6454 26936 6460 26988
rect 6512 26976 6518 26988
rect 7009 26979 7067 26985
rect 6512 26948 6960 26976
rect 6512 26936 6518 26948
rect 5350 26908 5356 26920
rect 5311 26880 5356 26908
rect 5350 26868 5356 26880
rect 5408 26908 5414 26920
rect 6822 26908 6828 26920
rect 5408 26880 6316 26908
rect 6783 26880 6828 26908
rect 5408 26868 5414 26880
rect 4982 26800 4988 26852
rect 5040 26840 5046 26852
rect 5721 26843 5779 26849
rect 5721 26840 5733 26843
rect 5040 26812 5733 26840
rect 5040 26800 5046 26812
rect 5721 26809 5733 26812
rect 5767 26809 5779 26843
rect 6288 26840 6316 26880
rect 6822 26868 6828 26880
rect 6880 26868 6886 26920
rect 6932 26908 6960 26948
rect 7009 26945 7021 26979
rect 7055 26976 7067 26979
rect 8110 26976 8116 26988
rect 7055 26948 8116 26976
rect 7055 26945 7067 26948
rect 7009 26939 7067 26945
rect 8110 26936 8116 26948
rect 8168 26936 8174 26988
rect 8478 26976 8484 26988
rect 8439 26948 8484 26976
rect 8478 26936 8484 26948
rect 8536 26936 8542 26988
rect 8573 26979 8631 26985
rect 8573 26945 8585 26979
rect 8619 26976 8631 26979
rect 9217 26979 9275 26985
rect 9217 26976 9229 26979
rect 8619 26948 9229 26976
rect 8619 26945 8631 26948
rect 8573 26939 8631 26945
rect 9217 26945 9229 26948
rect 9263 26945 9275 26979
rect 9217 26939 9275 26945
rect 9401 26979 9459 26985
rect 9401 26945 9413 26979
rect 9447 26976 9459 26979
rect 9950 26976 9956 26988
rect 9447 26948 9956 26976
rect 9447 26945 9459 26948
rect 9401 26939 9459 26945
rect 8588 26908 8616 26939
rect 9950 26936 9956 26948
rect 10008 26936 10014 26988
rect 10781 26979 10839 26985
rect 10781 26945 10793 26979
rect 10827 26976 10839 26979
rect 11974 26976 11980 26988
rect 10827 26948 11980 26976
rect 10827 26945 10839 26948
rect 10781 26939 10839 26945
rect 11974 26936 11980 26948
rect 12032 26936 12038 26988
rect 13262 26936 13268 26988
rect 13320 26976 13326 26988
rect 13648 26985 13676 27016
rect 18156 27016 20996 27044
rect 13357 26979 13415 26985
rect 13357 26976 13369 26979
rect 13320 26948 13369 26976
rect 13320 26936 13326 26948
rect 13357 26945 13369 26948
rect 13403 26945 13415 26979
rect 13357 26939 13415 26945
rect 13541 26979 13599 26985
rect 13541 26945 13553 26979
rect 13587 26945 13599 26979
rect 13541 26939 13599 26945
rect 13633 26979 13691 26985
rect 13633 26945 13645 26979
rect 13679 26945 13691 26979
rect 13633 26939 13691 26945
rect 14369 26979 14427 26985
rect 14369 26945 14381 26979
rect 14415 26976 14427 26979
rect 14458 26976 14464 26988
rect 14415 26948 14464 26976
rect 14415 26945 14427 26948
rect 14369 26939 14427 26945
rect 6932 26880 8616 26908
rect 9122 26868 9128 26920
rect 9180 26908 9186 26920
rect 10873 26911 10931 26917
rect 10873 26908 10885 26911
rect 9180 26880 10885 26908
rect 9180 26868 9186 26880
rect 10873 26877 10885 26880
rect 10919 26877 10931 26911
rect 10873 26871 10931 26877
rect 10962 26868 10968 26920
rect 11020 26908 11026 26920
rect 13556 26908 13584 26939
rect 14458 26936 14464 26948
rect 14516 26976 14522 26988
rect 16390 26976 16396 26988
rect 14516 26948 16396 26976
rect 14516 26936 14522 26948
rect 16390 26936 16396 26948
rect 16448 26936 16454 26988
rect 17034 26976 17040 26988
rect 16995 26948 17040 26976
rect 17034 26936 17040 26948
rect 17092 26936 17098 26988
rect 17310 26976 17316 26988
rect 17271 26948 17316 26976
rect 17310 26936 17316 26948
rect 17368 26936 17374 26988
rect 17678 26936 17684 26988
rect 17736 26976 17742 26988
rect 18156 26985 18184 27016
rect 20990 27004 20996 27016
rect 21048 27004 21054 27056
rect 22002 27044 22008 27056
rect 21963 27016 22008 27044
rect 22002 27004 22008 27016
rect 22060 27004 22066 27056
rect 22370 27044 22376 27056
rect 22204 27016 22376 27044
rect 17865 26979 17923 26985
rect 17865 26976 17877 26979
rect 17736 26948 17877 26976
rect 17736 26936 17742 26948
rect 17865 26945 17877 26948
rect 17911 26945 17923 26979
rect 17865 26939 17923 26945
rect 18141 26979 18199 26985
rect 18141 26945 18153 26979
rect 18187 26945 18199 26979
rect 18141 26939 18199 26945
rect 18877 26979 18935 26985
rect 18877 26945 18889 26979
rect 18923 26976 18935 26979
rect 19150 26976 19156 26988
rect 18923 26948 19156 26976
rect 18923 26945 18935 26948
rect 18877 26939 18935 26945
rect 19150 26936 19156 26948
rect 19208 26936 19214 26988
rect 19245 26979 19303 26985
rect 19245 26945 19257 26979
rect 19291 26945 19303 26979
rect 19978 26976 19984 26988
rect 19939 26948 19984 26976
rect 19245 26939 19303 26945
rect 14274 26908 14280 26920
rect 11020 26880 14280 26908
rect 11020 26868 11026 26880
rect 14274 26868 14280 26880
rect 14332 26868 14338 26920
rect 14642 26908 14648 26920
rect 14603 26880 14648 26908
rect 14642 26868 14648 26880
rect 14700 26868 14706 26920
rect 17218 26908 17224 26920
rect 17179 26880 17224 26908
rect 17218 26868 17224 26880
rect 17276 26868 17282 26920
rect 18690 26908 18696 26920
rect 17420 26880 18696 26908
rect 7193 26843 7251 26849
rect 7193 26840 7205 26843
rect 6288 26812 7205 26840
rect 5721 26803 5779 26809
rect 7193 26809 7205 26812
rect 7239 26809 7251 26843
rect 8662 26840 8668 26852
rect 8575 26812 8668 26840
rect 7193 26803 7251 26809
rect 8662 26800 8668 26812
rect 8720 26840 8726 26852
rect 9582 26840 9588 26852
rect 8720 26812 9588 26840
rect 8720 26800 8726 26812
rect 9582 26800 9588 26812
rect 9640 26800 9646 26852
rect 9858 26800 9864 26852
rect 9916 26840 9922 26852
rect 10778 26840 10784 26852
rect 9916 26812 10784 26840
rect 9916 26800 9922 26812
rect 10778 26800 10784 26812
rect 10836 26840 10842 26852
rect 11882 26840 11888 26852
rect 10836 26812 11888 26840
rect 10836 26800 10842 26812
rect 11882 26800 11888 26812
rect 11940 26800 11946 26852
rect 17126 26840 17132 26852
rect 17039 26812 17132 26840
rect 17126 26800 17132 26812
rect 17184 26840 17190 26852
rect 17420 26840 17448 26880
rect 18690 26868 18696 26880
rect 18748 26868 18754 26920
rect 18966 26868 18972 26920
rect 19024 26908 19030 26920
rect 19061 26911 19119 26917
rect 19061 26908 19073 26911
rect 19024 26880 19073 26908
rect 19024 26868 19030 26880
rect 19061 26877 19073 26880
rect 19107 26877 19119 26911
rect 19260 26908 19288 26939
rect 19978 26936 19984 26948
rect 20036 26936 20042 26988
rect 20162 26976 20168 26988
rect 20123 26948 20168 26976
rect 20162 26936 20168 26948
rect 20220 26936 20226 26988
rect 20806 26976 20812 26988
rect 20767 26948 20812 26976
rect 20806 26936 20812 26948
rect 20864 26936 20870 26988
rect 22204 26976 22232 27016
rect 22370 27004 22376 27016
rect 22428 27044 22434 27056
rect 23382 27044 23388 27056
rect 22428 27016 23388 27044
rect 22428 27004 22434 27016
rect 23382 27004 23388 27016
rect 23440 27004 23446 27056
rect 23474 27004 23480 27056
rect 23532 27044 23538 27056
rect 24026 27044 24032 27056
rect 23532 27016 24032 27044
rect 23532 27004 23538 27016
rect 24026 27004 24032 27016
rect 24084 27044 24090 27056
rect 24084 27016 24808 27044
rect 24084 27004 24090 27016
rect 21008 26948 22232 26976
rect 22281 26979 22339 26985
rect 20180 26908 20208 26936
rect 20898 26908 20904 26920
rect 19260 26880 20208 26908
rect 20859 26880 20904 26908
rect 19061 26871 19119 26877
rect 20898 26868 20904 26880
rect 20956 26868 20962 26920
rect 17184 26812 17448 26840
rect 17184 26800 17190 26812
rect 17494 26800 17500 26852
rect 17552 26840 17558 26852
rect 18141 26843 18199 26849
rect 18141 26840 18153 26843
rect 17552 26812 18153 26840
rect 17552 26800 17558 26812
rect 18141 26809 18153 26812
rect 18187 26809 18199 26843
rect 18141 26803 18199 26809
rect 19153 26843 19211 26849
rect 19153 26809 19165 26843
rect 19199 26840 19211 26843
rect 21008 26840 21036 26948
rect 22281 26945 22293 26979
rect 22327 26976 22339 26979
rect 22554 26976 22560 26988
rect 22327 26948 22560 26976
rect 22327 26945 22339 26948
rect 22281 26939 22339 26945
rect 22554 26936 22560 26948
rect 22612 26936 22618 26988
rect 22738 26936 22744 26988
rect 22796 26976 22802 26988
rect 22925 26979 22983 26985
rect 22925 26976 22937 26979
rect 22796 26948 22937 26976
rect 22796 26936 22802 26948
rect 22925 26945 22937 26948
rect 22971 26945 22983 26979
rect 22925 26939 22983 26945
rect 23201 26979 23259 26985
rect 23201 26945 23213 26979
rect 23247 26945 23259 26979
rect 23201 26939 23259 26945
rect 22097 26911 22155 26917
rect 22097 26877 22109 26911
rect 22143 26877 22155 26911
rect 22097 26871 22155 26877
rect 19199 26812 21036 26840
rect 21177 26843 21235 26849
rect 19199 26809 19211 26812
rect 19153 26803 19211 26809
rect 21177 26809 21189 26843
rect 21223 26840 21235 26843
rect 22112 26840 22140 26871
rect 22186 26868 22192 26920
rect 22244 26908 22250 26920
rect 23017 26911 23075 26917
rect 23017 26908 23029 26911
rect 22244 26880 23029 26908
rect 22244 26868 22250 26880
rect 23017 26877 23029 26880
rect 23063 26877 23075 26911
rect 23017 26871 23075 26877
rect 23106 26868 23112 26920
rect 23164 26868 23170 26920
rect 23216 26908 23244 26939
rect 24302 26936 24308 26988
rect 24360 26976 24366 26988
rect 24780 26985 24808 27016
rect 25424 26988 25452 27084
rect 25590 27072 25596 27124
rect 25648 27112 25654 27124
rect 26329 27115 26387 27121
rect 25648 27084 26280 27112
rect 25648 27072 25654 27084
rect 25774 27004 25780 27056
rect 25832 27044 25838 27056
rect 26145 27047 26203 27053
rect 26145 27044 26157 27047
rect 25832 27016 26157 27044
rect 25832 27004 25838 27016
rect 26145 27013 26157 27016
rect 26191 27013 26203 27047
rect 26252 27044 26280 27084
rect 26329 27081 26341 27115
rect 26375 27112 26387 27115
rect 27798 27112 27804 27124
rect 26375 27084 27804 27112
rect 26375 27081 26387 27084
rect 26329 27075 26387 27081
rect 27798 27072 27804 27084
rect 27856 27072 27862 27124
rect 29086 27112 29092 27124
rect 29047 27084 29092 27112
rect 29086 27072 29092 27084
rect 29144 27112 29150 27124
rect 31662 27112 31668 27124
rect 29144 27084 31668 27112
rect 29144 27072 29150 27084
rect 31662 27072 31668 27084
rect 31720 27072 31726 27124
rect 35986 27112 35992 27124
rect 34716 27084 35992 27112
rect 28442 27044 28448 27056
rect 26252 27016 28448 27044
rect 26145 27007 26203 27013
rect 24581 26979 24639 26985
rect 24581 26976 24593 26979
rect 24360 26948 24593 26976
rect 24360 26936 24366 26948
rect 24581 26945 24593 26948
rect 24627 26945 24639 26979
rect 24581 26939 24639 26945
rect 24765 26979 24823 26985
rect 24765 26945 24777 26979
rect 24811 26945 24823 26979
rect 25406 26976 25412 26988
rect 25319 26948 25412 26976
rect 24765 26939 24823 26945
rect 25406 26936 25412 26948
rect 25464 26976 25470 26988
rect 26694 26976 26700 26988
rect 25464 26948 26700 26976
rect 25464 26936 25470 26948
rect 26694 26936 26700 26948
rect 26752 26936 26758 26988
rect 27264 26985 27292 27016
rect 28442 27004 28448 27016
rect 28500 27004 28506 27056
rect 28626 27004 28632 27056
rect 28684 27044 28690 27056
rect 28684 27016 31340 27044
rect 28684 27004 28690 27016
rect 27249 26979 27307 26985
rect 27249 26945 27261 26979
rect 27295 26945 27307 26979
rect 28077 26979 28135 26985
rect 28077 26976 28089 26979
rect 27249 26939 27307 26945
rect 27540 26948 28089 26976
rect 25958 26908 25964 26920
rect 23216 26880 25964 26908
rect 25958 26868 25964 26880
rect 26016 26868 26022 26920
rect 26142 26868 26148 26920
rect 26200 26908 26206 26920
rect 27540 26908 27568 26948
rect 28077 26945 28089 26948
rect 28123 26976 28135 26979
rect 28994 26976 29000 26988
rect 28123 26948 29000 26976
rect 28123 26945 28135 26948
rect 28077 26939 28135 26945
rect 28994 26936 29000 26948
rect 29052 26976 29058 26988
rect 29089 26979 29147 26985
rect 29089 26976 29101 26979
rect 29052 26948 29101 26976
rect 29052 26936 29058 26948
rect 29089 26945 29101 26948
rect 29135 26945 29147 26979
rect 29089 26939 29147 26945
rect 29733 26979 29791 26985
rect 29733 26945 29745 26979
rect 29779 26945 29791 26979
rect 29733 26939 29791 26945
rect 26200 26880 27568 26908
rect 26200 26868 26206 26880
rect 27706 26868 27712 26920
rect 27764 26908 27770 26920
rect 29748 26908 29776 26939
rect 30650 26936 30656 26988
rect 30708 26976 30714 26988
rect 31021 26979 31079 26985
rect 31021 26976 31033 26979
rect 30708 26948 31033 26976
rect 30708 26936 30714 26948
rect 31021 26945 31033 26948
rect 31067 26945 31079 26979
rect 31021 26939 31079 26945
rect 31113 26979 31171 26985
rect 31113 26945 31125 26979
rect 31159 26976 31171 26979
rect 31202 26976 31208 26988
rect 31159 26948 31208 26976
rect 31159 26945 31171 26948
rect 31113 26939 31171 26945
rect 27764 26880 29776 26908
rect 27764 26868 27770 26880
rect 30374 26868 30380 26920
rect 30432 26908 30438 26920
rect 31128 26908 31156 26939
rect 31202 26936 31208 26948
rect 31260 26936 31266 26988
rect 31312 26985 31340 27016
rect 32030 27004 32036 27056
rect 32088 27044 32094 27056
rect 32950 27053 32956 27056
rect 32088 27016 32904 27044
rect 32088 27004 32094 27016
rect 31297 26979 31355 26985
rect 31297 26945 31309 26979
rect 31343 26945 31355 26979
rect 31297 26939 31355 26945
rect 31386 26936 31392 26988
rect 31444 26976 31450 26988
rect 32674 26976 32680 26988
rect 31444 26948 31489 26976
rect 32635 26948 32680 26976
rect 31444 26936 31450 26948
rect 32674 26936 32680 26948
rect 32732 26936 32738 26988
rect 32876 26976 32904 27016
rect 32944 27007 32956 27053
rect 33008 27044 33014 27056
rect 33008 27016 33044 27044
rect 32950 27004 32956 27007
rect 33008 27004 33014 27016
rect 34716 26976 34744 27084
rect 35986 27072 35992 27084
rect 36044 27072 36050 27124
rect 36173 27115 36231 27121
rect 36173 27081 36185 27115
rect 36219 27112 36231 27115
rect 36906 27112 36912 27124
rect 36219 27084 36912 27112
rect 36219 27081 36231 27084
rect 36173 27075 36231 27081
rect 36906 27072 36912 27084
rect 36964 27112 36970 27124
rect 37921 27115 37979 27121
rect 37921 27112 37933 27115
rect 36964 27084 37933 27112
rect 36964 27072 36970 27084
rect 37921 27081 37933 27084
rect 37967 27081 37979 27115
rect 37921 27075 37979 27081
rect 37826 27044 37832 27056
rect 35176 27016 37832 27044
rect 32876 26948 34744 26976
rect 30432 26880 31156 26908
rect 34716 26908 34744 26948
rect 34790 26936 34796 26988
rect 34848 26976 34854 26988
rect 35176 26985 35204 27016
rect 37826 27004 37832 27016
rect 37884 27004 37890 27056
rect 35161 26979 35219 26985
rect 35161 26976 35173 26979
rect 34848 26948 35173 26976
rect 34848 26936 34854 26948
rect 35161 26945 35173 26948
rect 35207 26945 35219 26979
rect 35161 26939 35219 26945
rect 35345 26979 35403 26985
rect 35345 26945 35357 26979
rect 35391 26945 35403 26979
rect 35345 26939 35403 26945
rect 35437 26979 35495 26985
rect 35437 26945 35449 26979
rect 35483 26945 35495 26979
rect 35437 26939 35495 26945
rect 35529 26979 35587 26985
rect 35529 26945 35541 26979
rect 35575 26976 35587 26979
rect 35802 26976 35808 26988
rect 35575 26948 35808 26976
rect 35575 26945 35587 26948
rect 35529 26939 35587 26945
rect 35360 26908 35388 26939
rect 34716 26880 35388 26908
rect 30432 26868 30438 26880
rect 21223 26812 22140 26840
rect 21223 26809 21235 26812
rect 21177 26803 21235 26809
rect 5534 26772 5540 26784
rect 5495 26744 5540 26772
rect 5534 26732 5540 26744
rect 5592 26732 5598 26784
rect 6822 26732 6828 26784
rect 6880 26772 6886 26784
rect 7374 26772 7380 26784
rect 6880 26744 7380 26772
rect 6880 26732 6886 26744
rect 7374 26732 7380 26744
rect 7432 26732 7438 26784
rect 9214 26772 9220 26784
rect 9175 26744 9220 26772
rect 9214 26732 9220 26744
rect 9272 26732 9278 26784
rect 10413 26775 10471 26781
rect 10413 26741 10425 26775
rect 10459 26772 10471 26775
rect 10870 26772 10876 26784
rect 10459 26744 10876 26772
rect 10459 26741 10471 26744
rect 10413 26735 10471 26741
rect 10870 26732 10876 26744
rect 10928 26732 10934 26784
rect 13170 26772 13176 26784
rect 13131 26744 13176 26772
rect 13170 26732 13176 26744
rect 13228 26732 13234 26784
rect 15562 26732 15568 26784
rect 15620 26772 15626 26784
rect 16853 26775 16911 26781
rect 16853 26772 16865 26775
rect 15620 26744 16865 26772
rect 15620 26732 15626 26744
rect 16853 26741 16865 26744
rect 16899 26741 16911 26775
rect 19058 26772 19064 26784
rect 19019 26744 19064 26772
rect 16853 26735 16911 26741
rect 19058 26732 19064 26744
rect 19116 26732 19122 26784
rect 20993 26775 21051 26781
rect 20993 26741 21005 26775
rect 21039 26772 21051 26775
rect 21910 26772 21916 26784
rect 21039 26744 21916 26772
rect 21039 26741 21051 26744
rect 20993 26735 21051 26741
rect 21910 26732 21916 26744
rect 21968 26732 21974 26784
rect 22281 26775 22339 26781
rect 22281 26741 22293 26775
rect 22327 26772 22339 26775
rect 22370 26772 22376 26784
rect 22327 26744 22376 26772
rect 22327 26741 22339 26744
rect 22281 26735 22339 26741
rect 22370 26732 22376 26744
rect 22428 26732 22434 26784
rect 23124 26781 23152 26868
rect 26513 26843 26571 26849
rect 26513 26809 26525 26843
rect 26559 26840 26571 26843
rect 32122 26840 32128 26852
rect 26559 26812 32128 26840
rect 26559 26809 26571 26812
rect 26513 26803 26571 26809
rect 32122 26800 32128 26812
rect 32180 26800 32186 26852
rect 33870 26800 33876 26852
rect 33928 26840 33934 26852
rect 34057 26843 34115 26849
rect 34057 26840 34069 26843
rect 33928 26812 34069 26840
rect 33928 26800 33934 26812
rect 34057 26809 34069 26812
rect 34103 26809 34115 26843
rect 34057 26803 34115 26809
rect 34606 26800 34612 26852
rect 34664 26840 34670 26852
rect 35452 26840 35480 26939
rect 35802 26936 35808 26948
rect 35860 26936 35866 26988
rect 36354 26976 36360 26988
rect 36315 26948 36360 26976
rect 36354 26936 36360 26948
rect 36412 26936 36418 26988
rect 36630 26976 36636 26988
rect 36591 26948 36636 26976
rect 36630 26936 36636 26948
rect 36688 26936 36694 26988
rect 38010 26908 38016 26920
rect 37971 26880 38016 26908
rect 38010 26868 38016 26880
rect 38068 26868 38074 26920
rect 34664 26812 35480 26840
rect 34664 26800 34670 26812
rect 23109 26775 23167 26781
rect 23109 26741 23121 26775
rect 23155 26741 23167 26775
rect 23109 26735 23167 26741
rect 23290 26732 23296 26784
rect 23348 26772 23354 26784
rect 23385 26775 23443 26781
rect 23385 26772 23397 26775
rect 23348 26744 23397 26772
rect 23348 26732 23354 26744
rect 23385 26741 23397 26744
rect 23431 26741 23443 26775
rect 23385 26735 23443 26741
rect 24578 26732 24584 26784
rect 24636 26772 24642 26784
rect 26329 26775 26387 26781
rect 26329 26772 26341 26775
rect 24636 26744 26341 26772
rect 24636 26732 24642 26744
rect 26329 26741 26341 26744
rect 26375 26741 26387 26775
rect 26329 26735 26387 26741
rect 26878 26732 26884 26784
rect 26936 26772 26942 26784
rect 28261 26775 28319 26781
rect 28261 26772 28273 26775
rect 26936 26744 28273 26772
rect 26936 26732 26942 26744
rect 28261 26741 28273 26744
rect 28307 26772 28319 26775
rect 30742 26772 30748 26784
rect 28307 26744 30748 26772
rect 28307 26741 28319 26744
rect 28261 26735 28319 26741
rect 30742 26732 30748 26744
rect 30800 26732 30806 26784
rect 30837 26775 30895 26781
rect 30837 26741 30849 26775
rect 30883 26772 30895 26775
rect 33410 26772 33416 26784
rect 30883 26744 33416 26772
rect 30883 26741 30895 26744
rect 30837 26735 30895 26741
rect 33410 26732 33416 26744
rect 33468 26732 33474 26784
rect 35713 26775 35771 26781
rect 35713 26741 35725 26775
rect 35759 26772 35771 26775
rect 35802 26772 35808 26784
rect 35759 26744 35808 26772
rect 35759 26741 35771 26744
rect 35713 26735 35771 26741
rect 35802 26732 35808 26744
rect 35860 26732 35866 26784
rect 36538 26772 36544 26784
rect 36499 26744 36544 26772
rect 36538 26732 36544 26744
rect 36596 26732 36602 26784
rect 37458 26772 37464 26784
rect 37419 26744 37464 26772
rect 37458 26732 37464 26744
rect 37516 26732 37522 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 4522 26528 4528 26580
rect 4580 26568 4586 26580
rect 4798 26568 4804 26580
rect 4580 26540 4804 26568
rect 4580 26528 4586 26540
rect 4798 26528 4804 26540
rect 4856 26528 4862 26580
rect 4893 26571 4951 26577
rect 4893 26537 4905 26571
rect 4939 26568 4951 26571
rect 5166 26568 5172 26580
rect 4939 26540 5172 26568
rect 4939 26537 4951 26540
rect 4893 26531 4951 26537
rect 5166 26528 5172 26540
rect 5224 26528 5230 26580
rect 5534 26528 5540 26580
rect 5592 26568 5598 26580
rect 5997 26571 6055 26577
rect 5997 26568 6009 26571
rect 5592 26540 6009 26568
rect 5592 26528 5598 26540
rect 5997 26537 6009 26540
rect 6043 26537 6055 26571
rect 9122 26568 9128 26580
rect 9083 26540 9128 26568
rect 5997 26531 6055 26537
rect 9122 26528 9128 26540
rect 9180 26528 9186 26580
rect 11238 26568 11244 26580
rect 9324 26540 11244 26568
rect 4430 26460 4436 26512
rect 4488 26500 4494 26512
rect 4488 26472 5212 26500
rect 4488 26460 4494 26472
rect 4341 26435 4399 26441
rect 4341 26401 4353 26435
rect 4387 26432 4399 26435
rect 4798 26432 4804 26444
rect 4387 26404 4804 26432
rect 4387 26401 4399 26404
rect 4341 26395 4399 26401
rect 4798 26392 4804 26404
rect 4856 26432 4862 26444
rect 5077 26435 5135 26441
rect 5077 26432 5089 26435
rect 4856 26404 5089 26432
rect 4856 26392 4862 26404
rect 5077 26401 5089 26404
rect 5123 26401 5135 26435
rect 5184 26432 5212 26472
rect 5258 26460 5264 26512
rect 5316 26500 5322 26512
rect 6270 26500 6276 26512
rect 5316 26472 6276 26500
rect 5316 26460 5322 26472
rect 6270 26460 6276 26472
rect 6328 26500 6334 26512
rect 7650 26500 7656 26512
rect 6328 26472 7656 26500
rect 6328 26460 6334 26472
rect 7650 26460 7656 26472
rect 7708 26460 7714 26512
rect 7006 26432 7012 26444
rect 5184 26404 5304 26432
rect 5077 26395 5135 26401
rect 4249 26367 4307 26373
rect 4249 26333 4261 26367
rect 4295 26333 4307 26367
rect 4249 26327 4307 26333
rect 4433 26367 4491 26373
rect 4433 26333 4445 26367
rect 4479 26333 4491 26367
rect 5166 26364 5172 26376
rect 5127 26336 5172 26364
rect 4433 26327 4491 26333
rect 4264 26228 4292 26327
rect 4448 26296 4476 26327
rect 5166 26324 5172 26336
rect 5224 26324 5230 26376
rect 5276 26373 5304 26404
rect 6196 26404 7012 26432
rect 5261 26367 5319 26373
rect 5261 26333 5273 26367
rect 5307 26333 5319 26367
rect 5261 26327 5319 26333
rect 5353 26367 5411 26373
rect 5353 26333 5365 26367
rect 5399 26364 5411 26367
rect 5534 26364 5540 26376
rect 5399 26336 5540 26364
rect 5399 26333 5411 26336
rect 5353 26327 5411 26333
rect 5534 26324 5540 26336
rect 5592 26324 5598 26376
rect 6196 26364 6224 26404
rect 7006 26392 7012 26404
rect 7064 26392 7070 26444
rect 6012 26336 6224 26364
rect 6012 26305 6040 26336
rect 6270 26324 6276 26376
rect 6328 26364 6334 26376
rect 6730 26364 6736 26376
rect 6328 26336 6373 26364
rect 6691 26336 6736 26364
rect 6328 26324 6334 26336
rect 6730 26324 6736 26336
rect 6788 26324 6794 26376
rect 6917 26367 6975 26373
rect 6917 26333 6929 26367
rect 6963 26364 6975 26367
rect 7190 26364 7196 26376
rect 6963 26336 7196 26364
rect 6963 26333 6975 26336
rect 6917 26327 6975 26333
rect 7190 26324 7196 26336
rect 7248 26324 7254 26376
rect 9324 26373 9352 26540
rect 11238 26528 11244 26540
rect 11296 26528 11302 26580
rect 11974 26568 11980 26580
rect 11935 26540 11980 26568
rect 11974 26528 11980 26540
rect 12032 26568 12038 26580
rect 13262 26568 13268 26580
rect 12032 26540 12434 26568
rect 13223 26540 13268 26568
rect 12032 26528 12038 26540
rect 9674 26460 9680 26512
rect 9732 26460 9738 26512
rect 9766 26460 9772 26512
rect 9824 26500 9830 26512
rect 10134 26500 10140 26512
rect 9824 26472 10140 26500
rect 9824 26460 9830 26472
rect 10134 26460 10140 26472
rect 10192 26460 10198 26512
rect 12406 26500 12434 26540
rect 13262 26528 13268 26540
rect 13320 26528 13326 26580
rect 16666 26528 16672 26580
rect 16724 26568 16730 26580
rect 17586 26568 17592 26580
rect 16724 26540 17592 26568
rect 16724 26528 16730 26540
rect 17586 26528 17592 26540
rect 17644 26528 17650 26580
rect 18414 26528 18420 26580
rect 18472 26568 18478 26580
rect 21818 26568 21824 26580
rect 18472 26540 21824 26568
rect 18472 26528 18478 26540
rect 21818 26528 21824 26540
rect 21876 26528 21882 26580
rect 22002 26528 22008 26580
rect 22060 26568 22066 26580
rect 22281 26571 22339 26577
rect 22281 26568 22293 26571
rect 22060 26540 22293 26568
rect 22060 26528 22066 26540
rect 22281 26537 22293 26540
rect 22327 26537 22339 26571
rect 22738 26568 22744 26580
rect 22699 26540 22744 26568
rect 22281 26531 22339 26537
rect 22738 26528 22744 26540
rect 22796 26528 22802 26580
rect 27525 26571 27583 26577
rect 27525 26537 27537 26571
rect 27571 26568 27583 26571
rect 28902 26568 28908 26580
rect 27571 26540 28908 26568
rect 27571 26537 27583 26540
rect 27525 26531 27583 26537
rect 28902 26528 28908 26540
rect 28960 26528 28966 26580
rect 30190 26528 30196 26580
rect 30248 26568 30254 26580
rect 34790 26568 34796 26580
rect 30248 26540 34796 26568
rect 30248 26528 30254 26540
rect 34790 26528 34796 26540
rect 34848 26528 34854 26580
rect 35253 26571 35311 26577
rect 35253 26537 35265 26571
rect 35299 26568 35311 26571
rect 36354 26568 36360 26580
rect 35299 26540 36360 26568
rect 35299 26537 35311 26540
rect 35253 26531 35311 26537
rect 36354 26528 36360 26540
rect 36412 26528 36418 26580
rect 37826 26528 37832 26580
rect 37884 26568 37890 26580
rect 38105 26571 38163 26577
rect 38105 26568 38117 26571
rect 37884 26540 38117 26568
rect 37884 26528 37890 26540
rect 38105 26537 38117 26540
rect 38151 26537 38163 26571
rect 38105 26531 38163 26537
rect 17310 26500 17316 26512
rect 12406 26472 17316 26500
rect 17310 26460 17316 26472
rect 17368 26460 17374 26512
rect 20254 26460 20260 26512
rect 20312 26500 20318 26512
rect 20312 26472 21128 26500
rect 20312 26460 20318 26472
rect 9692 26432 9720 26460
rect 10502 26432 10508 26444
rect 9692 26404 10508 26432
rect 10502 26392 10508 26404
rect 10560 26432 10566 26444
rect 10597 26435 10655 26441
rect 10597 26432 10609 26435
rect 10560 26404 10609 26432
rect 10560 26392 10566 26404
rect 10597 26401 10609 26404
rect 10643 26401 10655 26435
rect 10597 26395 10655 26401
rect 11790 26392 11796 26444
rect 11848 26432 11854 26444
rect 12250 26432 12256 26444
rect 11848 26404 12256 26432
rect 11848 26392 11854 26404
rect 12250 26392 12256 26404
rect 12308 26432 12314 26444
rect 15657 26435 15715 26441
rect 12308 26404 13768 26432
rect 12308 26392 12314 26404
rect 9309 26367 9367 26373
rect 9309 26333 9321 26367
rect 9355 26333 9367 26367
rect 9493 26367 9551 26373
rect 9493 26354 9505 26367
rect 9539 26354 9551 26367
rect 9769 26367 9827 26373
rect 9309 26327 9367 26333
rect 5997 26299 6055 26305
rect 5997 26296 6009 26299
rect 4448 26268 6009 26296
rect 5997 26265 6009 26268
rect 6043 26265 6055 26299
rect 5997 26259 6055 26265
rect 6181 26299 6239 26305
rect 6181 26265 6193 26299
rect 6227 26296 6239 26299
rect 6825 26299 6883 26305
rect 6825 26296 6837 26299
rect 6227 26268 6837 26296
rect 6227 26265 6239 26268
rect 6181 26259 6239 26265
rect 6825 26265 6837 26268
rect 6871 26265 6883 26299
rect 6825 26259 6883 26265
rect 8478 26256 8484 26308
rect 8536 26296 8542 26308
rect 9401 26299 9459 26305
rect 9490 26302 9496 26354
rect 9548 26302 9554 26354
rect 9769 26333 9781 26367
rect 9815 26364 9827 26367
rect 9858 26364 9864 26376
rect 9815 26336 9864 26364
rect 9815 26333 9827 26336
rect 9769 26327 9827 26333
rect 9858 26324 9864 26336
rect 9916 26324 9922 26376
rect 10870 26373 10876 26376
rect 10864 26364 10876 26373
rect 10831 26336 10876 26364
rect 10864 26327 10876 26336
rect 10870 26324 10876 26327
rect 10928 26324 10934 26376
rect 13449 26367 13507 26373
rect 13449 26333 13461 26367
rect 13495 26364 13507 26367
rect 13538 26364 13544 26376
rect 13495 26336 13544 26364
rect 13495 26333 13507 26336
rect 13449 26327 13507 26333
rect 13538 26324 13544 26336
rect 13596 26324 13602 26376
rect 13740 26373 13768 26404
rect 15657 26401 15669 26435
rect 15703 26432 15715 26435
rect 18138 26432 18144 26444
rect 15703 26404 16804 26432
rect 15703 26401 15715 26404
rect 15657 26395 15715 26401
rect 13725 26367 13783 26373
rect 13725 26333 13737 26367
rect 13771 26364 13783 26367
rect 14642 26364 14648 26376
rect 13771 26336 14648 26364
rect 13771 26333 13783 26336
rect 13725 26327 13783 26333
rect 14642 26324 14648 26336
rect 14700 26324 14706 26376
rect 15562 26364 15568 26376
rect 15523 26336 15568 26364
rect 15562 26324 15568 26336
rect 15620 26324 15626 26376
rect 15933 26367 15991 26373
rect 15933 26333 15945 26367
rect 15979 26333 15991 26367
rect 15933 26327 15991 26333
rect 9401 26296 9413 26299
rect 8536 26268 9413 26296
rect 8536 26256 8542 26268
rect 9401 26265 9413 26268
rect 9447 26265 9459 26299
rect 9401 26259 9459 26265
rect 9582 26256 9588 26308
rect 9640 26305 9646 26308
rect 9640 26299 9669 26305
rect 9657 26265 9669 26299
rect 9640 26259 9669 26265
rect 13633 26299 13691 26305
rect 13633 26265 13645 26299
rect 13679 26296 13691 26299
rect 14921 26299 14979 26305
rect 13679 26268 14780 26296
rect 13679 26265 13691 26268
rect 13633 26259 13691 26265
rect 9640 26256 9646 26259
rect 4706 26228 4712 26240
rect 4264 26200 4712 26228
rect 4706 26188 4712 26200
rect 4764 26228 4770 26240
rect 5166 26228 5172 26240
rect 4764 26200 5172 26228
rect 4764 26188 4770 26200
rect 5166 26188 5172 26200
rect 5224 26188 5230 26240
rect 5258 26188 5264 26240
rect 5316 26228 5322 26240
rect 8386 26228 8392 26240
rect 5316 26200 8392 26228
rect 5316 26188 5322 26200
rect 8386 26188 8392 26200
rect 8444 26188 8450 26240
rect 14752 26228 14780 26268
rect 14921 26265 14933 26299
rect 14967 26296 14979 26299
rect 15010 26296 15016 26308
rect 14967 26268 15016 26296
rect 14967 26265 14979 26268
rect 14921 26259 14979 26265
rect 15010 26256 15016 26268
rect 15068 26256 15074 26308
rect 15102 26256 15108 26308
rect 15160 26296 15166 26308
rect 15948 26296 15976 26327
rect 16022 26324 16028 26376
rect 16080 26364 16086 26376
rect 16080 26336 16125 26364
rect 16080 26324 16086 26336
rect 15160 26268 15976 26296
rect 16776 26296 16804 26404
rect 17420 26404 18144 26432
rect 16853 26367 16911 26373
rect 16853 26333 16865 26367
rect 16899 26364 16911 26367
rect 16942 26364 16948 26376
rect 16899 26336 16948 26364
rect 16899 26333 16911 26336
rect 16853 26327 16911 26333
rect 16942 26324 16948 26336
rect 17000 26324 17006 26376
rect 17126 26364 17132 26376
rect 17087 26336 17132 26364
rect 17126 26324 17132 26336
rect 17184 26324 17190 26376
rect 17218 26324 17224 26376
rect 17276 26364 17282 26376
rect 17420 26373 17448 26404
rect 18138 26392 18144 26404
rect 18196 26392 18202 26444
rect 17405 26367 17463 26373
rect 17405 26364 17417 26367
rect 17276 26336 17417 26364
rect 17276 26324 17282 26336
rect 17405 26333 17417 26336
rect 17451 26333 17463 26367
rect 17405 26327 17463 26333
rect 17586 26324 17592 26376
rect 17644 26364 17650 26376
rect 17773 26367 17831 26373
rect 17773 26364 17785 26367
rect 17644 26336 17785 26364
rect 17644 26324 17650 26336
rect 17773 26333 17785 26336
rect 17819 26333 17831 26367
rect 20622 26364 20628 26376
rect 20583 26336 20628 26364
rect 17773 26327 17831 26333
rect 20622 26324 20628 26336
rect 20680 26324 20686 26376
rect 20714 26324 20720 26376
rect 20772 26364 20778 26376
rect 20809 26367 20867 26373
rect 20809 26364 20821 26367
rect 20772 26336 20821 26364
rect 20772 26324 20778 26336
rect 20809 26333 20821 26336
rect 20855 26333 20867 26367
rect 21100 26364 21128 26472
rect 21266 26460 21272 26512
rect 21324 26500 21330 26512
rect 21324 26472 22324 26500
rect 21324 26460 21330 26472
rect 22002 26432 22008 26444
rect 21468 26404 22008 26432
rect 21468 26373 21496 26404
rect 22002 26392 22008 26404
rect 22060 26392 22066 26444
rect 21269 26367 21327 26373
rect 21269 26364 21281 26367
rect 21100 26336 21281 26364
rect 20809 26327 20867 26333
rect 21269 26333 21281 26336
rect 21315 26333 21327 26367
rect 21269 26327 21327 26333
rect 21453 26367 21511 26373
rect 21453 26333 21465 26367
rect 21499 26333 21511 26367
rect 21453 26327 21511 26333
rect 16776 26268 17816 26296
rect 15160 26256 15166 26268
rect 15120 26228 15148 26256
rect 17788 26237 17816 26268
rect 14752 26200 15148 26228
rect 17773 26231 17831 26237
rect 17773 26197 17785 26231
rect 17819 26228 17831 26231
rect 17862 26228 17868 26240
rect 17819 26200 17868 26228
rect 17819 26197 17831 26200
rect 17773 26191 17831 26197
rect 17862 26188 17868 26200
rect 17920 26188 17926 26240
rect 20717 26231 20775 26237
rect 20717 26197 20729 26231
rect 20763 26228 20775 26231
rect 21468 26228 21496 26327
rect 21542 26324 21548 26376
rect 21600 26364 21606 26376
rect 22296 26373 22324 26472
rect 28074 26460 28080 26512
rect 28132 26500 28138 26512
rect 28626 26500 28632 26512
rect 28132 26472 28632 26500
rect 28132 26460 28138 26472
rect 28626 26460 28632 26472
rect 28684 26460 28690 26512
rect 32766 26460 32772 26512
rect 32824 26500 32830 26512
rect 34241 26503 34299 26509
rect 34241 26500 34253 26503
rect 32824 26472 34253 26500
rect 32824 26460 32830 26472
rect 34241 26469 34253 26472
rect 34287 26469 34299 26503
rect 34241 26463 34299 26469
rect 22830 26392 22836 26444
rect 22888 26432 22894 26444
rect 22888 26404 24532 26432
rect 22888 26392 22894 26404
rect 21729 26367 21787 26373
rect 21729 26364 21741 26367
rect 21600 26336 21741 26364
rect 21600 26324 21606 26336
rect 21729 26333 21741 26336
rect 21775 26333 21787 26367
rect 21729 26327 21787 26333
rect 22281 26367 22339 26373
rect 22281 26333 22293 26367
rect 22327 26333 22339 26367
rect 22281 26327 22339 26333
rect 22370 26324 22376 26376
rect 22428 26364 22434 26376
rect 22465 26367 22523 26373
rect 22465 26364 22477 26367
rect 22428 26336 22477 26364
rect 22428 26324 22434 26336
rect 22465 26333 22477 26336
rect 22511 26333 22523 26367
rect 22465 26327 22523 26333
rect 22557 26367 22615 26373
rect 22557 26333 22569 26367
rect 22603 26333 22615 26367
rect 22557 26327 22615 26333
rect 22572 26296 22600 26327
rect 23014 26324 23020 26376
rect 23072 26364 23078 26376
rect 23201 26367 23259 26373
rect 23201 26364 23213 26367
rect 23072 26336 23213 26364
rect 23072 26324 23078 26336
rect 23201 26333 23213 26336
rect 23247 26333 23259 26367
rect 23382 26364 23388 26376
rect 23343 26336 23388 26364
rect 23201 26327 23259 26333
rect 23382 26324 23388 26336
rect 23440 26324 23446 26376
rect 24504 26364 24532 26404
rect 24670 26392 24676 26444
rect 24728 26432 24734 26444
rect 24857 26435 24915 26441
rect 24857 26432 24869 26435
rect 24728 26404 24869 26432
rect 24728 26392 24734 26404
rect 24857 26401 24869 26404
rect 24903 26401 24915 26435
rect 27614 26432 27620 26444
rect 24857 26395 24915 26401
rect 25240 26404 27620 26432
rect 24578 26364 24584 26376
rect 24491 26336 24584 26364
rect 24504 26334 24584 26336
rect 24578 26324 24584 26334
rect 24636 26324 24642 26376
rect 24769 26369 24827 26375
rect 24769 26335 24781 26369
rect 24815 26335 24827 26369
rect 24769 26329 24827 26335
rect 24780 26296 24808 26329
rect 24946 26324 24952 26376
rect 25004 26364 25010 26376
rect 25004 26336 25049 26364
rect 25004 26324 25010 26336
rect 25130 26324 25136 26376
rect 25188 26364 25194 26376
rect 25240 26364 25268 26404
rect 27614 26392 27620 26404
rect 27672 26392 27678 26444
rect 27985 26435 28043 26441
rect 27985 26401 27997 26435
rect 28031 26432 28043 26435
rect 28092 26432 28120 26460
rect 28534 26432 28540 26444
rect 28031 26404 28120 26432
rect 28495 26404 28540 26432
rect 28031 26401 28043 26404
rect 27985 26395 28043 26401
rect 28534 26392 28540 26404
rect 28592 26392 28598 26444
rect 31205 26435 31263 26441
rect 31205 26401 31217 26435
rect 31251 26432 31263 26435
rect 32217 26435 32275 26441
rect 32217 26432 32229 26435
rect 31251 26404 32229 26432
rect 31251 26401 31263 26404
rect 31205 26395 31263 26401
rect 32217 26401 32229 26404
rect 32263 26432 32275 26435
rect 32398 26432 32404 26444
rect 32263 26404 32404 26432
rect 32263 26401 32275 26404
rect 32217 26395 32275 26401
rect 32398 26392 32404 26404
rect 32456 26392 32462 26444
rect 32490 26392 32496 26444
rect 32548 26432 32554 26444
rect 32548 26404 33548 26432
rect 32548 26392 32554 26404
rect 25188 26336 25281 26364
rect 25188 26324 25194 26336
rect 26326 26324 26332 26376
rect 26384 26364 26390 26376
rect 27157 26367 27215 26373
rect 27157 26366 27169 26367
rect 27080 26364 27169 26366
rect 26384 26338 27169 26364
rect 26384 26336 27108 26338
rect 26384 26324 26390 26336
rect 27157 26333 27169 26338
rect 27203 26333 27215 26367
rect 27157 26327 27215 26333
rect 28074 26324 28080 26376
rect 28132 26364 28138 26376
rect 28169 26367 28227 26373
rect 28169 26364 28181 26367
rect 28132 26336 28181 26364
rect 28132 26324 28138 26336
rect 28169 26333 28181 26336
rect 28215 26333 28227 26367
rect 28169 26327 28227 26333
rect 31849 26367 31907 26373
rect 31849 26333 31861 26367
rect 31895 26364 31907 26367
rect 32122 26364 32128 26376
rect 31895 26336 32128 26364
rect 31895 26333 31907 26336
rect 31849 26327 31907 26333
rect 32122 26324 32128 26336
rect 32180 26324 32186 26376
rect 33134 26364 33140 26376
rect 33095 26336 33140 26364
rect 33134 26324 33140 26336
rect 33192 26324 33198 26376
rect 33226 26324 33232 26376
rect 33284 26364 33290 26376
rect 33410 26364 33416 26376
rect 33284 26336 33329 26364
rect 33371 26336 33416 26364
rect 33284 26324 33290 26336
rect 33410 26324 33416 26336
rect 33468 26324 33474 26376
rect 33520 26373 33548 26404
rect 33594 26392 33600 26444
rect 33652 26432 33658 26444
rect 33652 26404 35756 26432
rect 33652 26392 33658 26404
rect 33505 26367 33563 26373
rect 33505 26333 33517 26367
rect 33551 26333 33563 26367
rect 33962 26364 33968 26376
rect 33923 26336 33968 26364
rect 33505 26327 33563 26333
rect 33962 26324 33968 26336
rect 34020 26324 34026 26376
rect 34146 26364 34152 26376
rect 34107 26336 34152 26364
rect 34146 26324 34152 26336
rect 34204 26324 34210 26376
rect 35434 26364 35440 26376
rect 35395 26336 35440 26364
rect 35434 26324 35440 26336
rect 35492 26324 35498 26376
rect 35526 26324 35532 26376
rect 35584 26364 35590 26376
rect 35728 26373 35756 26404
rect 35713 26367 35771 26373
rect 35584 26336 35629 26364
rect 35584 26324 35590 26336
rect 35713 26333 35725 26367
rect 35759 26333 35771 26367
rect 35713 26327 35771 26333
rect 35802 26324 35808 26376
rect 35860 26364 35866 26376
rect 36725 26367 36783 26373
rect 35860 26336 35905 26364
rect 35860 26324 35866 26336
rect 36725 26333 36737 26367
rect 36771 26364 36783 26367
rect 36814 26364 36820 26376
rect 36771 26336 36820 26364
rect 36771 26333 36783 26336
rect 36725 26327 36783 26333
rect 36814 26324 36820 26336
rect 36872 26324 36878 26376
rect 36992 26367 37050 26373
rect 36992 26333 37004 26367
rect 37038 26364 37050 26367
rect 37458 26364 37464 26376
rect 37038 26336 37464 26364
rect 37038 26333 37050 26336
rect 36992 26327 37050 26333
rect 37458 26324 37464 26336
rect 37516 26324 37522 26376
rect 25774 26296 25780 26308
rect 22572 26268 23520 26296
rect 24780 26268 25452 26296
rect 25735 26268 25780 26296
rect 21634 26228 21640 26240
rect 20763 26200 21496 26228
rect 21595 26200 21640 26228
rect 20763 26197 20775 26200
rect 20717 26191 20775 26197
rect 21634 26188 21640 26200
rect 21692 26188 21698 26240
rect 23492 26237 23520 26268
rect 23477 26231 23535 26237
rect 23477 26197 23489 26231
rect 23523 26228 23535 26231
rect 24026 26228 24032 26240
rect 23523 26200 24032 26228
rect 23523 26197 23535 26200
rect 23477 26191 23535 26197
rect 24026 26188 24032 26200
rect 24084 26188 24090 26240
rect 25314 26228 25320 26240
rect 25275 26200 25320 26228
rect 25314 26188 25320 26200
rect 25372 26188 25378 26240
rect 25424 26228 25452 26268
rect 25774 26256 25780 26268
rect 25832 26256 25838 26308
rect 25958 26296 25964 26308
rect 25919 26268 25964 26296
rect 25958 26256 25964 26268
rect 26016 26296 26022 26308
rect 26418 26296 26424 26308
rect 26016 26268 26424 26296
rect 26016 26256 26022 26268
rect 26418 26256 26424 26268
rect 26476 26296 26482 26308
rect 27341 26299 27399 26305
rect 27341 26296 27353 26299
rect 26476 26268 27353 26296
rect 26476 26256 26482 26268
rect 27341 26265 27353 26268
rect 27387 26265 27399 26299
rect 27341 26259 27399 26265
rect 31021 26299 31079 26305
rect 31021 26265 31033 26299
rect 31067 26296 31079 26299
rect 32953 26299 33011 26305
rect 32953 26296 32965 26299
rect 31067 26268 32965 26296
rect 31067 26265 31079 26268
rect 31021 26259 31079 26265
rect 32953 26265 32965 26268
rect 32999 26296 33011 26299
rect 37090 26296 37096 26308
rect 32999 26268 37096 26296
rect 32999 26265 33011 26268
rect 32953 26259 33011 26265
rect 37090 26256 37096 26268
rect 37148 26256 37154 26308
rect 26142 26228 26148 26240
rect 25424 26200 26148 26228
rect 26142 26188 26148 26200
rect 26200 26188 26206 26240
rect 28442 26228 28448 26240
rect 28403 26200 28448 26228
rect 28442 26188 28448 26200
rect 28500 26188 28506 26240
rect 30558 26228 30564 26240
rect 30519 26200 30564 26228
rect 30558 26188 30564 26200
rect 30616 26188 30622 26240
rect 30926 26228 30932 26240
rect 30839 26200 30932 26228
rect 30926 26188 30932 26200
rect 30984 26228 30990 26240
rect 31294 26228 31300 26240
rect 30984 26200 31300 26228
rect 30984 26188 30990 26200
rect 31294 26188 31300 26200
rect 31352 26188 31358 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 5074 25984 5080 26036
rect 5132 26024 5138 26036
rect 5445 26027 5503 26033
rect 5445 26024 5457 26027
rect 5132 25996 5457 26024
rect 5132 25984 5138 25996
rect 5445 25993 5457 25996
rect 5491 26024 5503 26027
rect 7926 26024 7932 26036
rect 5491 25996 6684 26024
rect 5491 25993 5503 25996
rect 5445 25987 5503 25993
rect 6362 25956 6368 25968
rect 5276 25928 6368 25956
rect 5276 25897 5304 25928
rect 6362 25916 6368 25928
rect 6420 25956 6426 25968
rect 6549 25959 6607 25965
rect 6549 25956 6561 25959
rect 6420 25928 6561 25956
rect 6420 25916 6426 25928
rect 6549 25925 6561 25928
rect 6595 25925 6607 25959
rect 6656 25956 6684 25996
rect 7116 25996 7932 26024
rect 6656 25928 6860 25956
rect 6549 25919 6607 25925
rect 5261 25891 5319 25897
rect 5261 25857 5273 25891
rect 5307 25857 5319 25891
rect 5261 25851 5319 25857
rect 5537 25891 5595 25897
rect 5537 25857 5549 25891
rect 5583 25857 5595 25891
rect 6730 25888 6736 25900
rect 6691 25860 6736 25888
rect 5537 25851 5595 25857
rect 4890 25780 4896 25832
rect 4948 25820 4954 25832
rect 5552 25820 5580 25851
rect 6730 25848 6736 25860
rect 6788 25848 6794 25900
rect 6832 25897 6860 25928
rect 6825 25891 6883 25897
rect 6825 25857 6837 25891
rect 6871 25888 6883 25891
rect 7116 25888 7144 25996
rect 7926 25984 7932 25996
rect 7984 26024 7990 26036
rect 8037 26027 8095 26033
rect 8037 26024 8049 26027
rect 7984 25996 8049 26024
rect 7984 25984 7990 25996
rect 8037 25993 8049 25996
rect 8083 25993 8095 26027
rect 8037 25987 8095 25993
rect 7837 25959 7895 25965
rect 7837 25925 7849 25959
rect 7883 25925 7895 25959
rect 8052 25956 8080 25987
rect 8202 25984 8208 26036
rect 8260 26024 8266 26036
rect 9858 26024 9864 26036
rect 8260 25996 9864 26024
rect 8260 25984 8266 25996
rect 9858 25984 9864 25996
rect 9916 25984 9922 26036
rect 14553 26027 14611 26033
rect 14553 25993 14565 26027
rect 14599 26024 14611 26027
rect 15102 26024 15108 26036
rect 14599 25996 15108 26024
rect 14599 25993 14611 25996
rect 14553 25987 14611 25993
rect 15102 25984 15108 25996
rect 15160 25984 15166 26036
rect 16942 25984 16948 26036
rect 17000 25984 17006 26036
rect 18138 26024 18144 26036
rect 18099 25996 18144 26024
rect 18138 25984 18144 25996
rect 18196 25984 18202 26036
rect 18432 25996 20944 26024
rect 9398 25956 9404 25968
rect 8052 25928 9404 25956
rect 7837 25919 7895 25925
rect 6871 25860 7144 25888
rect 7852 25888 7880 25919
rect 9398 25916 9404 25928
rect 9456 25916 9462 25968
rect 13170 25916 13176 25968
rect 13228 25956 13234 25968
rect 13418 25959 13476 25965
rect 13418 25956 13430 25959
rect 13228 25928 13430 25956
rect 13228 25916 13234 25928
rect 13418 25925 13430 25928
rect 13464 25925 13476 25959
rect 16960 25956 16988 25984
rect 17129 25959 17187 25965
rect 17129 25956 17141 25959
rect 16960 25928 17141 25956
rect 13418 25919 13476 25925
rect 17129 25925 17141 25928
rect 17175 25925 17187 25959
rect 17129 25919 17187 25925
rect 8478 25888 8484 25900
rect 7852 25860 8484 25888
rect 6871 25857 6883 25860
rect 6825 25851 6883 25857
rect 8478 25848 8484 25860
rect 8536 25888 8542 25900
rect 9214 25888 9220 25900
rect 8536 25860 9220 25888
rect 8536 25848 8542 25860
rect 9214 25848 9220 25860
rect 9272 25848 9278 25900
rect 9950 25848 9956 25900
rect 10008 25888 10014 25900
rect 10137 25891 10195 25897
rect 10137 25888 10149 25891
rect 10008 25860 10149 25888
rect 10008 25848 10014 25860
rect 10137 25857 10149 25860
rect 10183 25857 10195 25891
rect 10137 25851 10195 25857
rect 10321 25891 10379 25897
rect 10321 25857 10333 25891
rect 10367 25888 10379 25891
rect 10594 25888 10600 25900
rect 10367 25860 10600 25888
rect 10367 25857 10379 25860
rect 10321 25851 10379 25857
rect 10594 25848 10600 25860
rect 10652 25888 10658 25900
rect 10870 25888 10876 25900
rect 10652 25860 10876 25888
rect 10652 25848 10658 25860
rect 10870 25848 10876 25860
rect 10928 25848 10934 25900
rect 16945 25891 17003 25897
rect 16945 25857 16957 25891
rect 16991 25888 17003 25891
rect 17034 25888 17040 25900
rect 16991 25860 17040 25888
rect 16991 25857 17003 25860
rect 16945 25851 17003 25857
rect 17034 25848 17040 25860
rect 17092 25848 17098 25900
rect 17678 25848 17684 25900
rect 17736 25888 17742 25900
rect 18325 25891 18383 25897
rect 18325 25888 18337 25891
rect 17736 25860 18337 25888
rect 17736 25848 17742 25860
rect 18325 25857 18337 25860
rect 18371 25888 18383 25891
rect 18432 25888 18460 25996
rect 19978 25956 19984 25968
rect 18616 25928 19984 25956
rect 18616 25900 18644 25928
rect 19978 25916 19984 25928
rect 20036 25916 20042 25968
rect 18598 25888 18604 25900
rect 18371 25860 18460 25888
rect 18511 25860 18604 25888
rect 18371 25857 18383 25860
rect 18325 25851 18383 25857
rect 18598 25848 18604 25860
rect 18656 25848 18662 25900
rect 19429 25891 19487 25897
rect 19429 25857 19441 25891
rect 19475 25888 19487 25891
rect 20346 25888 20352 25900
rect 19475 25860 20352 25888
rect 19475 25857 19487 25860
rect 19429 25851 19487 25857
rect 20346 25848 20352 25860
rect 20404 25848 20410 25900
rect 13170 25820 13176 25832
rect 4948 25792 5580 25820
rect 13131 25792 13176 25820
rect 4948 25780 4954 25792
rect 13170 25780 13176 25792
rect 13228 25780 13234 25832
rect 19613 25823 19671 25829
rect 19613 25789 19625 25823
rect 19659 25789 19671 25823
rect 19613 25783 19671 25789
rect 19889 25823 19947 25829
rect 19889 25789 19901 25823
rect 19935 25789 19947 25823
rect 19889 25783 19947 25789
rect 19981 25823 20039 25829
rect 19981 25789 19993 25823
rect 20027 25820 20039 25823
rect 20456 25820 20484 25996
rect 20916 25956 20944 25996
rect 21634 25984 21640 26036
rect 21692 26024 21698 26036
rect 22462 26024 22468 26036
rect 21692 25996 22468 26024
rect 21692 25984 21698 25996
rect 22462 25984 22468 25996
rect 22520 26024 22526 26036
rect 22557 26027 22615 26033
rect 22557 26024 22569 26027
rect 22520 25996 22569 26024
rect 22520 25984 22526 25996
rect 22557 25993 22569 25996
rect 22603 25993 22615 26027
rect 22557 25987 22615 25993
rect 23842 25984 23848 26036
rect 23900 26024 23906 26036
rect 24489 26027 24547 26033
rect 24489 26024 24501 26027
rect 23900 25996 24501 26024
rect 23900 25984 23906 25996
rect 24489 25993 24501 25996
rect 24535 25993 24547 26027
rect 24489 25987 24547 25993
rect 24578 25984 24584 26036
rect 24636 26024 24642 26036
rect 32122 26024 32128 26036
rect 24636 25996 32128 26024
rect 24636 25984 24642 25996
rect 32122 25984 32128 25996
rect 32180 25984 32186 26036
rect 32858 25984 32864 26036
rect 32916 26024 32922 26036
rect 33321 26027 33379 26033
rect 33321 26024 33333 26027
rect 32916 25996 33333 26024
rect 32916 25984 32922 25996
rect 33321 25993 33333 25996
rect 33367 25993 33379 26027
rect 33321 25987 33379 25993
rect 23014 25956 23020 25968
rect 20916 25928 23020 25956
rect 23014 25916 23020 25928
rect 23072 25916 23078 25968
rect 23124 25928 24716 25956
rect 20625 25891 20683 25897
rect 20625 25857 20637 25891
rect 20671 25857 20683 25891
rect 20625 25851 20683 25857
rect 20027 25792 20484 25820
rect 20640 25820 20668 25851
rect 20714 25848 20720 25900
rect 20772 25888 20778 25900
rect 20809 25891 20867 25897
rect 20809 25888 20821 25891
rect 20772 25860 20821 25888
rect 20772 25848 20778 25860
rect 20809 25857 20821 25860
rect 20855 25857 20867 25891
rect 20809 25851 20867 25857
rect 20898 25848 20904 25900
rect 20956 25888 20962 25900
rect 21177 25891 21235 25897
rect 21177 25888 21189 25891
rect 20956 25860 21189 25888
rect 20956 25848 20962 25860
rect 21177 25857 21189 25860
rect 21223 25888 21235 25891
rect 21450 25888 21456 25900
rect 21223 25860 21456 25888
rect 21223 25857 21235 25860
rect 21177 25851 21235 25857
rect 21450 25848 21456 25860
rect 21508 25848 21514 25900
rect 23124 25897 23152 25928
rect 24504 25900 24532 25928
rect 23109 25891 23167 25897
rect 23109 25857 23121 25891
rect 23155 25857 23167 25891
rect 23566 25888 23572 25900
rect 23109 25851 23167 25857
rect 23400 25860 23572 25888
rect 20990 25820 20996 25832
rect 20640 25792 20996 25820
rect 20027 25789 20039 25792
rect 19981 25783 20039 25789
rect 4430 25712 4436 25764
rect 4488 25752 4494 25764
rect 5077 25755 5135 25761
rect 5077 25752 5089 25755
rect 4488 25724 5089 25752
rect 4488 25712 4494 25724
rect 5077 25721 5089 25724
rect 5123 25752 5135 25755
rect 7466 25752 7472 25764
rect 5123 25724 7472 25752
rect 5123 25721 5135 25724
rect 5077 25715 5135 25721
rect 7466 25712 7472 25724
rect 7524 25712 7530 25764
rect 19334 25712 19340 25764
rect 19392 25752 19398 25764
rect 19628 25752 19656 25783
rect 19392 25724 19656 25752
rect 19904 25752 19932 25783
rect 20990 25780 20996 25792
rect 21048 25820 21054 25832
rect 23400 25820 23428 25860
rect 23566 25848 23572 25860
rect 23624 25848 23630 25900
rect 23661 25891 23719 25897
rect 23661 25857 23673 25891
rect 23707 25857 23719 25891
rect 23661 25851 23719 25857
rect 21048 25792 23428 25820
rect 23676 25820 23704 25851
rect 24486 25848 24492 25900
rect 24544 25848 24550 25900
rect 24688 25897 24716 25928
rect 25038 25916 25044 25968
rect 25096 25956 25102 25968
rect 30745 25959 30803 25965
rect 30745 25956 30757 25959
rect 25096 25928 30757 25956
rect 25096 25916 25102 25928
rect 30745 25925 30757 25928
rect 30791 25956 30803 25959
rect 31018 25956 31024 25968
rect 30791 25928 31024 25956
rect 30791 25925 30803 25928
rect 30745 25919 30803 25925
rect 31018 25916 31024 25928
rect 31076 25956 31082 25968
rect 35342 25956 35348 25968
rect 31076 25928 35348 25956
rect 31076 25916 31082 25928
rect 35342 25916 35348 25928
rect 35400 25916 35406 25968
rect 24673 25891 24731 25897
rect 24673 25857 24685 25891
rect 24719 25857 24731 25891
rect 24673 25851 24731 25857
rect 24949 25891 25007 25897
rect 24949 25857 24961 25891
rect 24995 25878 25007 25891
rect 25133 25891 25191 25897
rect 24995 25857 25084 25878
rect 24949 25851 25084 25857
rect 25133 25857 25145 25891
rect 25179 25888 25191 25891
rect 26142 25888 26148 25900
rect 25179 25860 26148 25888
rect 25179 25857 25191 25860
rect 25133 25851 25191 25857
rect 24964 25850 25084 25851
rect 25056 25820 25084 25850
rect 26142 25848 26148 25860
rect 26200 25848 26206 25900
rect 27522 25888 27528 25900
rect 27483 25860 27528 25888
rect 27522 25848 27528 25860
rect 27580 25848 27586 25900
rect 27709 25891 27767 25897
rect 27709 25857 27721 25891
rect 27755 25857 27767 25891
rect 27709 25851 27767 25857
rect 27801 25891 27859 25897
rect 27801 25857 27813 25891
rect 27847 25857 27859 25891
rect 27801 25851 27859 25857
rect 27893 25891 27951 25897
rect 27893 25857 27905 25891
rect 27939 25888 27951 25891
rect 27939 25860 28212 25888
rect 27939 25857 27951 25860
rect 27893 25851 27951 25857
rect 25406 25820 25412 25832
rect 23676 25792 24624 25820
rect 25056 25792 25412 25820
rect 21048 25780 21054 25792
rect 20070 25752 20076 25764
rect 19904 25724 20076 25752
rect 19392 25712 19398 25724
rect 20070 25712 20076 25724
rect 20128 25752 20134 25764
rect 20438 25752 20444 25764
rect 20128 25724 20444 25752
rect 20128 25712 20134 25724
rect 20438 25712 20444 25724
rect 20496 25712 20502 25764
rect 20622 25712 20628 25764
rect 20680 25752 20686 25764
rect 23676 25752 23704 25792
rect 24596 25764 24624 25792
rect 25406 25780 25412 25792
rect 25464 25780 25470 25832
rect 26694 25780 26700 25832
rect 26752 25820 26758 25832
rect 27154 25820 27160 25832
rect 26752 25792 27160 25820
rect 26752 25780 26758 25792
rect 27154 25780 27160 25792
rect 27212 25820 27218 25832
rect 27724 25820 27752 25851
rect 27212 25792 27752 25820
rect 27816 25820 27844 25851
rect 27982 25820 27988 25832
rect 27816 25792 27988 25820
rect 27212 25780 27218 25792
rect 27982 25780 27988 25792
rect 28040 25780 28046 25832
rect 28184 25820 28212 25860
rect 28442 25848 28448 25900
rect 28500 25888 28506 25900
rect 28537 25891 28595 25897
rect 28537 25888 28549 25891
rect 28500 25860 28549 25888
rect 28500 25848 28506 25860
rect 28537 25857 28549 25860
rect 28583 25857 28595 25891
rect 33134 25888 33140 25900
rect 33047 25860 33140 25888
rect 28537 25851 28595 25857
rect 33134 25848 33140 25860
rect 33192 25888 33198 25900
rect 34146 25888 34152 25900
rect 33192 25860 34152 25888
rect 33192 25848 33198 25860
rect 34146 25848 34152 25860
rect 34204 25848 34210 25900
rect 37829 25891 37887 25897
rect 37829 25857 37841 25891
rect 37875 25888 37887 25891
rect 37918 25888 37924 25900
rect 37875 25860 37924 25888
rect 37875 25857 37887 25860
rect 37829 25851 37887 25857
rect 37918 25848 37924 25860
rect 37976 25848 37982 25900
rect 28350 25820 28356 25832
rect 28184 25792 28356 25820
rect 20680 25724 23704 25752
rect 20680 25712 20686 25724
rect 24578 25712 24584 25764
rect 24636 25752 24642 25764
rect 24765 25755 24823 25761
rect 24765 25752 24777 25755
rect 24636 25724 24777 25752
rect 24636 25712 24642 25724
rect 24765 25721 24777 25724
rect 24811 25721 24823 25755
rect 24765 25715 24823 25721
rect 24854 25712 24860 25764
rect 24912 25752 24918 25764
rect 24912 25724 24957 25752
rect 24912 25712 24918 25724
rect 26234 25712 26240 25764
rect 26292 25752 26298 25764
rect 28184 25752 28212 25792
rect 28350 25780 28356 25792
rect 28408 25820 28414 25832
rect 28810 25820 28816 25832
rect 28408 25792 28816 25820
rect 28408 25780 28414 25792
rect 28810 25780 28816 25792
rect 28868 25780 28874 25832
rect 28994 25820 29000 25832
rect 28955 25792 29000 25820
rect 28994 25780 29000 25792
rect 29052 25780 29058 25832
rect 31573 25823 31631 25829
rect 31573 25789 31585 25823
rect 31619 25820 31631 25823
rect 31754 25820 31760 25832
rect 31619 25792 31760 25820
rect 31619 25789 31631 25792
rect 31573 25783 31631 25789
rect 31754 25780 31760 25792
rect 31812 25820 31818 25832
rect 32674 25820 32680 25832
rect 31812 25792 32680 25820
rect 31812 25780 31818 25792
rect 32674 25780 32680 25792
rect 32732 25780 32738 25832
rect 32953 25823 33011 25829
rect 32953 25789 32965 25823
rect 32999 25820 33011 25823
rect 33962 25820 33968 25832
rect 32999 25792 33968 25820
rect 32999 25789 33011 25792
rect 32953 25783 33011 25789
rect 33962 25780 33968 25792
rect 34020 25780 34026 25832
rect 38102 25820 38108 25832
rect 38063 25792 38108 25820
rect 38102 25780 38108 25792
rect 38160 25780 38166 25832
rect 26292 25724 28212 25752
rect 26292 25712 26298 25724
rect 4801 25687 4859 25693
rect 4801 25653 4813 25687
rect 4847 25684 4859 25687
rect 4890 25684 4896 25696
rect 4847 25656 4896 25684
rect 4847 25653 4859 25656
rect 4801 25647 4859 25653
rect 4890 25644 4896 25656
rect 4948 25644 4954 25696
rect 5166 25684 5172 25696
rect 5127 25656 5172 25684
rect 5166 25644 5172 25656
rect 5224 25644 5230 25696
rect 6454 25644 6460 25696
rect 6512 25684 6518 25696
rect 6549 25687 6607 25693
rect 6549 25684 6561 25687
rect 6512 25656 6561 25684
rect 6512 25644 6518 25656
rect 6549 25653 6561 25656
rect 6595 25653 6607 25687
rect 6549 25647 6607 25653
rect 8021 25687 8079 25693
rect 8021 25653 8033 25687
rect 8067 25684 8079 25687
rect 8110 25684 8116 25696
rect 8067 25656 8116 25684
rect 8067 25653 8079 25656
rect 8021 25647 8079 25653
rect 8110 25644 8116 25656
rect 8168 25684 8174 25696
rect 9306 25684 9312 25696
rect 8168 25656 9312 25684
rect 8168 25644 8174 25656
rect 9306 25644 9312 25656
rect 9364 25644 9370 25696
rect 10137 25687 10195 25693
rect 10137 25653 10149 25687
rect 10183 25684 10195 25687
rect 10594 25684 10600 25696
rect 10183 25656 10600 25684
rect 10183 25653 10195 25656
rect 10137 25647 10195 25653
rect 10594 25644 10600 25656
rect 10652 25644 10658 25696
rect 17218 25684 17224 25696
rect 17179 25656 17224 25684
rect 17218 25644 17224 25656
rect 17276 25644 17282 25696
rect 28077 25687 28135 25693
rect 28077 25653 28089 25687
rect 28123 25684 28135 25687
rect 28166 25684 28172 25696
rect 28123 25656 28172 25684
rect 28123 25653 28135 25656
rect 28077 25647 28135 25653
rect 28166 25644 28172 25656
rect 28224 25644 28230 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 5626 25440 5632 25492
rect 5684 25480 5690 25492
rect 6273 25483 6331 25489
rect 6273 25480 6285 25483
rect 5684 25452 6285 25480
rect 5684 25440 5690 25452
rect 6273 25449 6285 25452
rect 6319 25449 6331 25483
rect 6273 25443 6331 25449
rect 8386 25440 8392 25492
rect 8444 25480 8450 25492
rect 9309 25483 9367 25489
rect 9309 25480 9321 25483
rect 8444 25452 9321 25480
rect 8444 25440 8450 25452
rect 9309 25449 9321 25452
rect 9355 25480 9367 25483
rect 10318 25480 10324 25492
rect 9355 25452 10324 25480
rect 9355 25449 9367 25452
rect 9309 25443 9367 25449
rect 10318 25440 10324 25452
rect 10376 25440 10382 25492
rect 12897 25483 12955 25489
rect 12897 25480 12909 25483
rect 10796 25452 12909 25480
rect 5166 25372 5172 25424
rect 5224 25412 5230 25424
rect 7929 25415 7987 25421
rect 7929 25412 7941 25415
rect 5224 25384 7941 25412
rect 5224 25372 5230 25384
rect 7929 25381 7941 25384
rect 7975 25412 7987 25415
rect 8018 25412 8024 25424
rect 7975 25384 8024 25412
rect 7975 25381 7987 25384
rect 7929 25375 7987 25381
rect 8018 25372 8024 25384
rect 8076 25372 8082 25424
rect 4341 25347 4399 25353
rect 4341 25313 4353 25347
rect 4387 25344 4399 25347
rect 4706 25344 4712 25356
rect 4387 25316 4712 25344
rect 4387 25313 4399 25316
rect 4341 25307 4399 25313
rect 4706 25304 4712 25316
rect 4764 25304 4770 25356
rect 4890 25344 4896 25356
rect 4851 25316 4896 25344
rect 4890 25304 4896 25316
rect 4948 25304 4954 25356
rect 5261 25347 5319 25353
rect 5261 25313 5273 25347
rect 5307 25344 5319 25347
rect 5442 25344 5448 25356
rect 5307 25316 5448 25344
rect 5307 25313 5319 25316
rect 5261 25307 5319 25313
rect 5442 25304 5448 25316
rect 5500 25304 5506 25356
rect 6454 25344 6460 25356
rect 6415 25316 6460 25344
rect 6454 25304 6460 25316
rect 6512 25304 6518 25356
rect 6549 25347 6607 25353
rect 6549 25313 6561 25347
rect 6595 25344 6607 25347
rect 6914 25344 6920 25356
rect 6595 25316 6920 25344
rect 6595 25313 6607 25316
rect 6549 25307 6607 25313
rect 6914 25304 6920 25316
rect 6972 25304 6978 25356
rect 9674 25344 9680 25356
rect 8036 25316 9680 25344
rect 4154 25276 4160 25288
rect 4115 25248 4160 25276
rect 4154 25236 4160 25248
rect 4212 25236 4218 25288
rect 4430 25236 4436 25288
rect 4488 25276 4494 25288
rect 5350 25276 5356 25288
rect 4488 25248 4533 25276
rect 5311 25248 5356 25276
rect 4488 25236 4494 25248
rect 5350 25236 5356 25248
rect 5408 25236 5414 25288
rect 5460 25276 5488 25304
rect 6641 25279 6699 25285
rect 6641 25276 6653 25279
rect 5460 25248 6653 25276
rect 6641 25245 6653 25248
rect 6687 25245 6699 25279
rect 6641 25239 6699 25245
rect 6733 25279 6791 25285
rect 6733 25245 6745 25279
rect 6779 25276 6791 25279
rect 8036 25276 8064 25316
rect 9674 25304 9680 25316
rect 9732 25304 9738 25356
rect 6779 25248 8064 25276
rect 6779 25245 6791 25248
rect 6733 25239 6791 25245
rect 8110 25236 8116 25288
rect 8168 25276 8174 25288
rect 8386 25276 8392 25288
rect 8168 25248 8213 25276
rect 8347 25248 8392 25276
rect 8168 25236 8174 25248
rect 8386 25236 8392 25248
rect 8444 25236 8450 25288
rect 10505 25279 10563 25285
rect 10505 25276 10517 25279
rect 9508 25248 10517 25276
rect 9125 25211 9183 25217
rect 9125 25208 9137 25211
rect 8588 25180 9137 25208
rect 3970 25140 3976 25152
rect 3931 25112 3976 25140
rect 3970 25100 3976 25112
rect 4028 25100 4034 25152
rect 5534 25140 5540 25152
rect 5495 25112 5540 25140
rect 5534 25100 5540 25112
rect 5592 25100 5598 25152
rect 7466 25100 7472 25152
rect 7524 25140 7530 25152
rect 8588 25140 8616 25180
rect 9125 25177 9137 25180
rect 9171 25177 9183 25211
rect 9125 25171 9183 25177
rect 9508 25152 9536 25248
rect 10505 25245 10517 25248
rect 10551 25245 10563 25279
rect 10505 25239 10563 25245
rect 10594 25236 10600 25288
rect 10652 25276 10658 25288
rect 10796 25285 10824 25452
rect 12897 25449 12909 25452
rect 12943 25480 12955 25483
rect 19150 25480 19156 25492
rect 12943 25452 19156 25480
rect 12943 25449 12955 25452
rect 12897 25443 12955 25449
rect 19150 25440 19156 25452
rect 19208 25440 19214 25492
rect 21358 25440 21364 25492
rect 21416 25480 21422 25492
rect 21913 25483 21971 25489
rect 21913 25480 21925 25483
rect 21416 25452 21925 25480
rect 21416 25440 21422 25452
rect 21913 25449 21925 25452
rect 21959 25480 21971 25483
rect 26234 25480 26240 25492
rect 21959 25452 26240 25480
rect 21959 25449 21971 25452
rect 21913 25443 21971 25449
rect 26234 25440 26240 25452
rect 26292 25440 26298 25492
rect 27617 25483 27675 25489
rect 27617 25449 27629 25483
rect 27663 25480 27675 25483
rect 28074 25480 28080 25492
rect 27663 25452 28080 25480
rect 27663 25449 27675 25452
rect 27617 25443 27675 25449
rect 28074 25440 28080 25452
rect 28132 25440 28138 25492
rect 29914 25480 29920 25492
rect 28553 25452 29920 25480
rect 16574 25412 16580 25424
rect 16535 25384 16580 25412
rect 16574 25372 16580 25384
rect 16632 25372 16638 25424
rect 18506 25412 18512 25424
rect 16684 25384 18512 25412
rect 13722 25304 13728 25356
rect 13780 25344 13786 25356
rect 13780 25316 14320 25344
rect 13780 25304 13786 25316
rect 10689 25279 10747 25285
rect 10689 25276 10701 25279
rect 10652 25248 10701 25276
rect 10652 25236 10658 25248
rect 10689 25245 10701 25248
rect 10735 25245 10747 25279
rect 10689 25239 10747 25245
rect 10781 25279 10839 25285
rect 10781 25245 10793 25279
rect 10827 25245 10839 25279
rect 10781 25239 10839 25245
rect 10870 25236 10876 25288
rect 10928 25276 10934 25288
rect 11517 25279 11575 25285
rect 10928 25248 10973 25276
rect 10928 25236 10934 25248
rect 11517 25245 11529 25279
rect 11563 25276 11575 25279
rect 13170 25276 13176 25288
rect 11563 25248 13176 25276
rect 11563 25245 11575 25248
rect 11517 25239 11575 25245
rect 13170 25236 13176 25248
rect 13228 25276 13234 25288
rect 14182 25276 14188 25288
rect 13228 25248 14188 25276
rect 13228 25236 13234 25248
rect 14182 25236 14188 25248
rect 14240 25236 14246 25288
rect 14292 25285 14320 25316
rect 14277 25279 14335 25285
rect 14277 25245 14289 25279
rect 14323 25245 14335 25279
rect 14642 25276 14648 25288
rect 14603 25248 14648 25276
rect 14277 25239 14335 25245
rect 14642 25236 14648 25248
rect 14700 25236 14706 25288
rect 11762 25211 11820 25217
rect 11762 25208 11774 25211
rect 11072 25180 11774 25208
rect 7524 25112 8616 25140
rect 7524 25100 7530 25112
rect 9214 25100 9220 25152
rect 9272 25140 9278 25152
rect 9309 25143 9367 25149
rect 9309 25140 9321 25143
rect 9272 25112 9321 25140
rect 9272 25100 9278 25112
rect 9309 25109 9321 25112
rect 9355 25109 9367 25143
rect 9490 25140 9496 25152
rect 9451 25112 9496 25140
rect 9309 25103 9367 25109
rect 9490 25100 9496 25112
rect 9548 25100 9554 25152
rect 11072 25149 11100 25180
rect 11762 25177 11774 25180
rect 11808 25177 11820 25211
rect 11762 25171 11820 25177
rect 13538 25168 13544 25220
rect 13596 25208 13602 25220
rect 14461 25211 14519 25217
rect 14461 25208 14473 25211
rect 13596 25180 14473 25208
rect 13596 25168 13602 25180
rect 14461 25177 14473 25180
rect 14507 25177 14519 25211
rect 14461 25171 14519 25177
rect 14553 25211 14611 25217
rect 14553 25177 14565 25211
rect 14599 25208 14611 25211
rect 15654 25208 15660 25220
rect 14599 25180 15660 25208
rect 14599 25177 14611 25180
rect 14553 25171 14611 25177
rect 15654 25168 15660 25180
rect 15712 25168 15718 25220
rect 11057 25143 11115 25149
rect 11057 25109 11069 25143
rect 11103 25109 11115 25143
rect 14826 25140 14832 25152
rect 14787 25112 14832 25140
rect 11057 25103 11115 25109
rect 14826 25100 14832 25112
rect 14884 25100 14890 25152
rect 16684 25140 16712 25384
rect 18506 25372 18512 25384
rect 18564 25372 18570 25424
rect 18782 25372 18788 25424
rect 18840 25412 18846 25424
rect 19242 25412 19248 25424
rect 18840 25384 19248 25412
rect 18840 25372 18846 25384
rect 19242 25372 19248 25384
rect 19300 25412 19306 25424
rect 24762 25412 24768 25424
rect 19300 25384 24768 25412
rect 19300 25372 19306 25384
rect 18322 25344 18328 25356
rect 18283 25316 18328 25344
rect 18322 25304 18328 25316
rect 18380 25344 18386 25356
rect 18380 25316 19656 25344
rect 18380 25304 18386 25316
rect 16761 25279 16819 25285
rect 16761 25245 16773 25279
rect 16807 25276 16819 25279
rect 17678 25276 17684 25288
rect 16807 25248 17684 25276
rect 16807 25245 16819 25248
rect 16761 25239 16819 25245
rect 17678 25236 17684 25248
rect 17736 25236 17742 25288
rect 18509 25279 18567 25285
rect 18509 25245 18521 25279
rect 18555 25276 18567 25279
rect 18598 25276 18604 25288
rect 18555 25248 18604 25276
rect 18555 25245 18567 25248
rect 18509 25239 18567 25245
rect 18598 25236 18604 25248
rect 18656 25236 18662 25288
rect 18874 25276 18880 25288
rect 18835 25248 18880 25276
rect 18874 25236 18880 25248
rect 18932 25236 18938 25288
rect 19426 25236 19432 25288
rect 19484 25276 19490 25288
rect 19628 25285 19656 25316
rect 19521 25279 19579 25285
rect 19521 25276 19533 25279
rect 19484 25248 19533 25276
rect 19484 25236 19490 25248
rect 19521 25245 19533 25248
rect 19567 25245 19579 25279
rect 19521 25239 19579 25245
rect 19613 25279 19671 25285
rect 19613 25245 19625 25279
rect 19659 25245 19671 25279
rect 19613 25239 19671 25245
rect 20625 25279 20683 25285
rect 20625 25245 20637 25279
rect 20671 25245 20683 25279
rect 20990 25276 20996 25288
rect 20951 25248 20996 25276
rect 20625 25239 20683 25245
rect 16853 25211 16911 25217
rect 16853 25177 16865 25211
rect 16899 25208 16911 25211
rect 17862 25208 17868 25220
rect 16899 25180 17868 25208
rect 16899 25177 16911 25180
rect 16853 25171 16911 25177
rect 17862 25168 17868 25180
rect 17920 25168 17926 25220
rect 19536 25208 19564 25239
rect 20640 25208 20668 25239
rect 20990 25236 20996 25248
rect 21048 25236 21054 25288
rect 21634 25276 21640 25288
rect 21595 25248 21640 25276
rect 21634 25236 21640 25248
rect 21692 25236 21698 25288
rect 21818 25276 21824 25288
rect 21779 25248 21824 25276
rect 21818 25236 21824 25248
rect 21876 25236 21882 25288
rect 22940 25285 22968 25384
rect 24762 25372 24768 25384
rect 24820 25372 24826 25424
rect 24854 25372 24860 25424
rect 24912 25412 24918 25424
rect 26053 25415 26111 25421
rect 26053 25412 26065 25415
rect 24912 25384 26065 25412
rect 24912 25372 24918 25384
rect 26053 25381 26065 25384
rect 26099 25412 26111 25415
rect 28553 25412 28581 25452
rect 29914 25440 29920 25452
rect 29972 25440 29978 25492
rect 26099 25384 28581 25412
rect 28629 25415 28687 25421
rect 26099 25381 26111 25384
rect 26053 25375 26111 25381
rect 28629 25381 28641 25415
rect 28675 25412 28687 25415
rect 28902 25412 28908 25424
rect 28675 25384 28908 25412
rect 28675 25381 28687 25384
rect 28629 25375 28687 25381
rect 28902 25372 28908 25384
rect 28960 25372 28966 25424
rect 32861 25415 32919 25421
rect 32861 25381 32873 25415
rect 32907 25412 32919 25415
rect 33134 25412 33140 25424
rect 32907 25384 33140 25412
rect 32907 25381 32919 25384
rect 32861 25375 32919 25381
rect 33134 25372 33140 25384
rect 33192 25372 33198 25424
rect 25406 25304 25412 25356
rect 25464 25344 25470 25356
rect 25501 25347 25559 25353
rect 25501 25344 25513 25347
rect 25464 25316 25513 25344
rect 25464 25304 25470 25316
rect 25501 25313 25513 25316
rect 25547 25344 25559 25347
rect 25682 25344 25688 25356
rect 25547 25316 25688 25344
rect 25547 25313 25559 25316
rect 25501 25307 25559 25313
rect 25682 25304 25688 25316
rect 25740 25304 25746 25356
rect 25866 25304 25872 25356
rect 25924 25344 25930 25356
rect 30009 25347 30067 25353
rect 30009 25344 30021 25347
rect 25924 25316 30021 25344
rect 25924 25304 25930 25316
rect 30009 25313 30021 25316
rect 30055 25313 30067 25347
rect 33870 25344 33876 25356
rect 30009 25307 30067 25313
rect 32784 25316 33876 25344
rect 22741 25279 22799 25285
rect 22741 25245 22753 25279
rect 22787 25245 22799 25279
rect 22741 25239 22799 25245
rect 22925 25279 22983 25285
rect 22925 25245 22937 25279
rect 22971 25245 22983 25279
rect 24946 25276 24952 25288
rect 24907 25248 24952 25276
rect 22925 25239 22983 25245
rect 20714 25208 20720 25220
rect 19536 25180 20720 25208
rect 20714 25168 20720 25180
rect 20772 25208 20778 25220
rect 22756 25208 22784 25239
rect 24946 25236 24952 25248
rect 25004 25236 25010 25288
rect 25133 25279 25191 25285
rect 25133 25245 25145 25279
rect 25179 25276 25191 25279
rect 25222 25276 25228 25288
rect 25179 25248 25228 25276
rect 25179 25245 25191 25248
rect 25133 25239 25191 25245
rect 25222 25236 25228 25248
rect 25280 25276 25286 25288
rect 25961 25279 26019 25285
rect 25961 25276 25973 25279
rect 25280 25248 25973 25276
rect 25280 25236 25286 25248
rect 25961 25245 25973 25248
rect 26007 25245 26019 25279
rect 25961 25239 26019 25245
rect 26142 25236 26148 25288
rect 26200 25276 26206 25288
rect 26326 25276 26332 25288
rect 26200 25248 26332 25276
rect 26200 25236 26206 25248
rect 26326 25236 26332 25248
rect 26384 25276 26390 25288
rect 26513 25279 26571 25285
rect 26513 25276 26525 25279
rect 26384 25248 26525 25276
rect 26384 25236 26390 25248
rect 26513 25245 26525 25248
rect 26559 25245 26571 25279
rect 26513 25239 26571 25245
rect 26789 25279 26847 25285
rect 26789 25245 26801 25279
rect 26835 25245 26847 25279
rect 26789 25239 26847 25245
rect 20772 25180 22784 25208
rect 24964 25208 24992 25236
rect 25498 25208 25504 25220
rect 24964 25180 25504 25208
rect 20772 25168 20778 25180
rect 25498 25168 25504 25180
rect 25556 25168 25562 25220
rect 26050 25168 26056 25220
rect 26108 25208 26114 25220
rect 26804 25208 26832 25239
rect 26878 25236 26884 25288
rect 26936 25276 26942 25288
rect 27525 25279 27583 25285
rect 27525 25276 27537 25279
rect 26936 25248 27537 25276
rect 26936 25236 26942 25248
rect 27525 25245 27537 25248
rect 27571 25245 27583 25279
rect 28442 25276 28448 25288
rect 28403 25248 28448 25276
rect 27525 25239 27583 25245
rect 28442 25236 28448 25248
rect 28500 25236 28506 25288
rect 28537 25279 28595 25285
rect 28537 25245 28549 25279
rect 28583 25276 28595 25279
rect 28626 25276 28632 25288
rect 28583 25248 28632 25276
rect 28583 25245 28595 25248
rect 28537 25239 28595 25245
rect 28626 25236 28632 25248
rect 28684 25236 28690 25288
rect 28721 25279 28779 25285
rect 28721 25245 28733 25279
rect 28767 25276 28779 25279
rect 28994 25276 29000 25288
rect 28767 25248 29000 25276
rect 28767 25245 28779 25248
rect 28721 25239 28779 25245
rect 28994 25236 29000 25248
rect 29052 25236 29058 25288
rect 30024 25276 30052 25307
rect 32784 25288 32812 25316
rect 33870 25304 33876 25316
rect 33928 25304 33934 25356
rect 34054 25344 34060 25356
rect 34015 25316 34060 25344
rect 34054 25304 34060 25316
rect 34112 25304 34118 25356
rect 34333 25347 34391 25353
rect 34333 25313 34345 25347
rect 34379 25313 34391 25347
rect 34333 25307 34391 25313
rect 31754 25276 31760 25288
rect 30024 25248 31760 25276
rect 31754 25236 31760 25248
rect 31812 25236 31818 25288
rect 32401 25279 32459 25285
rect 32401 25245 32413 25279
rect 32447 25245 32459 25279
rect 32401 25239 32459 25245
rect 32585 25279 32643 25285
rect 32585 25245 32597 25279
rect 32631 25276 32643 25279
rect 32766 25276 32772 25288
rect 32631 25248 32772 25276
rect 32631 25245 32643 25248
rect 32585 25239 32643 25245
rect 26108 25180 26832 25208
rect 26108 25168 26114 25180
rect 27706 25168 27712 25220
rect 27764 25208 27770 25220
rect 29638 25208 29644 25220
rect 27764 25180 29644 25208
rect 27764 25168 27770 25180
rect 29638 25168 29644 25180
rect 29696 25168 29702 25220
rect 30276 25211 30334 25217
rect 30276 25177 30288 25211
rect 30322 25208 30334 25211
rect 30558 25208 30564 25220
rect 30322 25180 30564 25208
rect 30322 25177 30334 25180
rect 30276 25171 30334 25177
rect 30558 25168 30564 25180
rect 30616 25168 30622 25220
rect 16945 25143 17003 25149
rect 16945 25140 16957 25143
rect 16684 25112 16957 25140
rect 16945 25109 16957 25112
rect 16991 25109 17003 25143
rect 16945 25103 17003 25109
rect 17129 25143 17187 25149
rect 17129 25109 17141 25143
rect 17175 25140 17187 25143
rect 17310 25140 17316 25152
rect 17175 25112 17316 25140
rect 17175 25109 17187 25112
rect 17129 25103 17187 25109
rect 17310 25100 17316 25112
rect 17368 25100 17374 25152
rect 17770 25100 17776 25152
rect 17828 25140 17834 25152
rect 18785 25143 18843 25149
rect 18785 25140 18797 25143
rect 17828 25112 18797 25140
rect 17828 25100 17834 25112
rect 18785 25109 18797 25112
rect 18831 25140 18843 25143
rect 18966 25140 18972 25152
rect 18831 25112 18972 25140
rect 18831 25109 18843 25112
rect 18785 25103 18843 25109
rect 18966 25100 18972 25112
rect 19024 25100 19030 25152
rect 19426 25100 19432 25152
rect 19484 25140 19490 25152
rect 19521 25143 19579 25149
rect 19521 25140 19533 25143
rect 19484 25112 19533 25140
rect 19484 25100 19490 25112
rect 19521 25109 19533 25112
rect 19567 25109 19579 25143
rect 20530 25140 20536 25152
rect 20491 25112 20536 25140
rect 19521 25103 19579 25109
rect 20530 25100 20536 25112
rect 20588 25100 20594 25152
rect 23014 25140 23020 25152
rect 22975 25112 23020 25140
rect 23014 25100 23020 25112
rect 23072 25100 23078 25152
rect 24578 25100 24584 25152
rect 24636 25140 24642 25152
rect 26068 25140 26096 25168
rect 28258 25140 28264 25152
rect 24636 25112 26096 25140
rect 28219 25112 28264 25140
rect 24636 25100 24642 25112
rect 28258 25100 28264 25112
rect 28316 25100 28322 25152
rect 31294 25100 31300 25152
rect 31352 25140 31358 25152
rect 31389 25143 31447 25149
rect 31389 25140 31401 25143
rect 31352 25112 31401 25140
rect 31352 25100 31358 25112
rect 31389 25109 31401 25112
rect 31435 25109 31447 25143
rect 32416 25140 32444 25239
rect 32766 25236 32772 25248
rect 32824 25236 32830 25288
rect 32950 25276 32956 25288
rect 32911 25248 32956 25276
rect 32950 25236 32956 25248
rect 33008 25236 33014 25288
rect 33686 25236 33692 25288
rect 33744 25276 33750 25288
rect 33965 25279 34023 25285
rect 33965 25276 33977 25279
rect 33744 25248 33977 25276
rect 33744 25236 33750 25248
rect 33965 25245 33977 25248
rect 34011 25245 34023 25279
rect 33965 25239 34023 25245
rect 34348 25208 34376 25307
rect 34885 25279 34943 25285
rect 34885 25245 34897 25279
rect 34931 25276 34943 25279
rect 36814 25276 36820 25288
rect 34931 25248 36820 25276
rect 34931 25245 34943 25248
rect 34885 25239 34943 25245
rect 36814 25236 36820 25248
rect 36872 25236 36878 25288
rect 35130 25211 35188 25217
rect 35130 25208 35142 25211
rect 34348 25180 35142 25208
rect 35130 25177 35142 25180
rect 35176 25177 35188 25211
rect 35130 25171 35188 25177
rect 37084 25211 37142 25217
rect 37084 25177 37096 25211
rect 37130 25208 37142 25211
rect 37458 25208 37464 25220
rect 37130 25180 37464 25208
rect 37130 25177 37142 25180
rect 37084 25171 37142 25177
rect 37458 25168 37464 25180
rect 37516 25168 37522 25220
rect 32490 25140 32496 25152
rect 32403 25112 32496 25140
rect 31389 25103 31447 25109
rect 32490 25100 32496 25112
rect 32548 25140 32554 25152
rect 34606 25140 34612 25152
rect 32548 25112 34612 25140
rect 32548 25100 32554 25112
rect 34606 25100 34612 25112
rect 34664 25100 34670 25152
rect 36262 25140 36268 25152
rect 36223 25112 36268 25140
rect 36262 25100 36268 25112
rect 36320 25100 36326 25152
rect 37826 25100 37832 25152
rect 37884 25140 37890 25152
rect 38197 25143 38255 25149
rect 38197 25140 38209 25143
rect 37884 25112 38209 25140
rect 37884 25100 37890 25112
rect 38197 25109 38209 25112
rect 38243 25109 38255 25143
rect 38197 25103 38255 25109
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 4154 24896 4160 24948
rect 4212 24936 4218 24948
rect 4709 24939 4767 24945
rect 4709 24936 4721 24939
rect 4212 24908 4721 24936
rect 4212 24896 4218 24908
rect 4709 24905 4721 24908
rect 4755 24905 4767 24939
rect 4709 24899 4767 24905
rect 5442 24896 5448 24948
rect 5500 24936 5506 24948
rect 5905 24939 5963 24945
rect 5905 24936 5917 24939
rect 5500 24908 5917 24936
rect 5500 24896 5506 24908
rect 5905 24905 5917 24908
rect 5951 24905 5963 24939
rect 5905 24899 5963 24905
rect 8386 24896 8392 24948
rect 8444 24936 8450 24948
rect 8444 24908 9904 24936
rect 8444 24896 8450 24908
rect 2952 24871 3010 24877
rect 2952 24837 2964 24871
rect 2998 24868 3010 24871
rect 3970 24868 3976 24880
rect 2998 24840 3976 24868
rect 2998 24837 3010 24840
rect 2952 24831 3010 24837
rect 3970 24828 3976 24840
rect 4028 24828 4034 24880
rect 5074 24868 5080 24880
rect 5000 24840 5080 24868
rect 2685 24803 2743 24809
rect 2685 24769 2697 24803
rect 2731 24800 2743 24803
rect 2774 24800 2780 24812
rect 2731 24772 2780 24800
rect 2731 24769 2743 24772
rect 2685 24763 2743 24769
rect 2774 24760 2780 24772
rect 2832 24760 2838 24812
rect 4798 24760 4804 24812
rect 4856 24800 4862 24812
rect 5000 24809 5028 24840
rect 5074 24828 5080 24840
rect 5132 24828 5138 24880
rect 8202 24868 8208 24880
rect 6472 24840 7052 24868
rect 4893 24803 4951 24809
rect 4893 24800 4905 24803
rect 4856 24772 4905 24800
rect 4856 24760 4862 24772
rect 4893 24769 4905 24772
rect 4939 24769 4951 24803
rect 4893 24763 4951 24769
rect 4985 24803 5043 24809
rect 4985 24769 4997 24803
rect 5031 24769 5043 24803
rect 4985 24763 5043 24769
rect 5169 24803 5227 24809
rect 5169 24769 5181 24803
rect 5215 24800 5227 24803
rect 5626 24800 5632 24812
rect 5215 24772 5632 24800
rect 5215 24769 5227 24772
rect 5169 24763 5227 24769
rect 5626 24760 5632 24772
rect 5684 24760 5690 24812
rect 5813 24803 5871 24809
rect 5813 24769 5825 24803
rect 5859 24800 5871 24803
rect 5997 24803 6055 24809
rect 5859 24772 5948 24800
rect 5859 24769 5871 24772
rect 5813 24763 5871 24769
rect 5077 24735 5135 24741
rect 5077 24701 5089 24735
rect 5123 24732 5135 24735
rect 5920 24732 5948 24772
rect 5997 24769 6009 24803
rect 6043 24800 6055 24803
rect 6472 24800 6500 24840
rect 6043 24772 6500 24800
rect 6549 24803 6607 24809
rect 6043 24769 6055 24772
rect 5997 24763 6055 24769
rect 6549 24769 6561 24803
rect 6595 24769 6607 24803
rect 6730 24800 6736 24812
rect 6643 24772 6736 24800
rect 6549 24763 6607 24769
rect 5123 24704 5948 24732
rect 6564 24732 6592 24763
rect 6730 24760 6736 24772
rect 6788 24760 6794 24812
rect 6914 24800 6920 24812
rect 6875 24772 6920 24800
rect 6914 24760 6920 24772
rect 6972 24760 6978 24812
rect 7024 24800 7052 24840
rect 7668 24840 8208 24868
rect 7190 24800 7196 24812
rect 7024 24772 7196 24800
rect 7190 24760 7196 24772
rect 7248 24760 7254 24812
rect 7668 24809 7696 24840
rect 8202 24828 8208 24840
rect 8260 24828 8266 24880
rect 7653 24803 7711 24809
rect 7653 24769 7665 24803
rect 7699 24769 7711 24803
rect 7653 24763 7711 24769
rect 7742 24760 7748 24812
rect 7800 24800 7806 24812
rect 7837 24803 7895 24809
rect 7837 24800 7849 24803
rect 7800 24772 7849 24800
rect 7800 24760 7806 24772
rect 7837 24769 7849 24772
rect 7883 24800 7895 24803
rect 9306 24800 9312 24812
rect 7883 24772 9312 24800
rect 7883 24769 7895 24772
rect 7837 24763 7895 24769
rect 9306 24760 9312 24772
rect 9364 24760 9370 24812
rect 9585 24803 9643 24809
rect 9585 24769 9597 24803
rect 9631 24800 9643 24803
rect 9766 24800 9772 24812
rect 9631 24772 9772 24800
rect 9631 24769 9643 24772
rect 9585 24763 9643 24769
rect 9766 24760 9772 24772
rect 9824 24760 9830 24812
rect 9876 24809 9904 24908
rect 18874 24896 18880 24948
rect 18932 24936 18938 24948
rect 18932 24908 22608 24936
rect 18932 24896 18938 24908
rect 19242 24828 19248 24880
rect 19300 24868 19306 24880
rect 21082 24868 21088 24880
rect 19300 24840 19564 24868
rect 19300 24828 19306 24840
rect 9861 24803 9919 24809
rect 9861 24769 9873 24803
rect 9907 24769 9919 24803
rect 9861 24763 9919 24769
rect 10505 24803 10563 24809
rect 10505 24769 10517 24803
rect 10551 24800 10563 24803
rect 10594 24800 10600 24812
rect 10551 24772 10600 24800
rect 10551 24769 10563 24772
rect 10505 24763 10563 24769
rect 6638 24732 6644 24744
rect 6564 24704 6644 24732
rect 5123 24701 5135 24704
rect 5077 24695 5135 24701
rect 5920 24664 5948 24704
rect 6638 24692 6644 24704
rect 6696 24692 6702 24744
rect 6748 24732 6776 24760
rect 8570 24732 8576 24744
rect 6748 24704 8576 24732
rect 8570 24692 8576 24704
rect 8628 24692 8634 24744
rect 9674 24732 9680 24744
rect 9635 24704 9680 24732
rect 9674 24692 9680 24704
rect 9732 24692 9738 24744
rect 9876 24732 9904 24763
rect 10594 24760 10600 24772
rect 10652 24760 10658 24812
rect 10689 24803 10747 24809
rect 10689 24769 10701 24803
rect 10735 24769 10747 24803
rect 10689 24763 10747 24769
rect 10781 24803 10839 24809
rect 10781 24769 10793 24803
rect 10827 24769 10839 24803
rect 10781 24763 10839 24769
rect 9876 24704 10180 24732
rect 7742 24664 7748 24676
rect 5920 24636 7748 24664
rect 7742 24624 7748 24636
rect 7800 24624 7806 24676
rect 10152 24664 10180 24704
rect 10226 24692 10232 24744
rect 10284 24732 10290 24744
rect 10704 24732 10732 24763
rect 10284 24704 10732 24732
rect 10796 24732 10824 24763
rect 10870 24760 10876 24812
rect 10928 24800 10934 24812
rect 11146 24800 11152 24812
rect 10928 24772 11152 24800
rect 10928 24760 10934 24772
rect 11146 24760 11152 24772
rect 11204 24760 11210 24812
rect 14369 24803 14427 24809
rect 14369 24769 14381 24803
rect 14415 24800 14427 24803
rect 14826 24800 14832 24812
rect 14415 24772 14832 24800
rect 14415 24769 14427 24772
rect 14369 24763 14427 24769
rect 14826 24760 14832 24772
rect 14884 24760 14890 24812
rect 16850 24800 16856 24812
rect 16811 24772 16856 24800
rect 16850 24760 16856 24772
rect 16908 24760 16914 24812
rect 17678 24800 17684 24812
rect 17639 24772 17684 24800
rect 17678 24760 17684 24772
rect 17736 24760 17742 24812
rect 17862 24800 17868 24812
rect 17823 24772 17868 24800
rect 17862 24760 17868 24772
rect 17920 24760 17926 24812
rect 18506 24800 18512 24812
rect 18467 24772 18512 24800
rect 18506 24760 18512 24772
rect 18564 24760 18570 24812
rect 19150 24800 19156 24812
rect 19111 24772 19156 24800
rect 19150 24760 19156 24772
rect 19208 24760 19214 24812
rect 19429 24803 19487 24809
rect 19429 24800 19441 24803
rect 19260 24772 19441 24800
rect 12066 24732 12072 24744
rect 10796 24704 12072 24732
rect 10284 24692 10290 24704
rect 12066 24692 12072 24704
rect 12124 24692 12130 24744
rect 14093 24735 14151 24741
rect 14093 24701 14105 24735
rect 14139 24732 14151 24735
rect 14274 24732 14280 24744
rect 14139 24704 14280 24732
rect 14139 24701 14151 24704
rect 14093 24695 14151 24701
rect 14274 24692 14280 24704
rect 14332 24692 14338 24744
rect 15562 24692 15568 24744
rect 15620 24732 15626 24744
rect 19260 24732 19288 24772
rect 19429 24769 19441 24772
rect 19475 24769 19487 24803
rect 19429 24763 19487 24769
rect 15620 24704 19288 24732
rect 19337 24735 19395 24741
rect 15620 24692 15626 24704
rect 19337 24701 19349 24735
rect 19383 24732 19395 24735
rect 19536 24732 19564 24840
rect 20272 24840 21088 24868
rect 19613 24803 19671 24809
rect 19613 24769 19625 24803
rect 19659 24800 19671 24803
rect 20070 24800 20076 24812
rect 19659 24772 20076 24800
rect 19659 24769 19671 24772
rect 19613 24763 19671 24769
rect 20070 24760 20076 24772
rect 20128 24760 20134 24812
rect 20272 24809 20300 24840
rect 21082 24828 21088 24840
rect 21140 24828 21146 24880
rect 22580 24868 22608 24908
rect 22646 24896 22652 24948
rect 22704 24936 22710 24948
rect 23753 24939 23811 24945
rect 23753 24936 23765 24939
rect 22704 24908 23765 24936
rect 22704 24896 22710 24908
rect 23753 24905 23765 24908
rect 23799 24905 23811 24939
rect 23753 24899 23811 24905
rect 23845 24939 23903 24945
rect 23845 24905 23857 24939
rect 23891 24936 23903 24939
rect 25314 24936 25320 24948
rect 23891 24908 25320 24936
rect 23891 24905 23903 24908
rect 23845 24899 23903 24905
rect 25314 24896 25320 24908
rect 25372 24896 25378 24948
rect 26418 24896 26424 24948
rect 26476 24936 26482 24948
rect 32214 24936 32220 24948
rect 26476 24908 32220 24936
rect 26476 24896 26482 24908
rect 32214 24896 32220 24908
rect 32272 24896 32278 24948
rect 32950 24936 32956 24948
rect 32600 24908 32817 24936
rect 32911 24908 32956 24936
rect 24118 24868 24124 24880
rect 22580 24840 24124 24868
rect 24118 24828 24124 24840
rect 24176 24828 24182 24880
rect 25590 24868 25596 24880
rect 25056 24840 25596 24868
rect 20257 24803 20315 24809
rect 20257 24769 20269 24803
rect 20303 24769 20315 24803
rect 22741 24803 22799 24809
rect 22741 24800 22753 24803
rect 20257 24763 20315 24769
rect 20364 24772 22753 24800
rect 19383 24704 19564 24732
rect 19383 24701 19395 24704
rect 19337 24695 19395 24701
rect 19978 24692 19984 24744
rect 20036 24732 20042 24744
rect 20364 24732 20392 24772
rect 22741 24769 22753 24772
rect 22787 24769 22799 24803
rect 22741 24763 22799 24769
rect 23017 24803 23075 24809
rect 23017 24769 23029 24803
rect 23063 24800 23075 24803
rect 23474 24800 23480 24812
rect 23063 24772 23480 24800
rect 23063 24769 23075 24772
rect 23017 24763 23075 24769
rect 20036 24704 20392 24732
rect 20533 24735 20591 24741
rect 20036 24692 20042 24704
rect 20533 24701 20545 24735
rect 20579 24732 20591 24735
rect 22756 24732 22784 24763
rect 23474 24760 23480 24772
rect 23532 24760 23538 24812
rect 23934 24809 23940 24812
rect 23921 24803 23940 24809
rect 23921 24769 23933 24803
rect 23921 24763 23940 24769
rect 23934 24760 23940 24763
rect 23992 24760 23998 24812
rect 25056 24800 25084 24840
rect 25590 24828 25596 24840
rect 25648 24828 25654 24880
rect 27982 24868 27988 24880
rect 27448 24840 27988 24868
rect 25222 24800 25228 24812
rect 24228 24772 25084 24800
rect 25183 24772 25228 24800
rect 23106 24732 23112 24744
rect 20579 24704 22094 24732
rect 22756 24704 23112 24732
rect 20579 24701 20591 24704
rect 20533 24695 20591 24701
rect 18417 24667 18475 24673
rect 10152 24636 12434 24664
rect 4065 24599 4123 24605
rect 4065 24565 4077 24599
rect 4111 24596 4123 24599
rect 4430 24596 4436 24608
rect 4111 24568 4436 24596
rect 4111 24565 4123 24568
rect 4065 24559 4123 24565
rect 4430 24556 4436 24568
rect 4488 24596 4494 24608
rect 5166 24596 5172 24608
rect 4488 24568 5172 24596
rect 4488 24556 4494 24568
rect 5166 24556 5172 24568
rect 5224 24556 5230 24608
rect 7650 24596 7656 24608
rect 7611 24568 7656 24596
rect 7650 24556 7656 24568
rect 7708 24556 7714 24608
rect 9306 24556 9312 24608
rect 9364 24596 9370 24608
rect 9858 24596 9864 24608
rect 9364 24568 9864 24596
rect 9364 24556 9370 24568
rect 9858 24556 9864 24568
rect 9916 24556 9922 24608
rect 10045 24599 10103 24605
rect 10045 24565 10057 24599
rect 10091 24596 10103 24599
rect 10134 24596 10140 24608
rect 10091 24568 10140 24596
rect 10091 24565 10103 24568
rect 10045 24559 10103 24565
rect 10134 24556 10140 24568
rect 10192 24556 10198 24608
rect 10962 24556 10968 24608
rect 11020 24596 11026 24608
rect 11057 24599 11115 24605
rect 11057 24596 11069 24599
rect 11020 24568 11069 24596
rect 11020 24556 11026 24568
rect 11057 24565 11069 24568
rect 11103 24565 11115 24599
rect 12406 24596 12434 24636
rect 18417 24633 18429 24667
rect 18463 24664 18475 24667
rect 19058 24664 19064 24676
rect 18463 24636 19064 24664
rect 18463 24633 18475 24636
rect 18417 24627 18475 24633
rect 19058 24624 19064 24636
rect 19116 24624 19122 24676
rect 19242 24664 19248 24676
rect 19203 24636 19248 24664
rect 19242 24624 19248 24636
rect 19300 24624 19306 24676
rect 19886 24624 19892 24676
rect 19944 24664 19950 24676
rect 20438 24664 20444 24676
rect 19944 24636 20444 24664
rect 19944 24624 19950 24636
rect 20438 24624 20444 24636
rect 20496 24664 20502 24676
rect 20548 24664 20576 24695
rect 20496 24636 20576 24664
rect 22066 24664 22094 24704
rect 23106 24692 23112 24704
rect 23164 24692 23170 24744
rect 23566 24732 23572 24744
rect 23527 24704 23572 24732
rect 23566 24692 23572 24704
rect 23624 24692 23630 24744
rect 24228 24664 24256 24772
rect 25222 24760 25228 24772
rect 25280 24760 25286 24812
rect 25498 24800 25504 24812
rect 25459 24772 25504 24800
rect 25498 24760 25504 24772
rect 25556 24760 25562 24812
rect 27448 24800 27476 24840
rect 27982 24828 27988 24840
rect 28040 24828 28046 24880
rect 31662 24828 31668 24880
rect 31720 24868 31726 24880
rect 32600 24868 32628 24908
rect 31720 24840 32628 24868
rect 32789 24868 32817 24908
rect 32950 24896 32956 24908
rect 33008 24896 33014 24948
rect 33873 24939 33931 24945
rect 33873 24905 33885 24939
rect 33919 24936 33931 24939
rect 33962 24936 33968 24948
rect 33919 24908 33968 24936
rect 33919 24905 33931 24908
rect 33873 24899 33931 24905
rect 33962 24896 33968 24908
rect 34020 24896 34026 24948
rect 37458 24936 37464 24948
rect 37419 24908 37464 24936
rect 37458 24896 37464 24908
rect 37516 24896 37522 24948
rect 37826 24936 37832 24948
rect 37787 24908 37832 24936
rect 37826 24896 37832 24908
rect 37884 24896 37890 24948
rect 33226 24868 33232 24880
rect 31720 24828 31726 24840
rect 25608 24772 27476 24800
rect 27617 24803 27675 24809
rect 24305 24735 24363 24741
rect 24305 24701 24317 24735
rect 24351 24732 24363 24735
rect 25608 24732 25636 24772
rect 27617 24769 27629 24803
rect 27663 24769 27675 24803
rect 27617 24763 27675 24769
rect 24351 24704 25636 24732
rect 24351 24701 24363 24704
rect 24305 24695 24363 24701
rect 25682 24692 25688 24744
rect 25740 24732 25746 24744
rect 25740 24704 25785 24732
rect 25740 24692 25746 24704
rect 26786 24692 26792 24744
rect 26844 24732 26850 24744
rect 27632 24732 27660 24763
rect 27890 24760 27896 24812
rect 27948 24800 27954 24812
rect 28997 24803 29055 24809
rect 28997 24800 29009 24803
rect 27948 24772 29009 24800
rect 27948 24760 27954 24772
rect 28997 24769 29009 24772
rect 29043 24769 29055 24803
rect 28997 24763 29055 24769
rect 29181 24803 29239 24809
rect 29181 24769 29193 24803
rect 29227 24769 29239 24803
rect 29181 24763 29239 24769
rect 28445 24735 28503 24741
rect 26844 24704 27752 24732
rect 26844 24692 26850 24704
rect 22066 24636 24256 24664
rect 20496 24624 20502 24636
rect 14366 24596 14372 24608
rect 12406 24568 14372 24596
rect 11057 24559 11115 24565
rect 14366 24556 14372 24568
rect 14424 24556 14430 24608
rect 15654 24596 15660 24608
rect 15615 24568 15660 24596
rect 15654 24556 15660 24568
rect 15712 24556 15718 24608
rect 16758 24556 16764 24608
rect 16816 24596 16822 24608
rect 18138 24596 18144 24608
rect 16816 24568 18144 24596
rect 16816 24556 16822 24568
rect 18138 24556 18144 24568
rect 18196 24556 18202 24608
rect 18969 24599 19027 24605
rect 18969 24565 18981 24599
rect 19015 24596 19027 24599
rect 20254 24596 20260 24608
rect 19015 24568 20260 24596
rect 19015 24565 19027 24568
rect 18969 24559 19027 24565
rect 20254 24556 20260 24568
rect 20312 24556 20318 24608
rect 22554 24596 22560 24608
rect 22515 24568 22560 24596
rect 22554 24556 22560 24568
rect 22612 24556 22618 24608
rect 22738 24556 22744 24608
rect 22796 24596 22802 24608
rect 22925 24599 22983 24605
rect 22925 24596 22937 24599
rect 22796 24568 22937 24596
rect 22796 24556 22802 24568
rect 22925 24565 22937 24568
rect 22971 24565 22983 24599
rect 27724 24596 27752 24704
rect 28445 24701 28457 24735
rect 28491 24732 28503 24735
rect 28534 24732 28540 24744
rect 28491 24704 28540 24732
rect 28491 24701 28503 24704
rect 28445 24695 28503 24701
rect 28534 24692 28540 24704
rect 28592 24692 28598 24744
rect 29196 24732 29224 24763
rect 29270 24760 29276 24812
rect 29328 24800 29334 24812
rect 29328 24772 29373 24800
rect 29328 24760 29334 24772
rect 29638 24760 29644 24812
rect 29696 24800 29702 24812
rect 29733 24803 29791 24809
rect 29733 24800 29745 24803
rect 29696 24772 29745 24800
rect 29696 24760 29702 24772
rect 29733 24769 29745 24772
rect 29779 24769 29791 24803
rect 30006 24800 30012 24812
rect 29967 24772 30012 24800
rect 29733 24763 29791 24769
rect 30006 24760 30012 24772
rect 30064 24760 30070 24812
rect 32309 24803 32367 24809
rect 32309 24769 32321 24803
rect 32355 24769 32367 24803
rect 32309 24763 32367 24769
rect 28736 24704 29224 24732
rect 30469 24735 30527 24741
rect 28258 24624 28264 24676
rect 28316 24664 28322 24676
rect 28736 24664 28764 24704
rect 30469 24701 30481 24735
rect 30515 24732 30527 24735
rect 30515 24704 31754 24732
rect 30515 24701 30527 24704
rect 30469 24695 30527 24701
rect 28994 24664 29000 24676
rect 28316 24636 28764 24664
rect 28955 24636 29000 24664
rect 28316 24624 28322 24636
rect 28994 24624 29000 24636
rect 29052 24624 29058 24676
rect 29822 24664 29828 24676
rect 29783 24636 29828 24664
rect 29822 24624 29828 24636
rect 29880 24624 29886 24676
rect 31726 24664 31754 24704
rect 32030 24664 32036 24676
rect 31726 24636 32036 24664
rect 32030 24624 32036 24636
rect 32088 24624 32094 24676
rect 32324 24664 32352 24763
rect 32399 24760 32405 24812
rect 32457 24800 32463 24812
rect 32600 24809 32628 24840
rect 32585 24803 32643 24809
rect 32457 24772 32502 24800
rect 32457 24760 32463 24772
rect 32585 24769 32597 24803
rect 32631 24769 32643 24803
rect 32585 24763 32643 24769
rect 32674 24794 32680 24846
rect 32732 24794 32738 24846
rect 32789 24840 33232 24868
rect 33226 24828 33232 24840
rect 33284 24828 33290 24880
rect 33505 24871 33563 24877
rect 33505 24837 33517 24871
rect 33551 24868 33563 24871
rect 34054 24868 34060 24880
rect 33551 24840 34060 24868
rect 33551 24837 33563 24840
rect 33505 24831 33563 24837
rect 34054 24828 34060 24840
rect 34112 24828 34118 24880
rect 36081 24871 36139 24877
rect 36081 24837 36093 24871
rect 36127 24868 36139 24871
rect 36814 24868 36820 24880
rect 36127 24840 36820 24868
rect 36127 24837 36139 24840
rect 36081 24831 36139 24837
rect 36814 24828 36820 24840
rect 36872 24828 36878 24880
rect 32774 24803 32832 24809
rect 32674 24769 32686 24794
rect 32720 24769 32732 24794
rect 32674 24763 32732 24769
rect 32774 24769 32786 24803
rect 32820 24800 32832 24803
rect 33686 24800 33692 24812
rect 32820 24772 32904 24800
rect 33647 24772 33692 24800
rect 32820 24769 32832 24772
rect 32774 24763 32832 24769
rect 32674 24664 32680 24676
rect 32324 24636 32680 24664
rect 32674 24624 32680 24636
rect 32732 24624 32738 24676
rect 29730 24596 29736 24608
rect 27724 24568 29736 24596
rect 22925 24559 22983 24565
rect 29730 24556 29736 24568
rect 29788 24556 29794 24608
rect 30466 24556 30472 24608
rect 30524 24596 30530 24608
rect 32876 24596 32904 24772
rect 33686 24760 33692 24772
rect 33744 24760 33750 24812
rect 34330 24800 34336 24812
rect 34291 24772 34336 24800
rect 34330 24760 34336 24772
rect 34388 24760 34394 24812
rect 34514 24800 34520 24812
rect 34475 24772 34520 24800
rect 34514 24760 34520 24772
rect 34572 24760 34578 24812
rect 34606 24760 34612 24812
rect 34664 24800 34670 24812
rect 35253 24803 35311 24809
rect 34664 24772 34709 24800
rect 34664 24760 34670 24772
rect 35253 24769 35265 24803
rect 35299 24800 35311 24803
rect 35342 24800 35348 24812
rect 35299 24772 35348 24800
rect 35299 24769 35311 24772
rect 35253 24763 35311 24769
rect 35342 24760 35348 24772
rect 35400 24760 35406 24812
rect 37918 24732 37924 24744
rect 37879 24704 37924 24732
rect 37918 24692 37924 24704
rect 37976 24692 37982 24744
rect 38010 24692 38016 24744
rect 38068 24732 38074 24744
rect 38068 24704 38113 24732
rect 38068 24692 38074 24704
rect 34054 24624 34060 24676
rect 34112 24664 34118 24676
rect 34333 24667 34391 24673
rect 34333 24664 34345 24667
rect 34112 24636 34345 24664
rect 34112 24624 34118 24636
rect 34333 24633 34345 24636
rect 34379 24633 34391 24667
rect 34333 24627 34391 24633
rect 34514 24624 34520 24676
rect 34572 24664 34578 24676
rect 36262 24664 36268 24676
rect 34572 24636 36268 24664
rect 34572 24624 34578 24636
rect 36262 24624 36268 24636
rect 36320 24624 36326 24676
rect 30524 24568 32904 24596
rect 30524 24556 30530 24568
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 6825 24395 6883 24401
rect 6825 24361 6837 24395
rect 6871 24392 6883 24395
rect 8386 24392 8392 24404
rect 6871 24364 8392 24392
rect 6871 24361 6883 24364
rect 6825 24355 6883 24361
rect 8386 24352 8392 24364
rect 8444 24352 8450 24404
rect 9398 24352 9404 24404
rect 9456 24392 9462 24404
rect 9493 24395 9551 24401
rect 9493 24392 9505 24395
rect 9456 24364 9505 24392
rect 9456 24352 9462 24364
rect 9493 24361 9505 24364
rect 9539 24361 9551 24395
rect 10410 24392 10416 24404
rect 9493 24355 9551 24361
rect 9646 24364 10416 24392
rect 7190 24284 7196 24336
rect 7248 24324 7254 24336
rect 7926 24324 7932 24336
rect 7248 24296 7932 24324
rect 7248 24284 7254 24296
rect 7926 24284 7932 24296
rect 7984 24284 7990 24336
rect 7208 24256 7236 24284
rect 6656 24228 7236 24256
rect 8481 24259 8539 24265
rect 6656 24197 6684 24228
rect 8481 24225 8493 24259
rect 8527 24256 8539 24259
rect 9646 24256 9674 24364
rect 10410 24352 10416 24364
rect 10468 24352 10474 24404
rect 12066 24392 12072 24404
rect 12027 24364 12072 24392
rect 12066 24352 12072 24364
rect 12124 24392 12130 24404
rect 19242 24392 19248 24404
rect 12124 24364 19248 24392
rect 12124 24352 12130 24364
rect 19242 24352 19248 24364
rect 19300 24352 19306 24404
rect 19352 24364 22094 24392
rect 17678 24284 17684 24336
rect 17736 24324 17742 24336
rect 19352 24324 19380 24364
rect 17736 24296 19380 24324
rect 17736 24284 17742 24296
rect 19886 24284 19892 24336
rect 19944 24324 19950 24336
rect 20073 24327 20131 24333
rect 20073 24324 20085 24327
rect 19944 24296 20085 24324
rect 19944 24284 19950 24296
rect 20073 24293 20085 24296
rect 20119 24293 20131 24327
rect 20073 24287 20131 24293
rect 20165 24327 20223 24333
rect 20165 24293 20177 24327
rect 20211 24324 20223 24327
rect 20346 24324 20352 24336
rect 20211 24296 20352 24324
rect 20211 24293 20223 24296
rect 20165 24287 20223 24293
rect 20346 24284 20352 24296
rect 20404 24324 20410 24336
rect 20530 24324 20536 24336
rect 20404 24296 20536 24324
rect 20404 24284 20410 24296
rect 20530 24284 20536 24296
rect 20588 24284 20594 24336
rect 22066 24324 22094 24364
rect 22370 24352 22376 24404
rect 22428 24392 22434 24404
rect 23382 24392 23388 24404
rect 22428 24364 23388 24392
rect 22428 24352 22434 24364
rect 23382 24352 23388 24364
rect 23440 24352 23446 24404
rect 23845 24395 23903 24401
rect 23845 24361 23857 24395
rect 23891 24392 23903 24395
rect 23934 24392 23940 24404
rect 23891 24364 23940 24392
rect 23891 24361 23903 24364
rect 23845 24355 23903 24361
rect 23934 24352 23940 24364
rect 23992 24352 23998 24404
rect 24578 24352 24584 24404
rect 24636 24392 24642 24404
rect 26510 24392 26516 24404
rect 24636 24364 26516 24392
rect 24636 24352 24642 24364
rect 26510 24352 26516 24364
rect 26568 24352 26574 24404
rect 27890 24392 27896 24404
rect 27851 24364 27896 24392
rect 27890 24352 27896 24364
rect 27948 24352 27954 24404
rect 31294 24392 31300 24404
rect 29840 24364 31300 24392
rect 23566 24324 23572 24336
rect 22066 24296 23572 24324
rect 23566 24284 23572 24296
rect 23624 24324 23630 24336
rect 24857 24327 24915 24333
rect 24857 24324 24869 24327
rect 23624 24296 24869 24324
rect 23624 24284 23630 24296
rect 24857 24293 24869 24296
rect 24903 24293 24915 24327
rect 24857 24287 24915 24293
rect 26142 24284 26148 24336
rect 26200 24324 26206 24336
rect 29840 24324 29868 24364
rect 31294 24352 31300 24364
rect 31352 24352 31358 24404
rect 33597 24395 33655 24401
rect 33597 24361 33609 24395
rect 33643 24392 33655 24395
rect 34330 24392 34336 24404
rect 33643 24364 34336 24392
rect 33643 24361 33655 24364
rect 33597 24355 33655 24361
rect 34330 24352 34336 24364
rect 34388 24352 34394 24404
rect 35250 24324 35256 24336
rect 26200 24296 29868 24324
rect 32416 24296 35256 24324
rect 26200 24284 26206 24296
rect 8527 24228 9674 24256
rect 8527 24225 8539 24228
rect 8481 24219 8539 24225
rect 10502 24216 10508 24268
rect 10560 24256 10566 24268
rect 10689 24259 10747 24265
rect 10689 24256 10701 24259
rect 10560 24228 10701 24256
rect 10560 24216 10566 24228
rect 10689 24225 10701 24228
rect 10735 24225 10747 24259
rect 16758 24256 16764 24268
rect 16719 24228 16764 24256
rect 10689 24219 10747 24225
rect 16758 24216 16764 24228
rect 16816 24216 16822 24268
rect 17218 24256 17224 24268
rect 17131 24228 17224 24256
rect 6641 24191 6699 24197
rect 6641 24157 6653 24191
rect 6687 24157 6699 24191
rect 6641 24151 6699 24157
rect 6748 24160 8432 24188
rect 4154 24080 4160 24132
rect 4212 24120 4218 24132
rect 6748 24120 6776 24160
rect 4212 24092 6776 24120
rect 4212 24080 4218 24092
rect 6822 24080 6828 24132
rect 6880 24120 6886 24132
rect 8202 24120 8208 24132
rect 6880 24092 8208 24120
rect 6880 24080 6886 24092
rect 8202 24080 8208 24092
rect 8260 24080 8266 24132
rect 4798 24012 4804 24064
rect 4856 24052 4862 24064
rect 8113 24055 8171 24061
rect 8113 24052 8125 24055
rect 4856 24024 8125 24052
rect 4856 24012 4862 24024
rect 8113 24021 8125 24024
rect 8159 24021 8171 24055
rect 8294 24052 8300 24064
rect 8255 24024 8300 24052
rect 8113 24015 8171 24021
rect 8294 24012 8300 24024
rect 8352 24012 8358 24064
rect 8404 24052 8432 24160
rect 8754 24148 8760 24200
rect 8812 24188 8818 24200
rect 9214 24188 9220 24200
rect 8812 24160 9220 24188
rect 8812 24148 8818 24160
rect 9214 24148 9220 24160
rect 9272 24188 9278 24200
rect 10962 24197 10968 24200
rect 10956 24188 10968 24197
rect 9272 24160 9536 24188
rect 10923 24160 10968 24188
rect 9272 24148 9278 24160
rect 9306 24120 9312 24132
rect 9267 24092 9312 24120
rect 9306 24080 9312 24092
rect 9364 24080 9370 24132
rect 9508 24129 9536 24160
rect 10956 24151 10968 24160
rect 10962 24148 10968 24151
rect 11020 24148 11026 24200
rect 14274 24188 14280 24200
rect 14235 24160 14280 24188
rect 14274 24148 14280 24160
rect 14332 24148 14338 24200
rect 14366 24148 14372 24200
rect 14424 24188 14430 24200
rect 17144 24197 17172 24228
rect 17218 24216 17224 24228
rect 17276 24256 17282 24268
rect 22370 24256 22376 24268
rect 17276 24228 22376 24256
rect 17276 24216 17282 24228
rect 22370 24216 22376 24228
rect 22428 24216 22434 24268
rect 22848 24228 24072 24256
rect 14533 24191 14591 24197
rect 14533 24188 14545 24191
rect 14424 24160 14545 24188
rect 14424 24148 14430 24160
rect 14533 24157 14545 24160
rect 14579 24157 14591 24191
rect 14533 24151 14591 24157
rect 17129 24191 17187 24197
rect 17129 24157 17141 24191
rect 17175 24157 17187 24191
rect 17310 24188 17316 24200
rect 17271 24160 17316 24188
rect 17129 24151 17187 24157
rect 17310 24148 17316 24160
rect 17368 24148 17374 24200
rect 17497 24191 17555 24197
rect 17497 24157 17509 24191
rect 17543 24157 17555 24191
rect 17497 24151 17555 24157
rect 9493 24123 9551 24129
rect 9493 24089 9505 24123
rect 9539 24089 9551 24123
rect 17512 24120 17540 24151
rect 17586 24148 17592 24200
rect 17644 24188 17650 24200
rect 17681 24191 17739 24197
rect 17681 24188 17693 24191
rect 17644 24160 17693 24188
rect 17644 24148 17650 24160
rect 17681 24157 17693 24160
rect 17727 24157 17739 24191
rect 17681 24151 17739 24157
rect 18693 24191 18751 24197
rect 18693 24157 18705 24191
rect 18739 24188 18751 24191
rect 19150 24188 19156 24200
rect 18739 24160 19156 24188
rect 18739 24157 18751 24160
rect 18693 24151 18751 24157
rect 9493 24083 9551 24089
rect 9600 24092 17540 24120
rect 17696 24120 17724 24151
rect 19150 24148 19156 24160
rect 19208 24148 19214 24200
rect 19981 24191 20039 24197
rect 19981 24157 19993 24191
rect 20027 24157 20039 24191
rect 19981 24151 20039 24157
rect 19886 24120 19892 24132
rect 17696 24092 19892 24120
rect 9600 24052 9628 24092
rect 19886 24080 19892 24092
rect 19944 24080 19950 24132
rect 19996 24120 20024 24151
rect 20254 24148 20260 24200
rect 20312 24188 20318 24200
rect 20993 24191 21051 24197
rect 20312 24160 20357 24188
rect 20312 24148 20318 24160
rect 20993 24157 21005 24191
rect 21039 24188 21051 24191
rect 21818 24188 21824 24200
rect 21039 24160 21824 24188
rect 21039 24157 21051 24160
rect 20993 24151 21051 24157
rect 21818 24148 21824 24160
rect 21876 24148 21882 24200
rect 22649 24191 22707 24197
rect 22649 24157 22661 24191
rect 22695 24188 22707 24191
rect 22738 24188 22744 24200
rect 22695 24160 22744 24188
rect 22695 24157 22707 24160
rect 22649 24151 22707 24157
rect 22738 24148 22744 24160
rect 22796 24148 22802 24200
rect 22848 24197 22876 24228
rect 24044 24200 24072 24228
rect 26160 24228 26464 24256
rect 22833 24191 22891 24197
rect 22833 24157 22845 24191
rect 22879 24157 22891 24191
rect 23014 24188 23020 24200
rect 22975 24160 23020 24188
rect 22833 24151 22891 24157
rect 23014 24148 23020 24160
rect 23072 24148 23078 24200
rect 23290 24188 23296 24200
rect 23251 24160 23296 24188
rect 23290 24148 23296 24160
rect 23348 24148 23354 24200
rect 23382 24148 23388 24200
rect 23440 24188 23446 24200
rect 23845 24191 23903 24197
rect 23845 24188 23857 24191
rect 23440 24160 23857 24188
rect 23440 24148 23446 24160
rect 23845 24157 23857 24160
rect 23891 24157 23903 24191
rect 24026 24188 24032 24200
rect 23987 24160 24032 24188
rect 23845 24151 23903 24157
rect 24026 24148 24032 24160
rect 24084 24148 24090 24200
rect 24673 24191 24731 24197
rect 24673 24157 24685 24191
rect 24719 24157 24731 24191
rect 24673 24151 24731 24157
rect 20809 24123 20867 24129
rect 20809 24120 20821 24123
rect 19996 24092 20821 24120
rect 20809 24089 20821 24092
rect 20855 24120 20867 24123
rect 21358 24120 21364 24132
rect 20855 24092 21364 24120
rect 20855 24089 20867 24092
rect 20809 24083 20867 24089
rect 21358 24080 21364 24092
rect 21416 24120 21422 24132
rect 23032 24120 23060 24148
rect 21416 24092 23060 24120
rect 24688 24120 24716 24151
rect 24762 24148 24768 24200
rect 24820 24188 24826 24200
rect 25958 24188 25964 24200
rect 24820 24160 24865 24188
rect 25919 24160 25964 24188
rect 24820 24148 24826 24160
rect 25958 24148 25964 24160
rect 26016 24148 26022 24200
rect 26160 24197 26188 24228
rect 26145 24191 26203 24197
rect 26145 24157 26157 24191
rect 26191 24157 26203 24191
rect 26326 24188 26332 24200
rect 26287 24160 26332 24188
rect 26145 24151 26203 24157
rect 26326 24148 26332 24160
rect 26384 24148 26390 24200
rect 26436 24188 26464 24228
rect 26510 24216 26516 24268
rect 26568 24256 26574 24268
rect 29822 24256 29828 24268
rect 26568 24228 29828 24256
rect 26568 24216 26574 24228
rect 29822 24216 29828 24228
rect 29880 24256 29886 24268
rect 30009 24259 30067 24265
rect 30009 24256 30021 24259
rect 29880 24228 30021 24256
rect 29880 24216 29886 24228
rect 30009 24225 30021 24228
rect 30055 24225 30067 24259
rect 30558 24256 30564 24268
rect 30009 24219 30067 24225
rect 30116 24228 30564 24256
rect 26694 24188 26700 24200
rect 26436 24160 26700 24188
rect 26694 24148 26700 24160
rect 26752 24148 26758 24200
rect 27154 24148 27160 24200
rect 27212 24188 27218 24200
rect 27430 24197 27436 24200
rect 27249 24191 27307 24197
rect 27249 24188 27261 24191
rect 27212 24160 27261 24188
rect 27212 24148 27218 24160
rect 27249 24157 27261 24160
rect 27295 24157 27307 24191
rect 27249 24151 27307 24157
rect 27397 24191 27436 24197
rect 27397 24157 27409 24191
rect 27397 24151 27436 24157
rect 27430 24148 27436 24151
rect 27488 24148 27494 24200
rect 27798 24197 27804 24200
rect 27755 24191 27804 24197
rect 27755 24157 27767 24191
rect 27801 24157 27804 24191
rect 27755 24151 27804 24157
rect 27798 24148 27804 24151
rect 27856 24148 27862 24200
rect 27890 24148 27896 24200
rect 27948 24188 27954 24200
rect 29270 24188 29276 24200
rect 27948 24160 29276 24188
rect 27948 24148 27954 24160
rect 29270 24148 29276 24160
rect 29328 24148 29334 24200
rect 29917 24191 29975 24197
rect 29917 24157 29929 24191
rect 29963 24188 29975 24191
rect 30116 24188 30144 24228
rect 30558 24216 30564 24228
rect 30616 24216 30622 24268
rect 30653 24259 30711 24265
rect 30653 24225 30665 24259
rect 30699 24256 30711 24259
rect 31662 24256 31668 24268
rect 30699 24228 31668 24256
rect 30699 24225 30711 24228
rect 30653 24219 30711 24225
rect 31662 24216 31668 24228
rect 31720 24256 31726 24268
rect 32416 24256 32444 24296
rect 35250 24284 35256 24296
rect 35308 24284 35314 24336
rect 31720 24228 32444 24256
rect 31720 24216 31726 24228
rect 29963 24160 30144 24188
rect 30193 24191 30251 24197
rect 29963 24157 29975 24160
rect 29917 24151 29975 24157
rect 30193 24157 30205 24191
rect 30239 24157 30251 24191
rect 30193 24151 30251 24157
rect 31849 24191 31907 24197
rect 31849 24157 31861 24191
rect 31895 24157 31907 24191
rect 31849 24151 31907 24157
rect 24946 24120 24952 24132
rect 24688 24092 24952 24120
rect 21416 24080 21422 24092
rect 24946 24080 24952 24092
rect 25004 24080 25010 24132
rect 26237 24123 26295 24129
rect 26237 24089 26249 24123
rect 26283 24120 26295 24123
rect 26418 24120 26424 24132
rect 26283 24092 26424 24120
rect 26283 24089 26295 24092
rect 26237 24083 26295 24089
rect 26418 24080 26424 24092
rect 26476 24080 26482 24132
rect 27522 24120 27528 24132
rect 27483 24092 27528 24120
rect 27522 24080 27528 24092
rect 27580 24080 27586 24132
rect 27617 24123 27675 24129
rect 27617 24089 27629 24123
rect 27663 24120 27675 24123
rect 28074 24120 28080 24132
rect 27663 24092 28080 24120
rect 27663 24089 27675 24092
rect 27617 24083 27675 24089
rect 28074 24080 28080 24092
rect 28132 24080 28138 24132
rect 28350 24080 28356 24132
rect 28408 24120 28414 24132
rect 30006 24120 30012 24132
rect 28408 24092 30012 24120
rect 28408 24080 28414 24092
rect 30006 24080 30012 24092
rect 30064 24120 30070 24132
rect 30208 24120 30236 24151
rect 30064 24092 30236 24120
rect 31864 24120 31892 24151
rect 31938 24148 31944 24200
rect 31996 24188 32002 24200
rect 31996 24160 32041 24188
rect 31996 24148 32002 24160
rect 32122 24148 32128 24200
rect 32180 24188 32186 24200
rect 32370 24197 32398 24228
rect 32582 24216 32588 24268
rect 32640 24256 32646 24268
rect 32640 24228 33272 24256
rect 32640 24216 32646 24228
rect 32353 24191 32411 24197
rect 32180 24160 32225 24188
rect 32180 24148 32186 24160
rect 32353 24157 32365 24191
rect 32399 24157 32411 24191
rect 32353 24151 32411 24157
rect 32674 24148 32680 24200
rect 32732 24188 32738 24200
rect 33134 24197 33140 24200
rect 32953 24191 33011 24197
rect 32953 24188 32965 24191
rect 32732 24160 32965 24188
rect 32732 24148 32738 24160
rect 32953 24157 32965 24160
rect 32999 24157 33011 24191
rect 32953 24151 33011 24157
rect 33101 24191 33140 24197
rect 33101 24157 33113 24191
rect 33101 24151 33140 24157
rect 33134 24148 33140 24151
rect 33192 24148 33198 24200
rect 33244 24188 33272 24228
rect 33418 24191 33476 24197
rect 33418 24188 33430 24191
rect 33244 24160 33430 24188
rect 33418 24157 33430 24160
rect 33464 24157 33476 24191
rect 37826 24188 37832 24200
rect 37787 24160 37832 24188
rect 33418 24151 33476 24157
rect 37826 24148 37832 24160
rect 37884 24148 37890 24200
rect 32217 24123 32275 24129
rect 31864 24092 31984 24120
rect 30064 24080 30070 24092
rect 8404 24024 9628 24052
rect 9677 24055 9735 24061
rect 9677 24021 9689 24055
rect 9723 24052 9735 24055
rect 10226 24052 10232 24064
rect 9723 24024 10232 24052
rect 9723 24021 9735 24024
rect 9677 24015 9735 24021
rect 10226 24012 10232 24024
rect 10284 24012 10290 24064
rect 15657 24055 15715 24061
rect 15657 24021 15669 24055
rect 15703 24052 15715 24055
rect 17586 24052 17592 24064
rect 15703 24024 17592 24052
rect 15703 24021 15715 24024
rect 15657 24015 15715 24021
rect 17586 24012 17592 24024
rect 17644 24012 17650 24064
rect 18138 24052 18144 24064
rect 18099 24024 18144 24052
rect 18138 24012 18144 24024
rect 18196 24012 18202 24064
rect 18782 24052 18788 24064
rect 18743 24024 18788 24052
rect 18782 24012 18788 24024
rect 18840 24012 18846 24064
rect 19797 24055 19855 24061
rect 19797 24021 19809 24055
rect 19843 24052 19855 24055
rect 20990 24052 20996 24064
rect 19843 24024 20996 24052
rect 19843 24021 19855 24024
rect 19797 24015 19855 24021
rect 20990 24012 20996 24024
rect 21048 24012 21054 24064
rect 21082 24012 21088 24064
rect 21140 24052 21146 24064
rect 22646 24052 22652 24064
rect 21140 24024 21185 24052
rect 22607 24024 22652 24052
rect 21140 24012 21146 24024
rect 22646 24012 22652 24024
rect 22704 24012 22710 24064
rect 25498 24012 25504 24064
rect 25556 24052 25562 24064
rect 26513 24055 26571 24061
rect 26513 24052 26525 24055
rect 25556 24024 26525 24052
rect 25556 24012 25562 24024
rect 26513 24021 26525 24024
rect 26559 24021 26571 24055
rect 27540 24052 27568 24080
rect 31956 24064 31984 24092
rect 32217 24089 32229 24123
rect 32263 24120 32275 24123
rect 33226 24120 33232 24132
rect 32263 24092 32444 24120
rect 33187 24092 33232 24120
rect 32263 24089 32275 24092
rect 32217 24083 32275 24089
rect 32416 24064 32444 24092
rect 33226 24080 33232 24092
rect 33284 24080 33290 24132
rect 33318 24080 33324 24132
rect 33376 24120 33382 24132
rect 38102 24120 38108 24132
rect 33376 24092 33421 24120
rect 38063 24092 38108 24120
rect 33376 24080 33382 24092
rect 38102 24080 38108 24092
rect 38160 24080 38166 24132
rect 28534 24052 28540 24064
rect 27540 24024 28540 24052
rect 26513 24015 26571 24021
rect 28534 24012 28540 24024
rect 28592 24012 28598 24064
rect 29178 24012 29184 24064
rect 29236 24052 29242 24064
rect 29546 24052 29552 24064
rect 29236 24024 29552 24052
rect 29236 24012 29242 24024
rect 29546 24012 29552 24024
rect 29604 24012 29610 24064
rect 31938 24012 31944 24064
rect 31996 24012 32002 24064
rect 32398 24012 32404 24064
rect 32456 24012 32462 24064
rect 32493 24055 32551 24061
rect 32493 24021 32505 24055
rect 32539 24052 32551 24055
rect 32582 24052 32588 24064
rect 32539 24024 32588 24052
rect 32539 24021 32551 24024
rect 32493 24015 32551 24021
rect 32582 24012 32588 24024
rect 32640 24012 32646 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 4065 23851 4123 23857
rect 4065 23817 4077 23851
rect 4111 23848 4123 23851
rect 4154 23848 4160 23860
rect 4111 23820 4160 23848
rect 4111 23817 4123 23820
rect 4065 23811 4123 23817
rect 4154 23808 4160 23820
rect 4212 23808 4218 23860
rect 5534 23848 5540 23860
rect 5000 23820 5540 23848
rect 4614 23740 4620 23792
rect 4672 23780 4678 23792
rect 4672 23752 4844 23780
rect 4672 23740 4678 23752
rect 2685 23715 2743 23721
rect 2685 23681 2697 23715
rect 2731 23712 2743 23715
rect 2774 23712 2780 23724
rect 2731 23684 2780 23712
rect 2731 23681 2743 23684
rect 2685 23675 2743 23681
rect 2774 23672 2780 23684
rect 2832 23672 2838 23724
rect 2952 23715 3010 23721
rect 2952 23681 2964 23715
rect 2998 23712 3010 23715
rect 3970 23712 3976 23724
rect 2998 23684 3976 23712
rect 2998 23681 3010 23684
rect 2952 23675 3010 23681
rect 3970 23672 3976 23684
rect 4028 23672 4034 23724
rect 4706 23712 4712 23724
rect 4667 23684 4712 23712
rect 4706 23672 4712 23684
rect 4764 23672 4770 23724
rect 4816 23721 4844 23752
rect 5000 23721 5028 23820
rect 5534 23808 5540 23820
rect 5592 23808 5598 23860
rect 16850 23848 16856 23860
rect 5644 23820 16856 23848
rect 5166 23740 5172 23792
rect 5224 23780 5230 23792
rect 5644 23780 5672 23820
rect 16850 23808 16856 23820
rect 16908 23808 16914 23860
rect 18782 23808 18788 23860
rect 18840 23848 18846 23860
rect 21085 23851 21143 23857
rect 21085 23848 21097 23851
rect 18840 23820 21097 23848
rect 18840 23808 18846 23820
rect 21085 23817 21097 23820
rect 21131 23817 21143 23851
rect 21085 23811 21143 23817
rect 21174 23808 21180 23860
rect 21232 23848 21238 23860
rect 23290 23848 23296 23860
rect 21232 23820 23296 23848
rect 21232 23808 21238 23820
rect 23290 23808 23296 23820
rect 23348 23808 23354 23860
rect 23382 23808 23388 23860
rect 23440 23848 23446 23860
rect 23440 23820 25176 23848
rect 23440 23808 23446 23820
rect 7006 23780 7012 23792
rect 5224 23752 5672 23780
rect 6012 23752 7012 23780
rect 5224 23740 5230 23752
rect 4801 23715 4859 23721
rect 4801 23681 4813 23715
rect 4847 23681 4859 23715
rect 4801 23675 4859 23681
rect 4985 23715 5043 23721
rect 4985 23681 4997 23715
rect 5031 23681 5043 23715
rect 4985 23675 5043 23681
rect 5077 23715 5135 23721
rect 5077 23681 5089 23715
rect 5123 23712 5135 23715
rect 5537 23715 5595 23721
rect 5537 23712 5549 23715
rect 5123 23684 5549 23712
rect 5123 23681 5135 23684
rect 5077 23675 5135 23681
rect 5537 23681 5549 23684
rect 5583 23681 5595 23715
rect 5537 23675 5595 23681
rect 5721 23715 5779 23721
rect 5721 23681 5733 23715
rect 5767 23712 5779 23715
rect 5810 23712 5816 23724
rect 5767 23684 5816 23712
rect 5767 23681 5779 23684
rect 5721 23675 5779 23681
rect 4816 23576 4844 23675
rect 5810 23672 5816 23684
rect 5868 23672 5874 23724
rect 6012 23721 6040 23752
rect 7006 23740 7012 23752
rect 7064 23780 7070 23792
rect 7190 23780 7196 23792
rect 7064 23752 7196 23780
rect 7064 23740 7070 23752
rect 7190 23740 7196 23752
rect 7248 23740 7254 23792
rect 7285 23783 7343 23789
rect 7285 23749 7297 23783
rect 7331 23780 7343 23783
rect 7466 23780 7472 23792
rect 7331 23752 7472 23780
rect 7331 23749 7343 23752
rect 7285 23743 7343 23749
rect 5997 23715 6055 23721
rect 5997 23681 6009 23715
rect 6043 23681 6055 23715
rect 6822 23712 6828 23724
rect 5997 23675 6055 23681
rect 6564 23684 6828 23712
rect 5828 23644 5856 23672
rect 6564 23644 6592 23684
rect 6822 23672 6828 23684
rect 6880 23672 6886 23724
rect 7098 23712 7104 23724
rect 7059 23684 7104 23712
rect 7098 23672 7104 23684
rect 7156 23672 7162 23724
rect 5828 23616 6592 23644
rect 6638 23604 6644 23656
rect 6696 23644 6702 23656
rect 7300 23644 7328 23743
rect 7466 23740 7472 23752
rect 7524 23740 7530 23792
rect 15838 23780 15844 23792
rect 9324 23752 15844 23780
rect 7377 23715 7435 23721
rect 7377 23681 7389 23715
rect 7423 23681 7435 23715
rect 7377 23675 7435 23681
rect 6696 23616 7328 23644
rect 7392 23644 7420 23675
rect 8110 23672 8116 23724
rect 8168 23712 8174 23724
rect 8386 23712 8392 23724
rect 8168 23684 8392 23712
rect 8168 23672 8174 23684
rect 8386 23672 8392 23684
rect 8444 23672 8450 23724
rect 9324 23721 9352 23752
rect 15838 23740 15844 23752
rect 15896 23780 15902 23792
rect 16022 23780 16028 23792
rect 15896 23752 16028 23780
rect 15896 23740 15902 23752
rect 16022 23740 16028 23752
rect 16080 23740 16086 23792
rect 19705 23783 19763 23789
rect 19705 23749 19717 23783
rect 19751 23780 19763 23783
rect 21266 23780 21272 23792
rect 19751 23752 21272 23780
rect 19751 23749 19763 23752
rect 19705 23743 19763 23749
rect 21266 23740 21272 23752
rect 21324 23740 21330 23792
rect 23124 23752 23796 23780
rect 9309 23715 9367 23721
rect 9309 23681 9321 23715
rect 9355 23681 9367 23715
rect 9309 23675 9367 23681
rect 9674 23672 9680 23724
rect 9732 23712 9738 23724
rect 10413 23715 10471 23721
rect 10413 23712 10425 23715
rect 9732 23684 10425 23712
rect 9732 23672 9738 23684
rect 10413 23681 10425 23684
rect 10459 23712 10471 23715
rect 11146 23712 11152 23724
rect 10459 23684 11152 23712
rect 10459 23681 10471 23684
rect 10413 23675 10471 23681
rect 11146 23672 11152 23684
rect 11204 23672 11210 23724
rect 14458 23672 14464 23724
rect 14516 23712 14522 23724
rect 18046 23712 18052 23724
rect 14516 23684 18052 23712
rect 14516 23672 14522 23684
rect 18046 23672 18052 23684
rect 18104 23672 18110 23724
rect 19889 23715 19947 23721
rect 19889 23681 19901 23715
rect 19935 23681 19947 23715
rect 19889 23675 19947 23681
rect 20993 23715 21051 23721
rect 20993 23681 21005 23715
rect 21039 23712 21051 23715
rect 22830 23712 22836 23724
rect 21039 23684 22836 23712
rect 21039 23681 21051 23684
rect 20993 23675 21051 23681
rect 8662 23644 8668 23656
rect 7392 23616 8668 23644
rect 6696 23604 6702 23616
rect 8662 23604 8668 23616
rect 8720 23604 8726 23656
rect 9493 23647 9551 23653
rect 9493 23613 9505 23647
rect 9539 23613 9551 23647
rect 9493 23607 9551 23613
rect 10229 23647 10287 23653
rect 10229 23613 10241 23647
rect 10275 23644 10287 23647
rect 10275 23616 10732 23644
rect 10275 23613 10287 23616
rect 10229 23607 10287 23613
rect 8202 23576 8208 23588
rect 4816 23548 8208 23576
rect 8202 23536 8208 23548
rect 8260 23536 8266 23588
rect 9306 23536 9312 23588
rect 9364 23576 9370 23588
rect 9508 23576 9536 23607
rect 9364 23548 9536 23576
rect 9364 23536 9370 23548
rect 10704 23520 10732 23616
rect 19904 23576 19932 23675
rect 22830 23672 22836 23684
rect 22888 23672 22894 23724
rect 21269 23647 21327 23653
rect 21269 23613 21281 23647
rect 21315 23644 21327 23647
rect 21358 23644 21364 23656
rect 21315 23616 21364 23644
rect 21315 23613 21327 23616
rect 21269 23607 21327 23613
rect 21358 23604 21364 23616
rect 21416 23604 21422 23656
rect 23124 23576 23152 23752
rect 23768 23724 23796 23752
rect 24026 23740 24032 23792
rect 24084 23780 24090 23792
rect 24857 23783 24915 23789
rect 24857 23780 24869 23783
rect 24084 23752 24869 23780
rect 24084 23740 24090 23752
rect 24857 23749 24869 23752
rect 24903 23749 24915 23783
rect 24857 23743 24915 23749
rect 23201 23715 23259 23721
rect 23201 23681 23213 23715
rect 23247 23681 23259 23715
rect 23201 23675 23259 23681
rect 23216 23644 23244 23675
rect 23290 23672 23296 23724
rect 23348 23712 23354 23724
rect 23385 23715 23443 23721
rect 23385 23712 23397 23715
rect 23348 23684 23397 23712
rect 23348 23672 23354 23684
rect 23385 23681 23397 23684
rect 23431 23681 23443 23715
rect 23750 23712 23756 23724
rect 23711 23684 23756 23712
rect 23385 23675 23443 23681
rect 23750 23672 23756 23684
rect 23808 23672 23814 23724
rect 24946 23672 24952 23724
rect 25004 23712 25010 23724
rect 25041 23715 25099 23721
rect 25041 23712 25053 23715
rect 25004 23684 25053 23712
rect 25004 23672 25010 23684
rect 25041 23681 25053 23684
rect 25087 23681 25099 23715
rect 25148 23712 25176 23820
rect 25682 23808 25688 23860
rect 25740 23848 25746 23860
rect 26602 23848 26608 23860
rect 25740 23820 26608 23848
rect 25740 23808 25746 23820
rect 26602 23808 26608 23820
rect 26660 23848 26666 23860
rect 26660 23820 27476 23848
rect 26660 23808 26666 23820
rect 25225 23783 25283 23789
rect 25225 23749 25237 23783
rect 25271 23780 25283 23783
rect 26786 23780 26792 23792
rect 25271 23752 26792 23780
rect 25271 23749 25283 23752
rect 25225 23743 25283 23749
rect 26786 23740 26792 23752
rect 26844 23740 26850 23792
rect 27154 23780 27160 23792
rect 27115 23752 27160 23780
rect 27154 23740 27160 23752
rect 27212 23740 27218 23792
rect 27448 23780 27476 23820
rect 27706 23808 27712 23860
rect 27764 23848 27770 23860
rect 27764 23820 28304 23848
rect 27764 23808 27770 23820
rect 27890 23780 27896 23792
rect 27448 23752 27896 23780
rect 25685 23715 25743 23721
rect 25685 23712 25697 23715
rect 25148 23684 25697 23712
rect 25041 23675 25099 23681
rect 25685 23681 25697 23684
rect 25731 23681 25743 23715
rect 25685 23675 25743 23681
rect 26237 23715 26295 23721
rect 26237 23681 26249 23715
rect 26283 23712 26295 23715
rect 26326 23712 26332 23724
rect 26283 23684 26332 23712
rect 26283 23681 26295 23684
rect 26237 23675 26295 23681
rect 26326 23672 26332 23684
rect 26384 23712 26390 23724
rect 26970 23712 26976 23724
rect 26384 23684 26976 23712
rect 26384 23672 26390 23684
rect 26970 23672 26976 23684
rect 27028 23672 27034 23724
rect 27338 23672 27344 23724
rect 27396 23712 27402 23724
rect 27632 23721 27660 23752
rect 27890 23740 27896 23752
rect 27948 23740 27954 23792
rect 27617 23715 27675 23721
rect 27396 23684 27441 23712
rect 27396 23672 27402 23684
rect 27617 23681 27629 23715
rect 27663 23681 27675 23715
rect 28276 23712 28304 23820
rect 28810 23808 28816 23860
rect 28868 23808 28874 23860
rect 29454 23808 29460 23860
rect 29512 23848 29518 23860
rect 31294 23848 31300 23860
rect 29512 23820 31300 23848
rect 29512 23808 29518 23820
rect 31294 23808 31300 23820
rect 31352 23808 31358 23860
rect 31938 23808 31944 23860
rect 31996 23848 32002 23860
rect 33042 23848 33048 23860
rect 31996 23820 33048 23848
rect 31996 23808 32002 23820
rect 33042 23808 33048 23820
rect 33100 23808 33106 23860
rect 33134 23808 33140 23860
rect 33192 23848 33198 23860
rect 37734 23848 37740 23860
rect 33192 23820 37740 23848
rect 33192 23808 33198 23820
rect 28626 23740 28632 23792
rect 28684 23780 28690 23792
rect 28684 23752 28729 23780
rect 28684 23740 28690 23752
rect 28353 23715 28411 23721
rect 28353 23712 28365 23715
rect 28276 23684 28365 23712
rect 27617 23675 27675 23681
rect 28353 23681 28365 23684
rect 28399 23681 28411 23715
rect 28353 23675 28411 23681
rect 28491 23715 28549 23721
rect 28491 23681 28503 23715
rect 28537 23681 28549 23715
rect 28491 23675 28549 23681
rect 28745 23715 28803 23721
rect 28745 23681 28757 23715
rect 28791 23710 28803 23715
rect 28833 23710 28861 23808
rect 30653 23783 30711 23789
rect 30653 23749 30665 23783
rect 30699 23780 30711 23783
rect 31386 23780 31392 23792
rect 30699 23752 31392 23780
rect 30699 23749 30711 23752
rect 30653 23743 30711 23749
rect 31386 23740 31392 23752
rect 31444 23740 31450 23792
rect 32122 23740 32128 23792
rect 32180 23780 32186 23792
rect 32766 23780 32772 23792
rect 32180 23752 32772 23780
rect 32180 23740 32186 23752
rect 32766 23740 32772 23752
rect 32824 23780 32830 23792
rect 32824 23752 32996 23780
rect 32824 23740 32830 23752
rect 29914 23712 29920 23724
rect 28791 23682 28861 23710
rect 29875 23684 29920 23712
rect 28791 23681 28803 23682
rect 28745 23675 28803 23681
rect 24964 23644 24992 23672
rect 23216 23616 24992 23644
rect 26053 23647 26111 23653
rect 26053 23613 26065 23647
rect 26099 23613 26111 23647
rect 26053 23607 26111 23613
rect 26145 23647 26203 23653
rect 26145 23613 26157 23647
rect 26191 23644 26203 23647
rect 27062 23644 27068 23656
rect 26191 23616 27068 23644
rect 26191 23613 26203 23616
rect 26145 23607 26203 23613
rect 23658 23576 23664 23588
rect 19904 23548 23152 23576
rect 23619 23548 23664 23576
rect 23658 23536 23664 23548
rect 23716 23536 23722 23588
rect 26068 23576 26096 23607
rect 27062 23604 27068 23616
rect 27120 23604 27126 23656
rect 28516 23644 28544 23675
rect 29914 23672 29920 23684
rect 29972 23672 29978 23724
rect 30193 23715 30251 23721
rect 30193 23681 30205 23715
rect 30239 23681 30251 23715
rect 32582 23712 32588 23724
rect 32543 23684 32588 23712
rect 30193 23675 30251 23681
rect 29638 23644 29644 23656
rect 28516 23616 29644 23644
rect 29638 23604 29644 23616
rect 29696 23604 29702 23656
rect 29822 23604 29828 23656
rect 29880 23644 29886 23656
rect 30208 23644 30236 23675
rect 32582 23672 32588 23684
rect 32640 23672 32646 23724
rect 32968 23721 32996 23752
rect 32677 23715 32735 23721
rect 32677 23681 32689 23715
rect 32723 23681 32735 23715
rect 32677 23675 32735 23681
rect 32953 23715 33011 23721
rect 32953 23681 32965 23715
rect 32999 23681 33011 23715
rect 33060 23712 33088 23808
rect 34422 23740 34428 23792
rect 34480 23780 34486 23792
rect 35176 23789 35204 23820
rect 37734 23808 37740 23820
rect 37792 23808 37798 23860
rect 37826 23808 37832 23860
rect 37884 23808 37890 23860
rect 35069 23783 35127 23789
rect 35069 23780 35081 23783
rect 34480 23752 35081 23780
rect 34480 23740 34486 23752
rect 35069 23749 35081 23752
rect 35115 23749 35127 23783
rect 35069 23743 35127 23749
rect 35161 23783 35219 23789
rect 35161 23749 35173 23783
rect 35207 23749 35219 23783
rect 35161 23743 35219 23749
rect 35897 23783 35955 23789
rect 35897 23749 35909 23783
rect 35943 23780 35955 23783
rect 37844 23780 37872 23808
rect 37921 23783 37979 23789
rect 37921 23780 37933 23783
rect 35943 23752 37933 23780
rect 35943 23749 35955 23752
rect 35897 23743 35955 23749
rect 37921 23749 37933 23752
rect 37967 23749 37979 23783
rect 37921 23743 37979 23749
rect 34790 23712 34796 23724
rect 33060 23684 34796 23712
rect 32953 23675 33011 23681
rect 29880 23616 30236 23644
rect 29880 23604 29886 23616
rect 30650 23604 30656 23656
rect 30708 23644 30714 23656
rect 32692 23644 32720 23675
rect 34790 23672 34796 23684
rect 34848 23672 34854 23724
rect 34882 23672 34888 23724
rect 34940 23712 34946 23724
rect 35250 23712 35256 23724
rect 35308 23721 35314 23724
rect 34940 23684 34985 23712
rect 35216 23684 35256 23712
rect 34940 23672 34946 23684
rect 35250 23672 35256 23684
rect 35308 23675 35316 23721
rect 36081 23715 36139 23721
rect 36081 23712 36093 23715
rect 35452 23684 36093 23712
rect 35308 23672 35314 23675
rect 30708 23616 32720 23644
rect 30708 23604 30714 23616
rect 27890 23576 27896 23588
rect 26068 23548 27896 23576
rect 27890 23536 27896 23548
rect 27948 23536 27954 23588
rect 30006 23576 30012 23588
rect 28828 23548 30012 23576
rect 4525 23511 4583 23517
rect 4525 23477 4537 23511
rect 4571 23508 4583 23511
rect 4614 23508 4620 23520
rect 4571 23480 4620 23508
rect 4571 23477 4583 23480
rect 4525 23471 4583 23477
rect 4614 23468 4620 23480
rect 4672 23468 4678 23520
rect 5350 23468 5356 23520
rect 5408 23508 5414 23520
rect 5902 23508 5908 23520
rect 5408 23480 5908 23508
rect 5408 23468 5414 23480
rect 5902 23468 5908 23480
rect 5960 23468 5966 23520
rect 6914 23508 6920 23520
rect 6875 23480 6920 23508
rect 6914 23468 6920 23480
rect 6972 23468 6978 23520
rect 8481 23511 8539 23517
rect 8481 23477 8493 23511
rect 8527 23508 8539 23511
rect 8570 23508 8576 23520
rect 8527 23480 8576 23508
rect 8527 23477 8539 23480
rect 8481 23471 8539 23477
rect 8570 23468 8576 23480
rect 8628 23468 8634 23520
rect 10594 23508 10600 23520
rect 10555 23480 10600 23508
rect 10594 23468 10600 23480
rect 10652 23468 10658 23520
rect 10686 23468 10692 23520
rect 10744 23508 10750 23520
rect 12434 23508 12440 23520
rect 10744 23480 12440 23508
rect 10744 23468 10750 23480
rect 12434 23468 12440 23480
rect 12492 23468 12498 23520
rect 16298 23468 16304 23520
rect 16356 23508 16362 23520
rect 16482 23508 16488 23520
rect 16356 23480 16488 23508
rect 16356 23468 16362 23480
rect 16482 23468 16488 23480
rect 16540 23508 16546 23520
rect 19886 23508 19892 23520
rect 16540 23480 19892 23508
rect 16540 23468 16546 23480
rect 19886 23468 19892 23480
rect 19944 23468 19950 23520
rect 20070 23508 20076 23520
rect 20031 23480 20076 23508
rect 20070 23468 20076 23480
rect 20128 23468 20134 23520
rect 20530 23468 20536 23520
rect 20588 23508 20594 23520
rect 20625 23511 20683 23517
rect 20625 23508 20637 23511
rect 20588 23480 20637 23508
rect 20588 23468 20594 23480
rect 20625 23477 20637 23480
rect 20671 23477 20683 23511
rect 20625 23471 20683 23477
rect 26234 23468 26240 23520
rect 26292 23508 26298 23520
rect 27525 23511 27583 23517
rect 27525 23508 27537 23511
rect 26292 23480 27537 23508
rect 26292 23468 26298 23480
rect 27525 23477 27537 23480
rect 27571 23508 27583 23511
rect 28350 23508 28356 23520
rect 27571 23480 28356 23508
rect 27571 23477 27583 23480
rect 27525 23471 27583 23477
rect 28350 23468 28356 23480
rect 28408 23468 28414 23520
rect 28626 23468 28632 23520
rect 28684 23508 28690 23520
rect 28828 23508 28856 23548
rect 30006 23536 30012 23548
rect 30064 23536 30070 23588
rect 35452 23585 35480 23684
rect 36081 23681 36093 23684
rect 36127 23681 36139 23715
rect 36081 23675 36139 23681
rect 36170 23672 36176 23724
rect 36228 23712 36234 23724
rect 36449 23715 36507 23721
rect 36228 23684 36273 23712
rect 36228 23672 36234 23684
rect 36449 23681 36461 23715
rect 36495 23712 36507 23715
rect 36495 23684 36667 23712
rect 36495 23681 36507 23684
rect 36449 23675 36507 23681
rect 36357 23647 36415 23653
rect 36357 23613 36369 23647
rect 36403 23644 36415 23647
rect 36538 23644 36544 23656
rect 36403 23616 36544 23644
rect 36403 23613 36415 23616
rect 36357 23607 36415 23613
rect 36538 23604 36544 23616
rect 36596 23604 36602 23656
rect 32401 23579 32459 23585
rect 32401 23545 32413 23579
rect 32447 23576 32459 23579
rect 35437 23579 35495 23585
rect 32447 23548 35389 23576
rect 32447 23545 32459 23548
rect 32401 23539 32459 23545
rect 28948 23517 28954 23520
rect 28684 23480 28856 23508
rect 28905 23511 28954 23517
rect 28684 23468 28690 23480
rect 28905 23477 28917 23511
rect 28951 23477 28954 23511
rect 28905 23471 28954 23477
rect 28948 23468 28954 23471
rect 29006 23508 29012 23520
rect 32861 23511 32919 23517
rect 29006 23480 29053 23508
rect 29006 23468 29012 23480
rect 32861 23477 32873 23511
rect 32907 23508 32919 23511
rect 32950 23508 32956 23520
rect 32907 23480 32956 23508
rect 32907 23477 32919 23480
rect 32861 23471 32919 23477
rect 32950 23468 32956 23480
rect 33008 23468 33014 23520
rect 35361 23508 35389 23548
rect 35437 23545 35449 23579
rect 35483 23545 35495 23579
rect 35437 23539 35495 23545
rect 35618 23536 35624 23588
rect 35676 23576 35682 23588
rect 36262 23576 36268 23588
rect 35676 23548 36268 23576
rect 35676 23536 35682 23548
rect 36262 23536 36268 23548
rect 36320 23576 36326 23588
rect 36639 23576 36667 23684
rect 37734 23672 37740 23724
rect 37792 23712 37798 23724
rect 37829 23715 37887 23721
rect 37829 23712 37841 23715
rect 37792 23684 37841 23712
rect 37792 23672 37798 23684
rect 37829 23681 37841 23684
rect 37875 23681 37887 23715
rect 37829 23675 37887 23681
rect 38010 23644 38016 23656
rect 37971 23616 38016 23644
rect 38010 23604 38016 23616
rect 38068 23604 38074 23656
rect 37918 23576 37924 23588
rect 36320 23548 36667 23576
rect 36924 23548 37924 23576
rect 36320 23536 36326 23548
rect 36924 23508 36952 23548
rect 37918 23536 37924 23548
rect 37976 23536 37982 23588
rect 35361 23480 36952 23508
rect 36998 23468 37004 23520
rect 37056 23508 37062 23520
rect 37461 23511 37519 23517
rect 37461 23508 37473 23511
rect 37056 23480 37473 23508
rect 37056 23468 37062 23480
rect 37461 23477 37473 23480
rect 37507 23477 37519 23511
rect 37461 23471 37519 23477
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 3970 23304 3976 23316
rect 3931 23276 3976 23304
rect 3970 23264 3976 23276
rect 4028 23264 4034 23316
rect 5902 23264 5908 23316
rect 5960 23304 5966 23316
rect 10505 23307 10563 23313
rect 5960 23276 7788 23304
rect 5960 23264 5966 23276
rect 6914 23236 6920 23248
rect 6875 23208 6920 23236
rect 6914 23196 6920 23208
rect 6972 23196 6978 23248
rect 4525 23171 4583 23177
rect 4525 23137 4537 23171
rect 4571 23168 4583 23171
rect 4798 23168 4804 23180
rect 4571 23140 4804 23168
rect 4571 23137 4583 23140
rect 4525 23131 4583 23137
rect 4798 23128 4804 23140
rect 4856 23128 4862 23180
rect 5994 23128 6000 23180
rect 6052 23168 6058 23180
rect 6825 23171 6883 23177
rect 6052 23140 6776 23168
rect 6052 23128 6058 23140
rect 6748 23112 6776 23140
rect 6825 23137 6837 23171
rect 6871 23168 6883 23171
rect 7190 23168 7196 23180
rect 6871 23140 7196 23168
rect 6871 23137 6883 23140
rect 6825 23131 6883 23137
rect 7190 23128 7196 23140
rect 7248 23128 7254 23180
rect 4154 23060 4160 23112
rect 4212 23100 4218 23112
rect 4341 23103 4399 23109
rect 4341 23100 4353 23103
rect 4212 23072 4353 23100
rect 4212 23060 4218 23072
rect 4341 23069 4353 23072
rect 4387 23069 4399 23103
rect 4341 23063 4399 23069
rect 4433 23103 4491 23109
rect 4433 23069 4445 23103
rect 4479 23100 4491 23103
rect 4614 23100 4620 23112
rect 4479 23072 4620 23100
rect 4479 23069 4491 23072
rect 4433 23063 4491 23069
rect 4614 23060 4620 23072
rect 4672 23060 4678 23112
rect 4890 23060 4896 23112
rect 4948 23100 4954 23112
rect 5813 23103 5871 23109
rect 5813 23100 5825 23103
rect 4948 23072 5825 23100
rect 4948 23060 4954 23072
rect 5813 23069 5825 23072
rect 5859 23100 5871 23103
rect 6638 23100 6644 23112
rect 5859 23072 6644 23100
rect 5859 23069 5871 23072
rect 5813 23063 5871 23069
rect 6638 23060 6644 23072
rect 6696 23060 6702 23112
rect 6730 23060 6736 23112
rect 6788 23100 6794 23112
rect 6788 23072 6881 23100
rect 6788 23060 6794 23072
rect 6914 23060 6920 23112
rect 6972 23100 6978 23112
rect 7760 23109 7788 23276
rect 10505 23273 10517 23307
rect 10551 23304 10563 23307
rect 10686 23304 10692 23316
rect 10551 23276 10692 23304
rect 10551 23273 10563 23276
rect 10505 23267 10563 23273
rect 10686 23264 10692 23276
rect 10744 23264 10750 23316
rect 15654 23264 15660 23316
rect 15712 23304 15718 23316
rect 20714 23304 20720 23316
rect 15712 23276 20720 23304
rect 15712 23264 15718 23276
rect 20714 23264 20720 23276
rect 20772 23264 20778 23316
rect 21266 23304 21272 23316
rect 21227 23276 21272 23304
rect 21266 23264 21272 23276
rect 21324 23264 21330 23316
rect 22554 23304 22560 23316
rect 22515 23276 22560 23304
rect 22554 23264 22560 23276
rect 22612 23264 22618 23316
rect 34977 23307 35035 23313
rect 34977 23273 34989 23307
rect 35023 23304 35035 23307
rect 36170 23304 36176 23316
rect 35023 23276 36176 23304
rect 35023 23273 35035 23276
rect 34977 23267 35035 23273
rect 36170 23264 36176 23276
rect 36228 23264 36234 23316
rect 37734 23264 37740 23316
rect 37792 23304 37798 23316
rect 38105 23307 38163 23313
rect 38105 23304 38117 23307
rect 37792 23276 38117 23304
rect 37792 23264 37798 23276
rect 38105 23273 38117 23276
rect 38151 23273 38163 23307
rect 38105 23267 38163 23273
rect 15194 23196 15200 23248
rect 15252 23236 15258 23248
rect 15289 23239 15347 23245
rect 15289 23236 15301 23239
rect 15252 23208 15301 23236
rect 15252 23196 15258 23208
rect 15289 23205 15301 23208
rect 15335 23205 15347 23239
rect 23109 23239 23167 23245
rect 23109 23236 23121 23239
rect 15289 23199 15347 23205
rect 18708 23208 23121 23236
rect 14274 23128 14280 23180
rect 14332 23168 14338 23180
rect 14332 23140 16988 23168
rect 14332 23128 14338 23140
rect 7009 23103 7067 23109
rect 7009 23100 7021 23103
rect 6972 23072 7021 23100
rect 6972 23060 6978 23072
rect 7009 23069 7021 23072
rect 7055 23069 7067 23103
rect 7009 23063 7067 23069
rect 7745 23103 7803 23109
rect 7745 23069 7757 23103
rect 7791 23069 7803 23103
rect 7745 23063 7803 23069
rect 8021 23103 8079 23109
rect 8021 23069 8033 23103
rect 8067 23100 8079 23103
rect 8662 23100 8668 23112
rect 8067 23072 8668 23100
rect 8067 23069 8079 23072
rect 8021 23063 8079 23069
rect 8662 23060 8668 23072
rect 8720 23060 8726 23112
rect 9122 23100 9128 23112
rect 9083 23072 9128 23100
rect 9122 23060 9128 23072
rect 9180 23060 9186 23112
rect 12069 23103 12127 23109
rect 12069 23069 12081 23103
rect 12115 23100 12127 23103
rect 14292 23100 14320 23128
rect 12115 23072 14320 23100
rect 14645 23103 14703 23109
rect 12115 23069 12127 23072
rect 12069 23063 12127 23069
rect 14645 23069 14657 23103
rect 14691 23100 14703 23103
rect 15378 23100 15384 23112
rect 14691 23072 15384 23100
rect 14691 23069 14703 23072
rect 14645 23063 14703 23069
rect 5905 23035 5963 23041
rect 5905 23001 5917 23035
rect 5951 23032 5963 23035
rect 5951 23004 7972 23032
rect 5951 23001 5963 23004
rect 5905 22995 5963 23001
rect 6549 22967 6607 22973
rect 6549 22933 6561 22967
rect 6595 22964 6607 22967
rect 7190 22964 7196 22976
rect 6595 22936 7196 22964
rect 6595 22933 6607 22936
rect 6549 22927 6607 22933
rect 7190 22924 7196 22936
rect 7248 22924 7254 22976
rect 7558 22964 7564 22976
rect 7519 22936 7564 22964
rect 7558 22924 7564 22936
rect 7616 22924 7622 22976
rect 7944 22973 7972 23004
rect 8938 22992 8944 23044
rect 8996 23032 9002 23044
rect 12342 23041 12348 23044
rect 9370 23035 9428 23041
rect 9370 23032 9382 23035
rect 8996 23004 9382 23032
rect 8996 22992 9002 23004
rect 9370 23001 9382 23004
rect 9416 23001 9428 23035
rect 12336 23032 12348 23041
rect 12303 23004 12348 23032
rect 9370 22995 9428 23001
rect 12336 22995 12348 23004
rect 12342 22992 12348 22995
rect 12400 22992 12406 23044
rect 7929 22967 7987 22973
rect 7929 22933 7941 22967
rect 7975 22964 7987 22967
rect 9858 22964 9864 22976
rect 7975 22936 9864 22964
rect 7975 22933 7987 22936
rect 7929 22927 7987 22933
rect 9858 22924 9864 22936
rect 9916 22924 9922 22976
rect 12066 22924 12072 22976
rect 12124 22964 12130 22976
rect 13449 22967 13507 22973
rect 13449 22964 13461 22967
rect 12124 22936 13461 22964
rect 12124 22924 12130 22936
rect 13449 22933 13461 22936
rect 13495 22964 13507 22967
rect 14660 22964 14688 23063
rect 15378 23060 15384 23072
rect 15436 23060 15442 23112
rect 15565 23103 15623 23109
rect 15565 23069 15577 23103
rect 15611 23100 15623 23103
rect 15654 23100 15660 23112
rect 15611 23072 15660 23100
rect 15611 23069 15623 23072
rect 15565 23063 15623 23069
rect 15654 23060 15660 23072
rect 15712 23060 15718 23112
rect 15746 23060 15752 23112
rect 15804 23100 15810 23112
rect 16960 23109 16988 23140
rect 16025 23103 16083 23109
rect 16025 23100 16037 23103
rect 15804 23072 16037 23100
rect 15804 23060 15810 23072
rect 16025 23069 16037 23072
rect 16071 23069 16083 23103
rect 16025 23063 16083 23069
rect 16945 23103 17003 23109
rect 16945 23069 16957 23103
rect 16991 23100 17003 23103
rect 18414 23100 18420 23112
rect 16991 23072 18420 23100
rect 16991 23069 17003 23072
rect 16945 23063 17003 23069
rect 18414 23060 18420 23072
rect 18472 23060 18478 23112
rect 17218 23041 17224 23044
rect 15289 23035 15347 23041
rect 15289 23001 15301 23035
rect 15335 23032 15347 23035
rect 15335 23004 17172 23032
rect 15335 23001 15347 23004
rect 15289 22995 15347 23001
rect 13495 22936 14688 22964
rect 14737 22967 14795 22973
rect 13495 22933 13507 22936
rect 13449 22927 13507 22933
rect 14737 22933 14749 22967
rect 14783 22964 14795 22967
rect 15473 22967 15531 22973
rect 15473 22964 15485 22967
rect 14783 22936 15485 22964
rect 14783 22933 14795 22936
rect 14737 22927 14795 22933
rect 15473 22933 15485 22936
rect 15519 22933 15531 22967
rect 15473 22927 15531 22933
rect 16022 22924 16028 22976
rect 16080 22964 16086 22976
rect 16117 22967 16175 22973
rect 16117 22964 16129 22967
rect 16080 22936 16129 22964
rect 16080 22924 16086 22936
rect 16117 22933 16129 22936
rect 16163 22933 16175 22967
rect 17144 22964 17172 23004
rect 17212 22995 17224 23041
rect 17276 23032 17282 23044
rect 18708 23032 18736 23208
rect 23109 23205 23121 23208
rect 23155 23205 23167 23239
rect 23109 23199 23167 23205
rect 31938 23196 31944 23248
rect 31996 23236 32002 23248
rect 32950 23236 32956 23248
rect 31996 23208 32956 23236
rect 31996 23196 32002 23208
rect 32950 23196 32956 23208
rect 33008 23236 33014 23248
rect 36538 23236 36544 23248
rect 33008 23208 36544 23236
rect 33008 23196 33014 23208
rect 36538 23196 36544 23208
rect 36596 23196 36602 23248
rect 20530 23168 20536 23180
rect 20491 23140 20536 23168
rect 20530 23128 20536 23140
rect 20588 23128 20594 23180
rect 20622 23128 20628 23180
rect 20680 23168 20686 23180
rect 20898 23168 20904 23180
rect 20680 23140 20904 23168
rect 20680 23128 20686 23140
rect 20898 23128 20904 23140
rect 20956 23128 20962 23180
rect 20990 23128 20996 23180
rect 21048 23168 21054 23180
rect 21821 23171 21879 23177
rect 21821 23168 21833 23171
rect 21048 23140 21833 23168
rect 21048 23128 21054 23140
rect 21821 23137 21833 23140
rect 21867 23137 21879 23171
rect 23198 23168 23204 23180
rect 21821 23131 21879 23137
rect 22480 23140 23204 23168
rect 18966 23060 18972 23112
rect 19024 23100 19030 23112
rect 22480 23109 22508 23140
rect 23198 23128 23204 23140
rect 23256 23128 23262 23180
rect 25406 23128 25412 23180
rect 25464 23168 25470 23180
rect 26697 23171 26755 23177
rect 25464 23140 26648 23168
rect 25464 23128 25470 23140
rect 22465 23103 22523 23109
rect 19024 23072 21864 23100
rect 19024 23060 19030 23072
rect 21729 23035 21787 23041
rect 21729 23032 21741 23035
rect 17276 23004 17312 23032
rect 18156 23004 18736 23032
rect 20088 23004 21741 23032
rect 17218 22992 17224 22995
rect 17276 22992 17282 23004
rect 18156 22964 18184 23004
rect 18322 22964 18328 22976
rect 17144 22936 18184 22964
rect 18283 22936 18328 22964
rect 16117 22927 16175 22933
rect 18322 22924 18328 22936
rect 18380 22924 18386 22976
rect 20088 22973 20116 23004
rect 21729 23001 21741 23004
rect 21775 23001 21787 23035
rect 21836 23032 21864 23072
rect 22465 23069 22477 23103
rect 22511 23069 22523 23103
rect 22465 23063 22523 23069
rect 22741 23103 22799 23109
rect 22741 23069 22753 23103
rect 22787 23069 22799 23103
rect 22741 23063 22799 23069
rect 22925 23103 22983 23109
rect 22925 23069 22937 23103
rect 22971 23100 22983 23103
rect 24762 23100 24768 23112
rect 22971 23072 24768 23100
rect 22971 23069 22983 23072
rect 22925 23063 22983 23069
rect 22756 23032 22784 23063
rect 24762 23060 24768 23072
rect 24820 23060 24826 23112
rect 25961 23103 26019 23109
rect 25961 23069 25973 23103
rect 26007 23100 26019 23103
rect 26234 23100 26240 23112
rect 26007 23072 26240 23100
rect 26007 23069 26019 23072
rect 25961 23063 26019 23069
rect 26234 23060 26240 23072
rect 26292 23060 26298 23112
rect 26620 23109 26648 23140
rect 26697 23137 26709 23171
rect 26743 23168 26755 23171
rect 27338 23168 27344 23180
rect 26743 23140 27344 23168
rect 26743 23137 26755 23140
rect 26697 23131 26755 23137
rect 27338 23128 27344 23140
rect 27396 23128 27402 23180
rect 27890 23128 27896 23180
rect 27948 23168 27954 23180
rect 29638 23168 29644 23180
rect 27948 23140 28764 23168
rect 27948 23128 27954 23140
rect 28736 23112 28764 23140
rect 28966 23140 29644 23168
rect 28966 23112 28994 23140
rect 29638 23128 29644 23140
rect 29696 23128 29702 23180
rect 29914 23128 29920 23180
rect 29972 23168 29978 23180
rect 29972 23140 30696 23168
rect 29972 23128 29978 23140
rect 26605 23103 26663 23109
rect 26605 23069 26617 23103
rect 26651 23069 26663 23103
rect 26605 23063 26663 23069
rect 26786 23060 26792 23112
rect 26844 23100 26850 23112
rect 26881 23103 26939 23109
rect 26881 23100 26893 23103
rect 26844 23072 26893 23100
rect 26844 23060 26850 23072
rect 26881 23069 26893 23072
rect 26927 23069 26939 23103
rect 26881 23063 26939 23069
rect 27706 23060 27712 23112
rect 27764 23100 27770 23112
rect 27801 23103 27859 23109
rect 27801 23100 27813 23103
rect 27764 23072 27813 23100
rect 27764 23060 27770 23072
rect 27801 23069 27813 23072
rect 27847 23069 27859 23103
rect 27982 23100 27988 23112
rect 27943 23072 27988 23100
rect 27801 23063 27859 23069
rect 27982 23060 27988 23072
rect 28040 23060 28046 23112
rect 28626 23109 28632 23112
rect 28445 23103 28503 23109
rect 28445 23069 28457 23103
rect 28491 23069 28503 23103
rect 28445 23063 28503 23069
rect 28593 23103 28632 23109
rect 28593 23069 28605 23103
rect 28593 23063 28632 23069
rect 21836 23004 22784 23032
rect 27893 23035 27951 23041
rect 21729 22995 21787 23001
rect 27893 23001 27905 23035
rect 27939 23032 27951 23035
rect 28460 23032 28488 23063
rect 28626 23060 28632 23063
rect 28684 23060 28690 23112
rect 28718 23060 28724 23112
rect 28776 23100 28782 23112
rect 28776 23072 28869 23100
rect 28776 23060 28782 23072
rect 28902 23060 28908 23112
rect 28960 23100 28994 23112
rect 28960 23072 29053 23100
rect 28960 23063 28968 23072
rect 28960 23060 28966 23063
rect 29270 23060 29276 23112
rect 29328 23100 29334 23112
rect 29822 23100 29828 23112
rect 29328 23072 29828 23100
rect 29328 23060 29334 23072
rect 29822 23060 29828 23072
rect 29880 23060 29886 23112
rect 30006 23060 30012 23112
rect 30064 23100 30070 23112
rect 30668 23109 30696 23140
rect 31294 23128 31300 23180
rect 31352 23168 31358 23180
rect 35621 23171 35679 23177
rect 35621 23168 35633 23171
rect 31352 23140 35633 23168
rect 31352 23128 31358 23140
rect 35621 23137 35633 23140
rect 35667 23168 35679 23171
rect 35802 23168 35808 23180
rect 35667 23140 35808 23168
rect 35667 23137 35679 23140
rect 35621 23131 35679 23137
rect 35802 23128 35808 23140
rect 35860 23128 35866 23180
rect 30285 23103 30343 23109
rect 30285 23100 30297 23103
rect 30064 23072 30297 23100
rect 30064 23060 30070 23072
rect 30285 23069 30297 23072
rect 30331 23069 30343 23103
rect 30285 23063 30343 23069
rect 30653 23103 30711 23109
rect 30653 23069 30665 23103
rect 30699 23069 30711 23103
rect 30653 23063 30711 23069
rect 34514 23060 34520 23112
rect 34572 23100 34578 23112
rect 35161 23103 35219 23109
rect 35161 23100 35173 23103
rect 34572 23072 35173 23100
rect 34572 23060 34578 23072
rect 35161 23069 35173 23072
rect 35207 23069 35219 23103
rect 35161 23063 35219 23069
rect 35253 23103 35311 23109
rect 35253 23069 35265 23103
rect 35299 23069 35311 23103
rect 35526 23100 35532 23112
rect 35487 23072 35532 23100
rect 35253 23063 35311 23069
rect 27939 23004 28488 23032
rect 28813 23035 28871 23041
rect 27939 23001 27951 23004
rect 27893 22995 27951 23001
rect 28813 23001 28825 23035
rect 28859 23032 28871 23035
rect 31846 23032 31852 23044
rect 28859 23004 31852 23032
rect 28859 23001 28871 23004
rect 28813 22995 28871 23001
rect 31846 22992 31852 23004
rect 31904 22992 31910 23044
rect 20073 22967 20131 22973
rect 20073 22933 20085 22967
rect 20119 22933 20131 22967
rect 20438 22964 20444 22976
rect 20399 22936 20444 22964
rect 20073 22927 20131 22933
rect 20438 22924 20444 22936
rect 20496 22924 20502 22976
rect 21634 22964 21640 22976
rect 21595 22936 21640 22964
rect 21634 22924 21640 22936
rect 21692 22924 21698 22976
rect 24486 22924 24492 22976
rect 24544 22964 24550 22976
rect 29089 22967 29147 22973
rect 29089 22964 29101 22967
rect 24544 22936 29101 22964
rect 24544 22924 24550 22936
rect 29089 22933 29101 22936
rect 29135 22933 29147 22967
rect 29089 22927 29147 22933
rect 29454 22924 29460 22976
rect 29512 22964 29518 22976
rect 29914 22964 29920 22976
rect 29512 22936 29920 22964
rect 29512 22924 29518 22936
rect 29914 22924 29920 22936
rect 29972 22924 29978 22976
rect 30926 22964 30932 22976
rect 30887 22936 30932 22964
rect 30926 22924 30932 22936
rect 30984 22964 30990 22976
rect 35268 22964 35296 23063
rect 35526 23060 35532 23072
rect 35584 23060 35590 23112
rect 36725 23103 36783 23109
rect 36725 23069 36737 23103
rect 36771 23100 36783 23103
rect 36814 23100 36820 23112
rect 36771 23072 36820 23100
rect 36771 23069 36783 23072
rect 36725 23063 36783 23069
rect 36814 23060 36820 23072
rect 36872 23060 36878 23112
rect 36998 23109 37004 23112
rect 36992 23100 37004 23109
rect 36959 23072 37004 23100
rect 36992 23063 37004 23072
rect 36998 23060 37004 23063
rect 37056 23060 37062 23112
rect 35434 22964 35440 22976
rect 30984 22936 35440 22964
rect 30984 22924 30990 22936
rect 35434 22924 35440 22936
rect 35492 22924 35498 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 4706 22720 4712 22772
rect 4764 22760 4770 22772
rect 4801 22763 4859 22769
rect 4801 22760 4813 22763
rect 4764 22732 4813 22760
rect 4764 22720 4770 22732
rect 4801 22729 4813 22732
rect 4847 22729 4859 22763
rect 4801 22723 4859 22729
rect 6638 22720 6644 22772
rect 6696 22760 6702 22772
rect 7098 22760 7104 22772
rect 6696 22732 7104 22760
rect 6696 22720 6702 22732
rect 7098 22720 7104 22732
rect 7156 22720 7162 22772
rect 8938 22760 8944 22772
rect 8899 22732 8944 22760
rect 8938 22720 8944 22732
rect 8996 22720 9002 22772
rect 12342 22760 12348 22772
rect 12303 22732 12348 22760
rect 12342 22720 12348 22732
rect 12400 22720 12406 22772
rect 15654 22760 15660 22772
rect 15615 22732 15660 22760
rect 15654 22720 15660 22732
rect 15712 22720 15718 22772
rect 21082 22760 21088 22772
rect 18984 22732 21088 22760
rect 5074 22692 5080 22704
rect 4724 22664 5080 22692
rect 4724 22633 4752 22664
rect 5074 22652 5080 22664
rect 5132 22652 5138 22704
rect 7193 22695 7251 22701
rect 7193 22661 7205 22695
rect 7239 22692 7251 22695
rect 7834 22692 7840 22704
rect 7239 22664 7840 22692
rect 7239 22661 7251 22664
rect 7193 22655 7251 22661
rect 7834 22652 7840 22664
rect 7892 22652 7898 22704
rect 10410 22652 10416 22704
rect 10468 22692 10474 22704
rect 11057 22695 11115 22701
rect 10468 22664 10916 22692
rect 10468 22652 10474 22664
rect 4709 22627 4767 22633
rect 4709 22593 4721 22627
rect 4755 22593 4767 22627
rect 4890 22624 4896 22636
rect 4851 22596 4896 22624
rect 4709 22587 4767 22593
rect 4890 22584 4896 22596
rect 4948 22584 4954 22636
rect 7466 22624 7472 22636
rect 7427 22596 7472 22624
rect 7466 22584 7472 22596
rect 7524 22584 7530 22636
rect 8662 22584 8668 22636
rect 8720 22624 8726 22636
rect 9125 22627 9183 22633
rect 9125 22624 9137 22627
rect 8720 22596 9137 22624
rect 8720 22584 8726 22596
rect 9125 22593 9137 22596
rect 9171 22593 9183 22627
rect 9125 22587 9183 22593
rect 9401 22627 9459 22633
rect 9401 22593 9413 22627
rect 9447 22624 9459 22627
rect 10594 22624 10600 22636
rect 9447 22596 10600 22624
rect 9447 22593 9459 22596
rect 9401 22587 9459 22593
rect 10594 22584 10600 22596
rect 10652 22584 10658 22636
rect 10888 22633 10916 22664
rect 11057 22661 11069 22695
rect 11103 22692 11115 22695
rect 11698 22692 11704 22704
rect 11103 22664 11704 22692
rect 11103 22661 11115 22664
rect 11057 22655 11115 22661
rect 11698 22652 11704 22664
rect 11756 22652 11762 22704
rect 12066 22692 12072 22704
rect 12027 22664 12072 22692
rect 12066 22652 12072 22664
rect 12124 22652 12130 22704
rect 14274 22652 14280 22704
rect 14332 22692 14338 22704
rect 14332 22664 15056 22692
rect 14332 22652 14338 22664
rect 10873 22627 10931 22633
rect 10873 22593 10885 22627
rect 10919 22593 10931 22627
rect 11146 22624 11152 22636
rect 11107 22596 11152 22624
rect 10873 22587 10931 22593
rect 7282 22556 7288 22568
rect 7243 22528 7288 22556
rect 7282 22516 7288 22528
rect 7340 22516 7346 22568
rect 8018 22516 8024 22568
rect 8076 22556 8082 22568
rect 9217 22559 9275 22565
rect 9217 22556 9229 22559
rect 8076 22528 9229 22556
rect 8076 22516 8082 22528
rect 9217 22525 9229 22528
rect 9263 22525 9275 22559
rect 9217 22519 9275 22525
rect 9306 22516 9312 22568
rect 9364 22556 9370 22568
rect 10888 22556 10916 22587
rect 11146 22584 11152 22596
rect 11204 22584 11210 22636
rect 11790 22624 11796 22636
rect 11751 22596 11796 22624
rect 11790 22584 11796 22596
rect 11848 22584 11854 22636
rect 11977 22627 12035 22633
rect 11977 22593 11989 22627
rect 12023 22614 12035 22627
rect 12161 22627 12219 22633
rect 12023 22593 12112 22614
rect 11977 22587 12112 22593
rect 12161 22593 12173 22627
rect 12207 22624 12219 22627
rect 12250 22624 12256 22636
rect 12207 22596 12256 22624
rect 12207 22593 12219 22596
rect 12161 22587 12219 22593
rect 11992 22586 12112 22587
rect 12084 22556 12112 22586
rect 12250 22584 12256 22596
rect 12308 22584 12314 22636
rect 14366 22624 14372 22636
rect 14327 22596 14372 22624
rect 14366 22584 14372 22596
rect 14424 22584 14430 22636
rect 14550 22624 14556 22636
rect 14511 22596 14556 22624
rect 14550 22584 14556 22596
rect 14608 22584 14614 22636
rect 15028 22633 15056 22664
rect 15286 22652 15292 22704
rect 15344 22692 15350 22704
rect 15933 22695 15991 22701
rect 15933 22692 15945 22695
rect 15344 22664 15945 22692
rect 15344 22652 15350 22664
rect 15933 22661 15945 22664
rect 15979 22661 15991 22695
rect 15933 22655 15991 22661
rect 16143 22695 16201 22701
rect 16143 22661 16155 22695
rect 16189 22692 16201 22695
rect 16850 22692 16856 22704
rect 16189 22661 16206 22692
rect 16763 22664 16856 22692
rect 16143 22655 16206 22661
rect 15013 22627 15071 22633
rect 15013 22593 15025 22627
rect 15059 22624 15071 22627
rect 15102 22624 15108 22636
rect 15059 22596 15108 22624
rect 15059 22593 15071 22596
rect 15013 22587 15071 22593
rect 15102 22584 15108 22596
rect 15160 22584 15166 22636
rect 15841 22627 15899 22633
rect 15841 22593 15853 22627
rect 15887 22593 15899 22627
rect 15841 22587 15899 22593
rect 9364 22528 9409 22556
rect 10888 22528 12112 22556
rect 9364 22516 9370 22528
rect 5902 22448 5908 22500
rect 5960 22488 5966 22500
rect 15286 22488 15292 22500
rect 5960 22460 15292 22488
rect 5960 22448 5966 22460
rect 15286 22448 15292 22460
rect 15344 22448 15350 22500
rect 7190 22420 7196 22432
rect 7151 22392 7196 22420
rect 7190 22380 7196 22392
rect 7248 22380 7254 22432
rect 7653 22423 7711 22429
rect 7653 22389 7665 22423
rect 7699 22420 7711 22423
rect 8110 22420 8116 22432
rect 7699 22392 8116 22420
rect 7699 22389 7711 22392
rect 7653 22383 7711 22389
rect 8110 22380 8116 22392
rect 8168 22380 8174 22432
rect 10594 22380 10600 22432
rect 10652 22420 10658 22432
rect 10689 22423 10747 22429
rect 10689 22420 10701 22423
rect 10652 22392 10701 22420
rect 10652 22380 10658 22392
rect 10689 22389 10701 22392
rect 10735 22389 10747 22423
rect 14458 22420 14464 22432
rect 14419 22392 14464 22420
rect 10689 22383 10747 22389
rect 14458 22380 14464 22392
rect 14516 22380 14522 22432
rect 15105 22423 15163 22429
rect 15105 22389 15117 22423
rect 15151 22420 15163 22423
rect 15470 22420 15476 22432
rect 15151 22392 15476 22420
rect 15151 22389 15163 22392
rect 15105 22383 15163 22389
rect 15470 22380 15476 22392
rect 15528 22380 15534 22432
rect 15856 22420 15884 22587
rect 16023 22584 16029 22636
rect 16081 22624 16087 22636
rect 16178 22634 16206 22655
rect 16850 22652 16856 22664
rect 16908 22692 16914 22704
rect 18984 22692 19012 22732
rect 21082 22720 21088 22732
rect 21140 22720 21146 22772
rect 21177 22763 21235 22769
rect 21177 22729 21189 22763
rect 21223 22760 21235 22763
rect 21634 22760 21640 22772
rect 21223 22732 21640 22760
rect 21223 22729 21235 22732
rect 21177 22723 21235 22729
rect 21634 22720 21640 22732
rect 21692 22720 21698 22772
rect 27614 22760 27620 22772
rect 27264 22732 27620 22760
rect 20070 22701 20076 22704
rect 16908 22664 19012 22692
rect 19153 22695 19211 22701
rect 16908 22652 16914 22664
rect 19153 22661 19165 22695
rect 19199 22692 19211 22695
rect 20064 22692 20076 22701
rect 19199 22664 19932 22692
rect 20031 22664 20076 22692
rect 19199 22661 19211 22664
rect 19153 22655 19211 22661
rect 16178 22624 16252 22634
rect 16574 22624 16580 22636
rect 16081 22596 16126 22624
rect 16178 22606 16580 22624
rect 16224 22596 16580 22606
rect 16081 22584 16087 22596
rect 16574 22584 16580 22596
rect 16632 22624 16638 22636
rect 17037 22627 17095 22633
rect 17037 22624 17049 22627
rect 16632 22596 17049 22624
rect 16632 22584 16638 22596
rect 17037 22593 17049 22596
rect 17083 22624 17095 22627
rect 17126 22624 17132 22636
rect 17083 22596 17132 22624
rect 17083 22593 17095 22596
rect 17037 22587 17095 22593
rect 17126 22584 17132 22596
rect 17184 22624 17190 22636
rect 17494 22624 17500 22636
rect 17184 22596 17500 22624
rect 17184 22584 17190 22596
rect 17494 22584 17500 22596
rect 17552 22584 17558 22636
rect 18322 22624 18328 22636
rect 18283 22596 18328 22624
rect 18322 22584 18328 22596
rect 18380 22584 18386 22636
rect 18414 22584 18420 22636
rect 18472 22624 18478 22636
rect 19797 22627 19855 22633
rect 19797 22624 19809 22627
rect 18472 22596 19809 22624
rect 18472 22584 18478 22596
rect 19797 22593 19809 22596
rect 19843 22593 19855 22627
rect 19904 22624 19932 22664
rect 20064 22655 20076 22664
rect 20070 22652 20076 22655
rect 20128 22652 20134 22704
rect 21818 22652 21824 22704
rect 21876 22692 21882 22704
rect 21876 22664 24348 22692
rect 21876 22652 21882 22664
rect 21542 22624 21548 22636
rect 19904 22596 21548 22624
rect 19797 22587 19855 22593
rect 21542 22584 21548 22596
rect 21600 22584 21606 22636
rect 22646 22624 22652 22636
rect 22607 22596 22652 22624
rect 22646 22584 22652 22596
rect 22704 22584 22710 22636
rect 22922 22624 22928 22636
rect 22883 22596 22928 22624
rect 22922 22584 22928 22596
rect 22980 22584 22986 22636
rect 23569 22627 23627 22633
rect 23569 22593 23581 22627
rect 23615 22624 23627 22627
rect 23658 22624 23664 22636
rect 23615 22596 23664 22624
rect 23615 22593 23627 22596
rect 23569 22587 23627 22593
rect 23658 22584 23664 22596
rect 23716 22584 23722 22636
rect 16301 22559 16359 22565
rect 16301 22525 16313 22559
rect 16347 22556 16359 22559
rect 16482 22556 16488 22568
rect 16347 22528 16488 22556
rect 16347 22525 16359 22528
rect 16301 22519 16359 22525
rect 16482 22516 16488 22528
rect 16540 22516 16546 22568
rect 17402 22556 17408 22568
rect 17363 22528 17408 22556
rect 17402 22516 17408 22528
rect 17460 22516 17466 22568
rect 18506 22556 18512 22568
rect 18467 22528 18512 22556
rect 18506 22516 18512 22528
rect 18564 22516 18570 22568
rect 23382 22556 23388 22568
rect 23343 22528 23388 22556
rect 23382 22516 23388 22528
rect 23440 22516 23446 22568
rect 24320 22556 24348 22664
rect 24394 22652 24400 22704
rect 24452 22692 24458 22704
rect 24452 22664 24900 22692
rect 24452 22652 24458 22664
rect 24486 22624 24492 22636
rect 24447 22596 24492 22624
rect 24486 22584 24492 22596
rect 24544 22584 24550 22636
rect 24872 22633 24900 22664
rect 25314 22652 25320 22704
rect 25372 22692 25378 22704
rect 26418 22692 26424 22704
rect 25372 22664 26424 22692
rect 25372 22652 25378 22664
rect 26418 22652 26424 22664
rect 26476 22652 26482 22704
rect 24857 22627 24915 22633
rect 24857 22593 24869 22627
rect 24903 22624 24915 22627
rect 25590 22624 25596 22636
rect 24903 22596 25596 22624
rect 24903 22593 24915 22596
rect 24857 22587 24915 22593
rect 25590 22584 25596 22596
rect 25648 22584 25654 22636
rect 25317 22559 25375 22565
rect 24320 22528 25268 22556
rect 16206 22448 16212 22500
rect 16264 22488 16270 22500
rect 19794 22488 19800 22500
rect 16264 22460 19800 22488
rect 16264 22448 16270 22460
rect 19794 22448 19800 22460
rect 19852 22448 19858 22500
rect 24397 22491 24455 22497
rect 24397 22488 24409 22491
rect 22066 22460 24409 22488
rect 16850 22420 16856 22432
rect 15856 22392 16856 22420
rect 16850 22380 16856 22392
rect 16908 22380 16914 22432
rect 20162 22380 20168 22432
rect 20220 22420 20226 22432
rect 22066 22420 22094 22460
rect 24397 22457 24409 22460
rect 24443 22457 24455 22491
rect 25240 22488 25268 22528
rect 25317 22525 25329 22559
rect 25363 22556 25375 22559
rect 25774 22556 25780 22568
rect 25363 22528 25780 22556
rect 25363 22525 25375 22528
rect 25317 22519 25375 22525
rect 25774 22516 25780 22528
rect 25832 22556 25838 22568
rect 26142 22556 26148 22568
rect 25832 22528 26148 22556
rect 25832 22516 25838 22528
rect 26142 22516 26148 22528
rect 26200 22516 26206 22568
rect 27264 22488 27292 22732
rect 27614 22720 27620 22732
rect 27672 22720 27678 22772
rect 28261 22763 28319 22769
rect 28261 22729 28273 22763
rect 28307 22760 28319 22763
rect 28534 22760 28540 22772
rect 28307 22732 28540 22760
rect 28307 22729 28319 22732
rect 28261 22723 28319 22729
rect 28534 22720 28540 22732
rect 28592 22720 28598 22772
rect 29822 22720 29828 22772
rect 29880 22760 29886 22772
rect 30098 22760 30104 22772
rect 29880 22732 30104 22760
rect 29880 22720 29886 22732
rect 30098 22720 30104 22732
rect 30156 22720 30162 22772
rect 30742 22720 30748 22772
rect 30800 22760 30806 22772
rect 33505 22763 33563 22769
rect 30800 22732 31616 22760
rect 30800 22720 30806 22732
rect 27338 22652 27344 22704
rect 27396 22692 27402 22704
rect 29549 22695 29607 22701
rect 29549 22692 29561 22695
rect 27396 22664 29561 22692
rect 27396 22652 27402 22664
rect 29549 22661 29561 22664
rect 29595 22661 29607 22695
rect 29549 22655 29607 22661
rect 29641 22695 29699 22701
rect 29641 22661 29653 22695
rect 29687 22692 29699 22695
rect 30834 22692 30840 22704
rect 29687 22664 30840 22692
rect 29687 22661 29699 22664
rect 29641 22655 29699 22661
rect 30834 22652 30840 22664
rect 30892 22652 30898 22704
rect 31588 22636 31616 22732
rect 33505 22729 33517 22763
rect 33551 22760 33563 22763
rect 33686 22760 33692 22772
rect 33551 22732 33692 22760
rect 33551 22729 33563 22732
rect 33505 22723 33563 22729
rect 33686 22720 33692 22732
rect 33744 22720 33750 22772
rect 31757 22695 31815 22701
rect 31757 22661 31769 22695
rect 31803 22692 31815 22695
rect 32490 22692 32496 22704
rect 31803 22664 32496 22692
rect 31803 22661 31815 22664
rect 31757 22655 31815 22661
rect 32490 22652 32496 22664
rect 32548 22652 32554 22704
rect 35802 22692 35808 22704
rect 35763 22664 35808 22692
rect 35802 22652 35808 22664
rect 35860 22652 35866 22704
rect 27614 22624 27620 22636
rect 27575 22596 27620 22624
rect 27614 22584 27620 22596
rect 27672 22584 27678 22636
rect 27706 22584 27712 22636
rect 27764 22624 27770 22636
rect 27890 22624 27896 22636
rect 27764 22596 27809 22624
rect 27851 22596 27896 22624
rect 27764 22584 27770 22596
rect 27890 22584 27896 22596
rect 27948 22584 27954 22636
rect 27985 22627 28043 22633
rect 27985 22593 27997 22627
rect 28031 22593 28043 22627
rect 27985 22587 28043 22593
rect 28123 22627 28181 22633
rect 28123 22593 28135 22627
rect 28169 22624 28181 22627
rect 28258 22624 28264 22636
rect 28169 22596 28264 22624
rect 28169 22593 28181 22596
rect 28123 22587 28181 22593
rect 25240 22460 27292 22488
rect 24397 22451 24455 22457
rect 20220 22392 22094 22420
rect 28000 22420 28028 22587
rect 28258 22584 28264 22596
rect 28316 22624 28322 22636
rect 28902 22624 28908 22636
rect 28316 22596 28908 22624
rect 28316 22584 28322 22596
rect 28902 22584 28908 22596
rect 28960 22584 28966 22636
rect 29362 22624 29368 22636
rect 29323 22596 29368 22624
rect 29362 22584 29368 22596
rect 29420 22584 29426 22636
rect 29730 22624 29736 22636
rect 29691 22596 29736 22624
rect 29730 22584 29736 22596
rect 29788 22584 29794 22636
rect 30466 22584 30472 22636
rect 30524 22624 30530 22636
rect 31202 22624 31208 22636
rect 30524 22596 31208 22624
rect 30524 22584 30530 22596
rect 31202 22584 31208 22596
rect 31260 22584 31266 22636
rect 31570 22624 31576 22636
rect 31531 22596 31576 22624
rect 31570 22584 31576 22596
rect 31628 22584 31634 22636
rect 33134 22624 33140 22636
rect 33095 22596 33140 22624
rect 33134 22584 33140 22596
rect 33192 22584 33198 22636
rect 33321 22627 33379 22633
rect 33321 22593 33333 22627
rect 33367 22624 33379 22627
rect 33962 22624 33968 22636
rect 33367 22596 33968 22624
rect 33367 22593 33379 22596
rect 33321 22587 33379 22593
rect 33962 22584 33968 22596
rect 34020 22584 34026 22636
rect 35434 22624 35440 22636
rect 35395 22596 35440 22624
rect 35434 22584 35440 22596
rect 35492 22584 35498 22636
rect 35526 22584 35532 22636
rect 35584 22624 35590 22636
rect 35710 22624 35716 22636
rect 35584 22596 35716 22624
rect 35584 22584 35590 22596
rect 35710 22584 35716 22596
rect 35768 22584 35774 22636
rect 37734 22584 37740 22636
rect 37792 22624 37798 22636
rect 37829 22627 37887 22633
rect 37829 22624 37841 22627
rect 37792 22596 37841 22624
rect 37792 22584 37798 22596
rect 37829 22593 37841 22596
rect 37875 22593 37887 22627
rect 37829 22587 37887 22593
rect 29454 22516 29460 22568
rect 29512 22556 29518 22568
rect 30742 22556 30748 22568
rect 29512 22528 30748 22556
rect 29512 22516 29518 22528
rect 30742 22516 30748 22528
rect 30800 22516 30806 22568
rect 34606 22516 34612 22568
rect 34664 22556 34670 22568
rect 35345 22559 35403 22565
rect 35345 22556 35357 22559
rect 34664 22528 35357 22556
rect 34664 22516 34670 22528
rect 35345 22525 35357 22528
rect 35391 22525 35403 22559
rect 38102 22556 38108 22568
rect 38063 22528 38108 22556
rect 35345 22519 35403 22525
rect 38102 22516 38108 22528
rect 38160 22516 38166 22568
rect 31478 22488 31484 22500
rect 28184 22460 31484 22488
rect 28184 22420 28212 22460
rect 31478 22448 31484 22460
rect 31536 22448 31542 22500
rect 28000 22392 28212 22420
rect 20220 22380 20226 22392
rect 28994 22380 29000 22432
rect 29052 22420 29058 22432
rect 29917 22423 29975 22429
rect 29917 22420 29929 22423
rect 29052 22392 29929 22420
rect 29052 22380 29058 22392
rect 29917 22389 29929 22392
rect 29963 22389 29975 22423
rect 29917 22383 29975 22389
rect 35161 22423 35219 22429
rect 35161 22389 35173 22423
rect 35207 22420 35219 22423
rect 36354 22420 36360 22432
rect 35207 22392 36360 22420
rect 35207 22389 35219 22392
rect 35161 22383 35219 22389
rect 36354 22380 36360 22392
rect 36412 22380 36418 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 7193 22219 7251 22225
rect 7193 22185 7205 22219
rect 7239 22216 7251 22219
rect 7466 22216 7472 22228
rect 7239 22188 7472 22216
rect 7239 22185 7251 22188
rect 7193 22179 7251 22185
rect 7466 22176 7472 22188
rect 7524 22176 7530 22228
rect 11698 22176 11704 22228
rect 11756 22216 11762 22228
rect 11882 22216 11888 22228
rect 11756 22188 11888 22216
rect 11756 22176 11762 22188
rect 11882 22176 11888 22188
rect 11940 22176 11946 22228
rect 14366 22176 14372 22228
rect 14424 22216 14430 22228
rect 15105 22219 15163 22225
rect 15105 22216 15117 22219
rect 14424 22188 15117 22216
rect 14424 22176 14430 22188
rect 15105 22185 15117 22188
rect 15151 22185 15163 22219
rect 15105 22179 15163 22185
rect 16393 22219 16451 22225
rect 16393 22185 16405 22219
rect 16439 22216 16451 22219
rect 16482 22216 16488 22228
rect 16439 22188 16488 22216
rect 16439 22185 16451 22188
rect 16393 22179 16451 22185
rect 16482 22176 16488 22188
rect 16540 22176 16546 22228
rect 19794 22176 19800 22228
rect 19852 22216 19858 22228
rect 20438 22216 20444 22228
rect 19852 22188 20444 22216
rect 19852 22176 19858 22188
rect 20438 22176 20444 22188
rect 20496 22216 20502 22228
rect 20714 22216 20720 22228
rect 20496 22188 20720 22216
rect 20496 22176 20502 22188
rect 20714 22176 20720 22188
rect 20772 22216 20778 22228
rect 21818 22216 21824 22228
rect 20772 22188 21824 22216
rect 20772 22176 20778 22188
rect 21818 22176 21824 22188
rect 21876 22176 21882 22228
rect 22186 22216 22192 22228
rect 22066 22188 22192 22216
rect 9306 22148 9312 22160
rect 4632 22120 9312 22148
rect 4632 22092 4660 22120
rect 9306 22108 9312 22120
rect 9364 22108 9370 22160
rect 15304 22120 15884 22148
rect 4614 22080 4620 22092
rect 4527 22052 4620 22080
rect 4614 22040 4620 22052
rect 4672 22040 4678 22092
rect 15194 22080 15200 22092
rect 7576 22052 8294 22080
rect 4433 22015 4491 22021
rect 4433 21981 4445 22015
rect 4479 22012 4491 22015
rect 4706 22012 4712 22024
rect 4479 21984 4712 22012
rect 4479 21981 4491 21984
rect 4433 21975 4491 21981
rect 4706 21972 4712 21984
rect 4764 21972 4770 22024
rect 7098 21972 7104 22024
rect 7156 22012 7162 22024
rect 7466 22012 7472 22024
rect 7156 21984 7472 22012
rect 7156 21972 7162 21984
rect 7466 21972 7472 21984
rect 7524 21972 7530 22024
rect 7576 22021 7604 22052
rect 7944 22024 7972 22052
rect 7561 22015 7619 22021
rect 7561 21981 7573 22015
rect 7607 21981 7619 22015
rect 7561 21975 7619 21981
rect 7653 22015 7711 22021
rect 7653 21981 7665 22015
rect 7699 21981 7711 22015
rect 7834 22012 7840 22024
rect 7795 21984 7840 22012
rect 7653 21975 7711 21981
rect 6730 21904 6736 21956
rect 6788 21944 6794 21956
rect 7190 21944 7196 21956
rect 6788 21916 7196 21944
rect 6788 21904 6794 21916
rect 7190 21904 7196 21916
rect 7248 21944 7254 21956
rect 7668 21944 7696 21975
rect 7834 21972 7840 21984
rect 7892 21972 7898 22024
rect 7926 21972 7932 22024
rect 7984 21972 7990 22024
rect 8266 22012 8294 22052
rect 14292 22052 15200 22080
rect 8386 22012 8392 22024
rect 8266 21984 8392 22012
rect 8386 21972 8392 21984
rect 8444 22012 8450 22024
rect 9214 22012 9220 22024
rect 8444 21984 9220 22012
rect 8444 21972 8450 21984
rect 9214 21972 9220 21984
rect 9272 21972 9278 22024
rect 9309 22015 9367 22021
rect 9309 21981 9321 22015
rect 9355 21981 9367 22015
rect 9309 21975 9367 21981
rect 10505 22015 10563 22021
rect 10505 21981 10517 22015
rect 10551 22012 10563 22015
rect 12158 22012 12164 22024
rect 10551 21984 12164 22012
rect 10551 21981 10563 21984
rect 10505 21975 10563 21981
rect 7248 21916 7696 21944
rect 7852 21944 7880 21972
rect 9324 21944 9352 21975
rect 12158 21972 12164 21984
rect 12216 22012 12222 22024
rect 14292 22021 14320 22052
rect 15194 22040 15200 22052
rect 15252 22040 15258 22092
rect 12345 22015 12403 22021
rect 12345 22012 12357 22015
rect 12216 21984 12357 22012
rect 12216 21972 12222 21984
rect 12345 21981 12357 21984
rect 12391 21981 12403 22015
rect 12345 21975 12403 21981
rect 14277 22015 14335 22021
rect 14277 21981 14289 22015
rect 14323 21981 14335 22015
rect 14458 22012 14464 22024
rect 14419 21984 14464 22012
rect 14277 21975 14335 21981
rect 14458 21972 14464 21984
rect 14516 21972 14522 22024
rect 15304 22021 15332 22120
rect 15378 22040 15384 22092
rect 15436 22080 15442 22092
rect 15749 22083 15807 22089
rect 15749 22080 15761 22083
rect 15436 22052 15761 22080
rect 15436 22040 15442 22052
rect 15749 22049 15761 22052
rect 15795 22049 15807 22083
rect 15856 22080 15884 22120
rect 15930 22108 15936 22160
rect 15988 22148 15994 22160
rect 17402 22148 17408 22160
rect 15988 22120 17408 22148
rect 15988 22108 15994 22120
rect 17402 22108 17408 22120
rect 17460 22148 17466 22160
rect 22066 22148 22094 22188
rect 22186 22176 22192 22188
rect 22244 22216 22250 22228
rect 22462 22216 22468 22228
rect 22244 22188 22468 22216
rect 22244 22176 22250 22188
rect 22462 22176 22468 22188
rect 22520 22176 22526 22228
rect 27614 22176 27620 22228
rect 27672 22216 27678 22228
rect 27893 22219 27951 22225
rect 27893 22216 27905 22219
rect 27672 22188 27905 22216
rect 27672 22176 27678 22188
rect 27893 22185 27905 22188
rect 27939 22185 27951 22219
rect 27893 22179 27951 22185
rect 31202 22176 31208 22228
rect 31260 22216 31266 22228
rect 33042 22216 33048 22228
rect 31260 22188 33048 22216
rect 31260 22176 31266 22188
rect 33042 22176 33048 22188
rect 33100 22176 33106 22228
rect 35526 22216 35532 22228
rect 34532 22188 35532 22216
rect 17460 22120 22094 22148
rect 23293 22151 23351 22157
rect 17460 22108 17466 22120
rect 23293 22117 23305 22151
rect 23339 22148 23351 22151
rect 24302 22148 24308 22160
rect 23339 22120 24308 22148
rect 23339 22117 23351 22120
rect 23293 22111 23351 22117
rect 24302 22108 24308 22120
rect 24360 22108 24366 22160
rect 26050 22148 26056 22160
rect 24412 22120 26056 22148
rect 16574 22080 16580 22092
rect 15856 22052 16580 22080
rect 15749 22043 15807 22049
rect 16574 22040 16580 22052
rect 16632 22040 16638 22092
rect 23014 22080 23020 22092
rect 22975 22052 23020 22080
rect 23014 22040 23020 22052
rect 23072 22040 23078 22092
rect 24412 22080 24440 22120
rect 26050 22108 26056 22120
rect 26108 22108 26114 22160
rect 27706 22108 27712 22160
rect 27764 22148 27770 22160
rect 31754 22148 31760 22160
rect 27764 22120 28994 22148
rect 27764 22108 27770 22120
rect 25774 22080 25780 22092
rect 23860 22052 24440 22080
rect 24872 22052 25452 22080
rect 25735 22052 25780 22080
rect 15289 22015 15347 22021
rect 15289 21981 15301 22015
rect 15335 21981 15347 22015
rect 15470 22012 15476 22024
rect 15431 21984 15476 22012
rect 15289 21975 15347 21981
rect 15470 21972 15476 21984
rect 15528 21972 15534 22024
rect 16206 22012 16212 22024
rect 16167 21984 16212 22012
rect 16206 21972 16212 21984
rect 16264 21972 16270 22024
rect 16393 22015 16451 22021
rect 16393 21981 16405 22015
rect 16439 22012 16451 22015
rect 16758 22012 16764 22024
rect 16439 21984 16764 22012
rect 16439 21981 16451 21984
rect 16393 21975 16451 21981
rect 16758 21972 16764 21984
rect 16816 21972 16822 22024
rect 22922 22012 22928 22024
rect 22883 21984 22928 22012
rect 22922 21972 22928 21984
rect 22980 21972 22986 22024
rect 23860 22021 23888 22052
rect 23845 22015 23903 22021
rect 23845 21981 23857 22015
rect 23891 21981 23903 22015
rect 23845 21975 23903 21981
rect 24029 22015 24087 22021
rect 24029 21981 24041 22015
rect 24075 22012 24087 22015
rect 24118 22012 24124 22024
rect 24075 21984 24124 22012
rect 24075 21981 24087 21984
rect 24029 21975 24087 21981
rect 24118 21972 24124 21984
rect 24176 21972 24182 22024
rect 24872 22021 24900 22052
rect 24857 22015 24915 22021
rect 24857 21981 24869 22015
rect 24903 21981 24915 22015
rect 24857 21975 24915 21981
rect 24946 21972 24952 22024
rect 25004 22012 25010 22024
rect 25130 22012 25136 22024
rect 25004 21984 25136 22012
rect 25004 21972 25010 21984
rect 25130 21972 25136 21984
rect 25188 21972 25194 22024
rect 25222 21972 25228 22024
rect 25280 22012 25286 22024
rect 25317 22015 25375 22021
rect 25317 22012 25329 22015
rect 25280 21984 25329 22012
rect 25280 21972 25286 21984
rect 25317 21981 25329 21984
rect 25363 21981 25375 22015
rect 25424 22012 25452 22052
rect 25774 22040 25780 22052
rect 25832 22040 25838 22092
rect 28534 22080 28540 22092
rect 26528 22052 28540 22080
rect 26528 22012 26556 22052
rect 28534 22040 28540 22052
rect 28592 22040 28598 22092
rect 28810 22040 28816 22092
rect 28868 22080 28874 22092
rect 28966 22080 28994 22120
rect 31220 22120 31760 22148
rect 28868 22052 28994 22080
rect 28868 22040 28874 22052
rect 29454 22040 29460 22092
rect 29512 22080 29518 22092
rect 31220 22089 31248 22120
rect 31754 22108 31760 22120
rect 31812 22108 31818 22160
rect 32674 22148 32680 22160
rect 32600 22120 32680 22148
rect 31205 22083 31263 22089
rect 31205 22080 31217 22083
rect 29512 22052 31217 22080
rect 29512 22040 29518 22052
rect 31205 22049 31217 22052
rect 31251 22049 31263 22083
rect 31205 22043 31263 22049
rect 31294 22040 31300 22092
rect 31352 22080 31358 22092
rect 31352 22052 31397 22080
rect 31352 22040 31358 22052
rect 26786 22012 26792 22024
rect 25424 21984 26556 22012
rect 26747 21984 26792 22012
rect 25317 21975 25375 21981
rect 26786 21972 26792 21984
rect 26844 21972 26850 22024
rect 27157 22015 27215 22021
rect 27157 21981 27169 22015
rect 27203 22012 27215 22015
rect 27706 22012 27712 22024
rect 27203 21984 27712 22012
rect 27203 21981 27215 21984
rect 27157 21975 27215 21981
rect 27706 21972 27712 21984
rect 27764 21972 27770 22024
rect 27890 22012 27896 22024
rect 27851 21984 27896 22012
rect 27890 21972 27896 21984
rect 27948 21972 27954 22024
rect 27982 21972 27988 22024
rect 28040 22012 28046 22024
rect 28077 22015 28135 22021
rect 28077 22012 28089 22015
rect 28040 21984 28089 22012
rect 28040 21972 28046 21984
rect 28077 21981 28089 21984
rect 28123 22012 28135 22015
rect 28350 22012 28356 22024
rect 28123 21984 28356 22012
rect 28123 21981 28135 21984
rect 28077 21975 28135 21981
rect 28350 21972 28356 21984
rect 28408 21972 28414 22024
rect 28442 21972 28448 22024
rect 28500 22012 28506 22024
rect 30837 22015 30895 22021
rect 30837 22012 30849 22015
rect 28500 21984 30849 22012
rect 28500 21972 28506 21984
rect 30837 21981 30849 21984
rect 30883 21981 30895 22015
rect 30837 21975 30895 21981
rect 30926 21972 30932 22024
rect 30984 22012 30990 22024
rect 31110 22012 31116 22024
rect 30984 21984 31116 22012
rect 30984 21972 30990 21984
rect 31110 21972 31116 21984
rect 31168 21972 31174 22024
rect 32490 21972 32496 22024
rect 32548 22012 32554 22024
rect 32600 22021 32628 22120
rect 32674 22108 32680 22120
rect 32732 22108 32738 22160
rect 33134 22108 33140 22160
rect 33192 22148 33198 22160
rect 34532 22148 34560 22188
rect 35526 22176 35532 22188
rect 35584 22176 35590 22228
rect 33192 22120 33824 22148
rect 33192 22108 33198 22120
rect 33686 22080 33692 22092
rect 32968 22052 33692 22080
rect 32585 22015 32643 22021
rect 32585 22012 32597 22015
rect 32548 21984 32597 22012
rect 32548 21972 32554 21984
rect 32585 21981 32597 21984
rect 32631 21981 32643 22015
rect 32585 21975 32643 21981
rect 32733 22015 32791 22021
rect 32733 21981 32745 22015
rect 32779 22012 32791 22015
rect 32968 22012 32996 22052
rect 33686 22040 33692 22052
rect 33744 22040 33750 22092
rect 33796 22089 33824 22120
rect 34164 22120 34560 22148
rect 33781 22083 33839 22089
rect 33781 22049 33793 22083
rect 33827 22080 33839 22083
rect 33827 22052 33861 22080
rect 33827 22049 33839 22052
rect 33781 22043 33839 22049
rect 32779 21984 32996 22012
rect 32779 21981 32791 21984
rect 32733 21975 32791 21981
rect 33042 21972 33048 22024
rect 33100 22021 33106 22024
rect 33100 22012 33108 22021
rect 33873 22015 33931 22021
rect 33100 21984 33145 22012
rect 33100 21975 33108 21984
rect 33873 21981 33885 22015
rect 33919 22012 33931 22015
rect 33962 22012 33968 22024
rect 33919 21984 33968 22012
rect 33919 21981 33931 21984
rect 33873 21975 33931 21981
rect 33100 21972 33106 21975
rect 33962 21972 33968 21984
rect 34020 21972 34026 22024
rect 34164 22012 34192 22120
rect 34241 22083 34299 22089
rect 34241 22049 34253 22083
rect 34287 22080 34299 22083
rect 34287 22052 34836 22080
rect 34287 22049 34299 22052
rect 34241 22043 34299 22049
rect 34072 21984 34192 22012
rect 7852 21916 9352 21944
rect 9493 21947 9551 21953
rect 7248 21904 7254 21916
rect 9493 21913 9505 21947
rect 9539 21944 9551 21947
rect 9674 21944 9680 21956
rect 9539 21916 9680 21944
rect 9539 21913 9551 21916
rect 9493 21907 9551 21913
rect 9674 21904 9680 21916
rect 9732 21944 9738 21956
rect 10042 21944 10048 21956
rect 9732 21916 10048 21944
rect 9732 21904 9738 21916
rect 10042 21904 10048 21916
rect 10100 21904 10106 21956
rect 10594 21904 10600 21956
rect 10652 21944 10658 21956
rect 10750 21947 10808 21953
rect 10750 21944 10762 21947
rect 10652 21916 10762 21944
rect 10652 21904 10658 21916
rect 10750 21913 10762 21916
rect 10796 21913 10808 21947
rect 12590 21947 12648 21953
rect 12590 21944 12602 21947
rect 10750 21907 10808 21913
rect 12406 21916 12602 21944
rect 3970 21876 3976 21888
rect 3931 21848 3976 21876
rect 3970 21836 3976 21848
rect 4028 21836 4034 21888
rect 4338 21876 4344 21888
rect 4299 21848 4344 21876
rect 4338 21836 4344 21848
rect 4396 21836 4402 21888
rect 6638 21836 6644 21888
rect 6696 21876 6702 21888
rect 7558 21876 7564 21888
rect 6696 21848 7564 21876
rect 6696 21836 6702 21848
rect 7558 21836 7564 21848
rect 7616 21836 7622 21888
rect 8570 21836 8576 21888
rect 8628 21876 8634 21888
rect 12406 21876 12434 21916
rect 12590 21913 12602 21916
rect 12636 21913 12648 21947
rect 14642 21944 14648 21956
rect 14603 21916 14648 21944
rect 12590 21907 12648 21913
rect 14642 21904 14648 21916
rect 14700 21904 14706 21956
rect 15381 21947 15439 21953
rect 15381 21913 15393 21947
rect 15427 21913 15439 21947
rect 15381 21907 15439 21913
rect 15611 21947 15669 21953
rect 15611 21913 15623 21947
rect 15657 21944 15669 21947
rect 15930 21944 15936 21956
rect 15657 21916 15936 21944
rect 15657 21913 15669 21916
rect 15611 21907 15669 21913
rect 13722 21876 13728 21888
rect 8628 21848 12434 21876
rect 13683 21848 13728 21876
rect 8628 21836 8634 21848
rect 13722 21836 13728 21848
rect 13780 21836 13786 21888
rect 15396 21876 15424 21907
rect 15930 21904 15936 21916
rect 15988 21904 15994 21956
rect 17218 21904 17224 21956
rect 17276 21944 17282 21956
rect 26694 21944 26700 21956
rect 17276 21916 26700 21944
rect 17276 21904 17282 21916
rect 26694 21904 26700 21916
rect 26752 21904 26758 21956
rect 26973 21947 27031 21953
rect 26973 21913 26985 21947
rect 27019 21913 27031 21947
rect 26973 21907 27031 21913
rect 16022 21876 16028 21888
rect 15396 21848 16028 21876
rect 16022 21836 16028 21848
rect 16080 21836 16086 21888
rect 16574 21876 16580 21888
rect 16535 21848 16580 21876
rect 16574 21836 16580 21848
rect 16632 21836 16638 21888
rect 23937 21879 23995 21885
rect 23937 21845 23949 21879
rect 23983 21876 23995 21879
rect 24670 21876 24676 21888
rect 23983 21848 24676 21876
rect 23983 21845 23995 21848
rect 23937 21839 23995 21845
rect 24670 21836 24676 21848
rect 24728 21836 24734 21888
rect 24857 21879 24915 21885
rect 24857 21845 24869 21879
rect 24903 21876 24915 21879
rect 24946 21876 24952 21888
rect 24903 21848 24952 21876
rect 24903 21845 24915 21848
rect 24857 21839 24915 21845
rect 24946 21836 24952 21848
rect 25004 21836 25010 21888
rect 25774 21836 25780 21888
rect 25832 21876 25838 21888
rect 26988 21876 27016 21907
rect 27062 21904 27068 21956
rect 27120 21944 27126 21956
rect 32122 21944 32128 21956
rect 27120 21916 32128 21944
rect 27120 21904 27126 21916
rect 32122 21904 32128 21916
rect 32180 21904 32186 21956
rect 32858 21944 32864 21956
rect 32819 21916 32864 21944
rect 32858 21904 32864 21916
rect 32916 21904 32922 21956
rect 32953 21947 33011 21953
rect 32953 21913 32965 21947
rect 32999 21944 33011 21947
rect 34072 21944 34100 21984
rect 32999 21916 34100 21944
rect 34808 21944 34836 22052
rect 34885 22015 34943 22021
rect 34885 21981 34897 22015
rect 34931 22012 34943 22015
rect 36814 22012 36820 22024
rect 34931 21984 36820 22012
rect 34931 21981 34943 21984
rect 34885 21975 34943 21981
rect 36814 21972 36820 21984
rect 36872 22012 36878 22024
rect 36909 22015 36967 22021
rect 36909 22012 36921 22015
rect 36872 21984 36921 22012
rect 36872 21972 36878 21984
rect 36909 21981 36921 21984
rect 36955 21981 36967 22015
rect 36909 21975 36967 21981
rect 35130 21947 35188 21953
rect 35130 21944 35142 21947
rect 34808 21916 35142 21944
rect 32999 21913 33011 21916
rect 32953 21907 33011 21913
rect 35130 21913 35142 21916
rect 35176 21913 35188 21947
rect 35130 21907 35188 21913
rect 37176 21947 37234 21953
rect 37176 21913 37188 21947
rect 37222 21944 37234 21947
rect 37458 21944 37464 21956
rect 37222 21916 37464 21944
rect 37222 21913 37234 21916
rect 37176 21907 37234 21913
rect 27246 21876 27252 21888
rect 25832 21848 27252 21876
rect 25832 21836 25838 21848
rect 27246 21836 27252 21848
rect 27304 21836 27310 21888
rect 27341 21879 27399 21885
rect 27341 21845 27353 21879
rect 27387 21876 27399 21879
rect 27522 21876 27528 21888
rect 27387 21848 27528 21876
rect 27387 21845 27399 21848
rect 27341 21839 27399 21845
rect 27522 21836 27528 21848
rect 27580 21836 27586 21888
rect 27982 21836 27988 21888
rect 28040 21876 28046 21888
rect 28626 21876 28632 21888
rect 28040 21848 28632 21876
rect 28040 21836 28046 21848
rect 28626 21836 28632 21848
rect 28684 21836 28690 21888
rect 30650 21876 30656 21888
rect 30611 21848 30656 21876
rect 30650 21836 30656 21848
rect 30708 21836 30714 21888
rect 31386 21836 31392 21888
rect 31444 21876 31450 21888
rect 31754 21876 31760 21888
rect 31444 21848 31760 21876
rect 31444 21836 31450 21848
rect 31754 21836 31760 21848
rect 31812 21836 31818 21888
rect 32214 21836 32220 21888
rect 32272 21876 32278 21888
rect 32968 21876 32996 21907
rect 37458 21904 37464 21916
rect 37516 21904 37522 21956
rect 33226 21876 33232 21888
rect 32272 21848 32996 21876
rect 33187 21848 33232 21876
rect 32272 21836 32278 21848
rect 33226 21836 33232 21848
rect 33284 21836 33290 21888
rect 35526 21836 35532 21888
rect 35584 21876 35590 21888
rect 36265 21879 36323 21885
rect 36265 21876 36277 21879
rect 35584 21848 36277 21876
rect 35584 21836 35590 21848
rect 36265 21845 36277 21848
rect 36311 21876 36323 21879
rect 36630 21876 36636 21888
rect 36311 21848 36636 21876
rect 36311 21845 36323 21848
rect 36265 21839 36323 21845
rect 36630 21836 36636 21848
rect 36688 21836 36694 21888
rect 38286 21876 38292 21888
rect 38247 21848 38292 21876
rect 38286 21836 38292 21848
rect 38344 21836 38350 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 5902 21632 5908 21684
rect 5960 21672 5966 21684
rect 5960 21644 6868 21672
rect 5960 21632 5966 21644
rect 3044 21607 3102 21613
rect 3044 21573 3056 21607
rect 3090 21604 3102 21607
rect 3970 21604 3976 21616
rect 3090 21576 3976 21604
rect 3090 21573 3102 21576
rect 3044 21567 3102 21573
rect 3970 21564 3976 21576
rect 4028 21564 4034 21616
rect 6638 21604 6644 21616
rect 6564 21576 6644 21604
rect 2774 21496 2780 21548
rect 2832 21536 2838 21548
rect 5721 21539 5779 21545
rect 2832 21508 2877 21536
rect 2832 21496 2838 21508
rect 5721 21505 5733 21539
rect 5767 21536 5779 21539
rect 5810 21536 5816 21548
rect 5767 21508 5816 21536
rect 5767 21505 5779 21508
rect 5721 21499 5779 21505
rect 5810 21496 5816 21508
rect 5868 21496 5874 21548
rect 6564 21545 6592 21576
rect 6638 21564 6644 21576
rect 6696 21564 6702 21616
rect 6840 21613 6868 21644
rect 7466 21632 7472 21684
rect 7524 21672 7530 21684
rect 9243 21675 9301 21681
rect 7524 21644 9168 21672
rect 7524 21632 7530 21644
rect 6825 21607 6883 21613
rect 6825 21573 6837 21607
rect 6871 21573 6883 21607
rect 6825 21567 6883 21573
rect 9033 21607 9091 21613
rect 9033 21573 9045 21607
rect 9079 21573 9091 21607
rect 9140 21604 9168 21644
rect 9243 21641 9255 21675
rect 9289 21672 9301 21675
rect 9398 21672 9404 21684
rect 9289 21644 9404 21672
rect 9289 21641 9301 21644
rect 9243 21635 9301 21641
rect 9398 21632 9404 21644
rect 9456 21672 9462 21684
rect 9861 21675 9919 21681
rect 9861 21672 9873 21675
rect 9456 21644 9873 21672
rect 9456 21632 9462 21644
rect 9861 21641 9873 21644
rect 9907 21641 9919 21675
rect 9861 21635 9919 21641
rect 12434 21632 12440 21684
rect 12492 21672 12498 21684
rect 22094 21672 22100 21684
rect 12492 21644 15884 21672
rect 22007 21644 22100 21672
rect 12492 21632 12498 21644
rect 10137 21607 10195 21613
rect 10137 21604 10149 21607
rect 9140 21576 10149 21604
rect 9033 21567 9091 21573
rect 10137 21573 10149 21576
rect 10183 21573 10195 21607
rect 10137 21567 10195 21573
rect 6549 21539 6607 21545
rect 6549 21505 6561 21539
rect 6595 21505 6607 21539
rect 6730 21536 6736 21548
rect 6691 21508 6736 21536
rect 6549 21499 6607 21505
rect 6730 21496 6736 21508
rect 6788 21496 6794 21548
rect 6914 21496 6920 21548
rect 6972 21536 6978 21548
rect 7837 21539 7895 21545
rect 6972 21508 7017 21536
rect 6972 21496 6978 21508
rect 7837 21505 7849 21539
rect 7883 21536 7895 21539
rect 8202 21536 8208 21548
rect 7883 21508 8208 21536
rect 7883 21505 7895 21508
rect 7837 21499 7895 21505
rect 8202 21496 8208 21508
rect 8260 21496 8266 21548
rect 4614 21428 4620 21480
rect 4672 21468 4678 21480
rect 5537 21471 5595 21477
rect 5537 21468 5549 21471
rect 4672 21440 5549 21468
rect 4672 21428 4678 21440
rect 5537 21437 5549 21440
rect 5583 21437 5595 21471
rect 5537 21431 5595 21437
rect 5905 21471 5963 21477
rect 5905 21437 5917 21471
rect 5951 21468 5963 21471
rect 6748 21468 6776 21496
rect 7926 21468 7932 21480
rect 5951 21440 6776 21468
rect 7887 21440 7932 21468
rect 5951 21437 5963 21440
rect 5905 21431 5963 21437
rect 7926 21428 7932 21440
rect 7984 21428 7990 21480
rect 8021 21471 8079 21477
rect 8021 21437 8033 21471
rect 8067 21437 8079 21471
rect 8021 21431 8079 21437
rect 4157 21403 4215 21409
rect 4157 21369 4169 21403
rect 4203 21400 4215 21403
rect 4338 21400 4344 21412
rect 4203 21372 4344 21400
rect 4203 21369 4215 21372
rect 4157 21363 4215 21369
rect 4338 21360 4344 21372
rect 4396 21400 4402 21412
rect 4396 21372 7788 21400
rect 4396 21360 4402 21372
rect 5994 21292 6000 21344
rect 6052 21332 6058 21344
rect 7101 21335 7159 21341
rect 7101 21332 7113 21335
rect 6052 21304 7113 21332
rect 6052 21292 6058 21304
rect 7101 21301 7113 21304
rect 7147 21301 7159 21335
rect 7650 21332 7656 21344
rect 7611 21304 7656 21332
rect 7101 21295 7159 21301
rect 7650 21292 7656 21304
rect 7708 21292 7714 21344
rect 7760 21332 7788 21372
rect 7834 21360 7840 21412
rect 7892 21400 7898 21412
rect 8036 21400 8064 21431
rect 8110 21428 8116 21480
rect 8168 21468 8174 21480
rect 8168 21440 8213 21468
rect 8168 21428 8174 21440
rect 9048 21400 9076 21567
rect 11882 21564 11888 21616
rect 11940 21604 11946 21616
rect 15746 21604 15752 21616
rect 11940 21576 15752 21604
rect 11940 21564 11946 21576
rect 15746 21564 15752 21576
rect 15804 21564 15810 21616
rect 9766 21496 9772 21548
rect 9824 21536 9830 21548
rect 9861 21539 9919 21545
rect 9861 21536 9873 21539
rect 9824 21508 9873 21536
rect 9824 21496 9830 21508
rect 9861 21505 9873 21508
rect 9907 21505 9919 21539
rect 9861 21499 9919 21505
rect 13814 21496 13820 21548
rect 13872 21536 13878 21548
rect 14737 21539 14795 21545
rect 14737 21536 14749 21539
rect 13872 21508 14749 21536
rect 13872 21496 13878 21508
rect 14737 21505 14749 21508
rect 14783 21505 14795 21539
rect 14737 21499 14795 21505
rect 15013 21539 15071 21545
rect 15013 21505 15025 21539
rect 15059 21536 15071 21539
rect 15654 21536 15660 21548
rect 15059 21508 15660 21536
rect 15059 21505 15071 21508
rect 15013 21499 15071 21505
rect 15654 21496 15660 21508
rect 15712 21496 15718 21548
rect 9214 21428 9220 21480
rect 9272 21468 9278 21480
rect 9953 21471 10011 21477
rect 9953 21468 9965 21471
rect 9272 21440 9965 21468
rect 9272 21428 9278 21440
rect 9953 21437 9965 21440
rect 9999 21437 10011 21471
rect 9953 21431 10011 21437
rect 11882 21428 11888 21480
rect 11940 21468 11946 21480
rect 14550 21468 14556 21480
rect 11940 21440 14556 21468
rect 11940 21428 11946 21440
rect 14550 21428 14556 21440
rect 14608 21428 14614 21480
rect 14918 21468 14924 21480
rect 14879 21440 14924 21468
rect 14918 21428 14924 21440
rect 14976 21428 14982 21480
rect 15764 21468 15792 21564
rect 15856 21545 15884 21644
rect 16942 21564 16948 21616
rect 17000 21604 17006 21616
rect 17000 21576 19564 21604
rect 17000 21564 17006 21576
rect 15841 21539 15899 21545
rect 15841 21505 15853 21539
rect 15887 21505 15899 21539
rect 15841 21499 15899 21505
rect 15933 21539 15991 21545
rect 15933 21505 15945 21539
rect 15979 21536 15991 21539
rect 16666 21536 16672 21548
rect 15979 21508 16672 21536
rect 15979 21505 15991 21508
rect 15933 21499 15991 21505
rect 16666 21496 16672 21508
rect 16724 21496 16730 21548
rect 16853 21539 16911 21545
rect 16853 21505 16865 21539
rect 16899 21536 16911 21539
rect 19426 21536 19432 21548
rect 16899 21508 19432 21536
rect 16899 21505 16911 21508
rect 16853 21499 16911 21505
rect 19426 21496 19432 21508
rect 19484 21496 19490 21548
rect 16206 21468 16212 21480
rect 15764 21440 16212 21468
rect 16206 21428 16212 21440
rect 16264 21428 16270 21480
rect 16301 21471 16359 21477
rect 16301 21437 16313 21471
rect 16347 21468 16359 21471
rect 17589 21471 17647 21477
rect 17589 21468 17601 21471
rect 16347 21440 17601 21468
rect 16347 21437 16359 21440
rect 16301 21431 16359 21437
rect 17589 21437 17601 21440
rect 17635 21468 17647 21471
rect 18414 21468 18420 21480
rect 17635 21440 18420 21468
rect 17635 21437 17647 21440
rect 17589 21431 17647 21437
rect 18414 21428 18420 21440
rect 18472 21428 18478 21480
rect 19536 21468 19564 21576
rect 22020 21545 22048 21644
rect 22094 21632 22100 21644
rect 22152 21672 22158 21684
rect 24578 21672 24584 21684
rect 22152 21644 24584 21672
rect 22152 21632 22158 21644
rect 24578 21632 24584 21644
rect 24636 21632 24642 21684
rect 26513 21675 26571 21681
rect 26513 21641 26525 21675
rect 26559 21672 26571 21675
rect 26878 21672 26884 21684
rect 26559 21644 26884 21672
rect 26559 21641 26571 21644
rect 26513 21635 26571 21641
rect 26878 21632 26884 21644
rect 26936 21632 26942 21684
rect 27246 21632 27252 21684
rect 27304 21672 27310 21684
rect 32861 21675 32919 21681
rect 32861 21672 32873 21675
rect 27304 21644 27568 21672
rect 27304 21632 27310 21644
rect 22281 21607 22339 21613
rect 22281 21573 22293 21607
rect 22327 21604 22339 21607
rect 27062 21604 27068 21616
rect 22327 21576 27068 21604
rect 22327 21573 22339 21576
rect 22281 21567 22339 21573
rect 27062 21564 27068 21576
rect 27120 21564 27126 21616
rect 27430 21604 27436 21616
rect 27391 21576 27436 21604
rect 27430 21564 27436 21576
rect 27488 21564 27494 21616
rect 27540 21604 27568 21644
rect 28736 21644 32873 21672
rect 27614 21604 27620 21616
rect 27540 21576 27620 21604
rect 22005 21539 22063 21545
rect 22005 21505 22017 21539
rect 22051 21505 22063 21539
rect 22186 21536 22192 21548
rect 22147 21508 22192 21536
rect 22005 21499 22063 21505
rect 22186 21496 22192 21508
rect 22244 21496 22250 21548
rect 22370 21496 22376 21548
rect 22428 21545 22434 21548
rect 22428 21536 22436 21545
rect 22428 21508 22473 21536
rect 22428 21499 22436 21508
rect 22428 21496 22434 21499
rect 24670 21496 24676 21548
rect 24728 21536 24734 21548
rect 24765 21539 24823 21545
rect 24765 21536 24777 21539
rect 24728 21508 24777 21536
rect 24728 21496 24734 21508
rect 24765 21505 24777 21508
rect 24811 21505 24823 21539
rect 26326 21536 26332 21548
rect 26287 21508 26332 21536
rect 24765 21499 24823 21505
rect 26326 21496 26332 21508
rect 26384 21496 26390 21548
rect 26602 21536 26608 21548
rect 26563 21508 26608 21536
rect 26602 21496 26608 21508
rect 26660 21496 26666 21548
rect 26694 21496 26700 21548
rect 26752 21536 26758 21548
rect 27540 21545 27568 21576
rect 27614 21564 27620 21576
rect 27672 21604 27678 21616
rect 28626 21604 28632 21616
rect 27672 21576 28632 21604
rect 27672 21564 27678 21576
rect 28626 21564 28632 21576
rect 28684 21564 28690 21616
rect 28534 21545 28540 21548
rect 27157 21539 27215 21545
rect 27157 21536 27169 21539
rect 26752 21508 27169 21536
rect 26752 21496 26758 21508
rect 27157 21505 27169 21508
rect 27203 21505 27215 21539
rect 27157 21499 27215 21505
rect 27341 21539 27399 21545
rect 27341 21505 27353 21539
rect 27387 21505 27399 21539
rect 27341 21499 27399 21505
rect 27525 21539 27583 21545
rect 27525 21505 27537 21539
rect 27571 21505 27583 21539
rect 27525 21499 27583 21505
rect 28353 21539 28411 21545
rect 28353 21505 28365 21539
rect 28399 21505 28411 21539
rect 28353 21499 28411 21505
rect 28501 21539 28540 21545
rect 28501 21505 28513 21539
rect 28501 21499 28540 21505
rect 26145 21471 26203 21477
rect 19536 21440 22094 21468
rect 7892 21372 9076 21400
rect 9140 21372 9812 21400
rect 7892 21360 7898 21372
rect 9140 21332 9168 21372
rect 7760 21304 9168 21332
rect 9214 21292 9220 21344
rect 9272 21332 9278 21344
rect 9401 21335 9459 21341
rect 9272 21304 9317 21332
rect 9272 21292 9278 21304
rect 9401 21301 9413 21335
rect 9447 21332 9459 21335
rect 9582 21332 9588 21344
rect 9447 21304 9588 21332
rect 9447 21301 9459 21304
rect 9401 21295 9459 21301
rect 9582 21292 9588 21304
rect 9640 21292 9646 21344
rect 9784 21332 9812 21372
rect 10962 21360 10968 21412
rect 11020 21400 11026 21412
rect 13538 21400 13544 21412
rect 11020 21372 13544 21400
rect 11020 21360 11026 21372
rect 13538 21360 13544 21372
rect 13596 21360 13602 21412
rect 13630 21360 13636 21412
rect 13688 21400 13694 21412
rect 21818 21400 21824 21412
rect 13688 21372 21824 21400
rect 13688 21360 13694 21372
rect 21818 21360 21824 21372
rect 21876 21360 21882 21412
rect 22066 21400 22094 21440
rect 26145 21437 26157 21471
rect 26191 21468 26203 21471
rect 27246 21468 27252 21480
rect 26191 21440 27252 21468
rect 26191 21437 26203 21440
rect 26145 21431 26203 21437
rect 27246 21428 27252 21440
rect 27304 21468 27310 21480
rect 27356 21468 27384 21499
rect 28368 21468 28396 21499
rect 28534 21496 28540 21499
rect 28592 21496 28598 21548
rect 28736 21545 28764 21644
rect 32861 21641 32873 21644
rect 32907 21672 32919 21675
rect 35526 21672 35532 21684
rect 32907 21644 35532 21672
rect 32907 21641 32919 21644
rect 32861 21635 32919 21641
rect 35526 21632 35532 21644
rect 35584 21632 35590 21684
rect 35621 21675 35679 21681
rect 35621 21641 35633 21675
rect 35667 21641 35679 21675
rect 37458 21672 37464 21684
rect 37419 21644 37464 21672
rect 35621 21635 35679 21641
rect 32490 21604 32496 21616
rect 30484 21576 32496 21604
rect 30484 21548 30512 21576
rect 32490 21564 32496 21576
rect 32548 21564 32554 21616
rect 32677 21607 32735 21613
rect 32677 21573 32689 21607
rect 32723 21604 32735 21607
rect 33226 21604 33232 21616
rect 32723 21576 33232 21604
rect 32723 21573 32735 21576
rect 32677 21567 32735 21573
rect 33226 21564 33232 21576
rect 33284 21564 33290 21616
rect 33686 21564 33692 21616
rect 33744 21604 33750 21616
rect 35345 21607 35403 21613
rect 35345 21604 35357 21607
rect 33744 21576 35357 21604
rect 33744 21564 33750 21576
rect 35345 21573 35357 21576
rect 35391 21573 35403 21607
rect 35345 21567 35403 21573
rect 28721 21539 28779 21545
rect 28721 21505 28733 21539
rect 28767 21505 28779 21539
rect 28721 21499 28779 21505
rect 28818 21539 28876 21545
rect 28818 21505 28830 21539
rect 28864 21505 28876 21539
rect 30466 21536 30472 21548
rect 30379 21508 30472 21536
rect 28818 21499 28876 21505
rect 27304 21440 28396 21468
rect 27304 21428 27310 21440
rect 22557 21403 22615 21409
rect 22557 21400 22569 21403
rect 22066 21372 22569 21400
rect 22557 21369 22569 21372
rect 22603 21369 22615 21403
rect 22557 21363 22615 21369
rect 24578 21360 24584 21412
rect 24636 21400 24642 21412
rect 28736 21400 28764 21499
rect 24636 21372 28764 21400
rect 24636 21360 24642 21372
rect 14274 21332 14280 21344
rect 9784 21304 14280 21332
rect 14274 21292 14280 21304
rect 14332 21292 14338 21344
rect 14734 21332 14740 21344
rect 14695 21304 14740 21332
rect 14734 21292 14740 21304
rect 14792 21292 14798 21344
rect 15194 21332 15200 21344
rect 15155 21304 15200 21332
rect 15194 21292 15200 21304
rect 15252 21292 15258 21344
rect 15378 21292 15384 21344
rect 15436 21332 15442 21344
rect 15657 21335 15715 21341
rect 15657 21332 15669 21335
rect 15436 21304 15669 21332
rect 15436 21292 15442 21304
rect 15657 21301 15669 21304
rect 15703 21301 15715 21335
rect 15657 21295 15715 21301
rect 15838 21292 15844 21344
rect 15896 21332 15902 21344
rect 19334 21332 19340 21344
rect 15896 21304 19340 21332
rect 15896 21292 15902 21304
rect 19334 21292 19340 21304
rect 19392 21292 19398 21344
rect 25041 21335 25099 21341
rect 25041 21301 25053 21335
rect 25087 21332 25099 21335
rect 25130 21332 25136 21344
rect 25087 21304 25136 21332
rect 25087 21301 25099 21304
rect 25041 21295 25099 21301
rect 25130 21292 25136 21304
rect 25188 21292 25194 21344
rect 27430 21292 27436 21344
rect 27488 21332 27494 21344
rect 27709 21335 27767 21341
rect 27709 21332 27721 21335
rect 27488 21304 27721 21332
rect 27488 21292 27494 21304
rect 27709 21301 27721 21304
rect 27755 21301 27767 21335
rect 27709 21295 27767 21301
rect 27798 21292 27804 21344
rect 27856 21332 27862 21344
rect 28828 21332 28856 21499
rect 30466 21496 30472 21508
rect 30524 21496 30530 21548
rect 30742 21536 30748 21548
rect 30703 21508 30748 21536
rect 30742 21496 30748 21508
rect 30800 21496 30806 21548
rect 31202 21536 31208 21548
rect 31163 21508 31208 21536
rect 31202 21496 31208 21508
rect 31260 21496 31266 21548
rect 31478 21496 31484 21548
rect 31536 21536 31542 21548
rect 31573 21539 31631 21545
rect 31573 21536 31585 21539
rect 31536 21508 31585 21536
rect 31536 21496 31542 21508
rect 31573 21505 31585 21508
rect 31619 21505 31631 21539
rect 31573 21499 31631 21505
rect 32582 21496 32588 21548
rect 32640 21536 32646 21548
rect 32950 21536 32956 21548
rect 32640 21508 32956 21536
rect 32640 21496 32646 21508
rect 32950 21496 32956 21508
rect 33008 21496 33014 21548
rect 34790 21496 34796 21548
rect 34848 21536 34854 21548
rect 34977 21539 35035 21545
rect 34977 21536 34989 21539
rect 34848 21508 34989 21536
rect 34848 21496 34854 21508
rect 34977 21505 34989 21508
rect 35023 21505 35035 21539
rect 34977 21499 35035 21505
rect 35070 21539 35128 21545
rect 35070 21505 35082 21539
rect 35116 21505 35128 21539
rect 35250 21536 35256 21548
rect 35211 21508 35256 21536
rect 35070 21499 35128 21505
rect 30558 21428 30564 21480
rect 30616 21468 30622 21480
rect 31021 21471 31079 21477
rect 31021 21468 31033 21471
rect 30616 21440 31033 21468
rect 30616 21428 30622 21440
rect 31021 21437 31033 21440
rect 31067 21437 31079 21471
rect 34422 21468 34428 21480
rect 31021 21431 31079 21437
rect 31312 21440 34428 21468
rect 31312 21412 31340 21440
rect 34422 21428 34428 21440
rect 34480 21428 34486 21480
rect 34514 21428 34520 21480
rect 34572 21468 34578 21480
rect 35084 21468 35112 21499
rect 35250 21496 35256 21508
rect 35308 21496 35314 21548
rect 34572 21440 35112 21468
rect 35360 21468 35388 21567
rect 35526 21545 35532 21548
rect 35483 21539 35532 21545
rect 35483 21505 35495 21539
rect 35529 21505 35532 21539
rect 35483 21499 35532 21505
rect 35526 21496 35532 21499
rect 35584 21496 35590 21548
rect 35636 21536 35664 21635
rect 37458 21632 37464 21644
rect 37516 21632 37522 21684
rect 36081 21607 36139 21613
rect 36081 21573 36093 21607
rect 36127 21604 36139 21607
rect 37734 21604 37740 21616
rect 36127 21576 37740 21604
rect 36127 21573 36139 21576
rect 36081 21567 36139 21573
rect 37734 21564 37740 21576
rect 37792 21604 37798 21616
rect 37921 21607 37979 21613
rect 37921 21604 37933 21607
rect 37792 21576 37933 21604
rect 37792 21564 37798 21576
rect 37921 21573 37933 21576
rect 37967 21573 37979 21607
rect 37921 21567 37979 21573
rect 36265 21539 36323 21545
rect 36265 21536 36277 21539
rect 35636 21508 36277 21536
rect 36265 21505 36277 21508
rect 36311 21505 36323 21539
rect 36265 21499 36323 21505
rect 36354 21496 36360 21548
rect 36412 21536 36418 21548
rect 36630 21536 36636 21548
rect 36412 21508 36457 21536
rect 36591 21508 36636 21536
rect 36412 21496 36418 21508
rect 36630 21496 36636 21508
rect 36688 21496 36694 21548
rect 37829 21539 37887 21545
rect 37829 21505 37841 21539
rect 37875 21536 37887 21539
rect 38286 21536 38292 21548
rect 37875 21508 38292 21536
rect 37875 21505 37887 21508
rect 37829 21499 37887 21505
rect 37844 21468 37872 21499
rect 38286 21496 38292 21508
rect 38344 21496 38350 21548
rect 38010 21468 38016 21480
rect 35360 21440 37872 21468
rect 37971 21440 38016 21468
rect 34572 21428 34578 21440
rect 29086 21360 29092 21412
rect 29144 21400 29150 21412
rect 31294 21400 31300 21412
rect 29144 21372 31300 21400
rect 29144 21360 29150 21372
rect 31294 21360 31300 21372
rect 31352 21360 31358 21412
rect 32677 21403 32735 21409
rect 32677 21369 32689 21403
rect 32723 21400 32735 21403
rect 33134 21400 33140 21412
rect 32723 21372 33140 21400
rect 32723 21369 32735 21372
rect 32677 21363 32735 21369
rect 33134 21360 33140 21372
rect 33192 21360 33198 21412
rect 35084 21400 35112 21440
rect 38010 21428 38016 21440
rect 38068 21428 38074 21480
rect 35342 21400 35348 21412
rect 35084 21372 35348 21400
rect 35342 21360 35348 21372
rect 35400 21360 35406 21412
rect 36538 21400 36544 21412
rect 36499 21372 36544 21400
rect 36538 21360 36544 21372
rect 36596 21360 36602 21412
rect 27856 21304 28856 21332
rect 28997 21335 29055 21341
rect 27856 21292 27862 21304
rect 28997 21301 29009 21335
rect 29043 21332 29055 21335
rect 29730 21332 29736 21344
rect 29043 21304 29736 21332
rect 29043 21301 29055 21304
rect 28997 21295 29055 21301
rect 29730 21292 29736 21304
rect 29788 21292 29794 21344
rect 34422 21292 34428 21344
rect 34480 21332 34486 21344
rect 35250 21332 35256 21344
rect 34480 21304 35256 21332
rect 34480 21292 34486 21304
rect 35250 21292 35256 21304
rect 35308 21292 35314 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 5902 21128 5908 21140
rect 5863 21100 5908 21128
rect 5902 21088 5908 21100
rect 5960 21088 5966 21140
rect 9582 21088 9588 21140
rect 9640 21128 9646 21140
rect 10686 21128 10692 21140
rect 9640 21100 10692 21128
rect 9640 21088 9646 21100
rect 10686 21088 10692 21100
rect 10744 21088 10750 21140
rect 10962 21128 10968 21140
rect 10923 21100 10968 21128
rect 10962 21088 10968 21100
rect 11020 21088 11026 21140
rect 14550 21088 14556 21140
rect 14608 21128 14614 21140
rect 15838 21128 15844 21140
rect 14608 21100 15844 21128
rect 14608 21088 14614 21100
rect 15838 21088 15844 21100
rect 15896 21088 15902 21140
rect 18506 21128 18512 21140
rect 18467 21100 18512 21128
rect 18506 21088 18512 21100
rect 18564 21088 18570 21140
rect 21818 21128 21824 21140
rect 21779 21100 21824 21128
rect 21818 21088 21824 21100
rect 21876 21128 21882 21140
rect 25038 21128 25044 21140
rect 21876 21100 25044 21128
rect 21876 21088 21882 21100
rect 25038 21088 25044 21100
rect 25096 21088 25102 21140
rect 25314 21088 25320 21140
rect 25372 21128 25378 21140
rect 25682 21128 25688 21140
rect 25372 21100 25688 21128
rect 25372 21088 25378 21100
rect 25682 21088 25688 21100
rect 25740 21088 25746 21140
rect 26326 21088 26332 21140
rect 26384 21128 26390 21140
rect 30466 21128 30472 21140
rect 26384 21100 30472 21128
rect 26384 21088 26390 21100
rect 30466 21088 30472 21100
rect 30524 21088 30530 21140
rect 31386 21088 31392 21140
rect 31444 21128 31450 21140
rect 31573 21131 31631 21137
rect 31573 21128 31585 21131
rect 31444 21100 31585 21128
rect 31444 21088 31450 21100
rect 31573 21097 31585 21100
rect 31619 21097 31631 21131
rect 31938 21128 31944 21140
rect 31899 21100 31944 21128
rect 31573 21091 31631 21097
rect 31938 21088 31944 21100
rect 31996 21088 32002 21140
rect 13722 21020 13728 21072
rect 13780 21060 13786 21072
rect 13780 21032 17080 21060
rect 13780 21020 13786 21032
rect 2774 20952 2780 21004
rect 2832 20992 2838 21004
rect 3970 20992 3976 21004
rect 2832 20964 3976 20992
rect 2832 20952 2838 20964
rect 3970 20952 3976 20964
rect 4028 20992 4034 21004
rect 4525 20995 4583 21001
rect 4525 20992 4537 20995
rect 4028 20964 4537 20992
rect 4028 20952 4034 20964
rect 4525 20961 4537 20964
rect 4571 20961 4583 20995
rect 9214 20992 9220 21004
rect 4525 20955 4583 20961
rect 7208 20964 9220 20992
rect 7208 20936 7236 20964
rect 9214 20952 9220 20964
rect 9272 20952 9278 21004
rect 14921 20995 14979 21001
rect 14921 20961 14933 20995
rect 14967 20992 14979 20995
rect 15286 20992 15292 21004
rect 14967 20964 15292 20992
rect 14967 20961 14979 20964
rect 14921 20955 14979 20961
rect 15286 20952 15292 20964
rect 15344 20952 15350 21004
rect 16758 20992 16764 21004
rect 15396 20964 16764 20992
rect 4792 20927 4850 20933
rect 4792 20893 4804 20927
rect 4838 20924 4850 20927
rect 5994 20924 6000 20936
rect 4838 20896 6000 20924
rect 4838 20893 4850 20896
rect 4792 20887 4850 20893
rect 5994 20884 6000 20896
rect 6052 20884 6058 20936
rect 6825 20927 6883 20933
rect 6825 20893 6837 20927
rect 6871 20924 6883 20927
rect 7006 20924 7012 20936
rect 6871 20896 7012 20924
rect 6871 20893 6883 20896
rect 6825 20887 6883 20893
rect 7006 20884 7012 20896
rect 7064 20884 7070 20936
rect 7101 20927 7159 20933
rect 7101 20893 7113 20927
rect 7147 20924 7159 20927
rect 7190 20924 7196 20936
rect 7147 20896 7196 20924
rect 7147 20893 7159 20896
rect 7101 20887 7159 20893
rect 7190 20884 7196 20896
rect 7248 20884 7254 20936
rect 9122 20884 9128 20936
rect 9180 20924 9186 20936
rect 9585 20927 9643 20933
rect 9585 20924 9597 20927
rect 9180 20896 9597 20924
rect 9180 20884 9186 20896
rect 9585 20893 9597 20896
rect 9631 20893 9643 20927
rect 9585 20887 9643 20893
rect 13538 20884 13544 20936
rect 13596 20924 13602 20936
rect 15396 20924 15424 20964
rect 16758 20952 16764 20964
rect 16816 20952 16822 21004
rect 17052 20978 17080 21032
rect 28902 21020 28908 21072
rect 28960 21060 28966 21072
rect 30190 21060 30196 21072
rect 28960 21032 30196 21060
rect 28960 21020 28966 21032
rect 30190 21020 30196 21032
rect 30248 21020 30254 21072
rect 32585 21063 32643 21069
rect 32585 21029 32597 21063
rect 32631 21060 32643 21063
rect 33594 21060 33600 21072
rect 32631 21032 33600 21060
rect 32631 21029 32643 21032
rect 32585 21023 32643 21029
rect 33594 21020 33600 21032
rect 33652 21020 33658 21072
rect 24118 20952 24124 21004
rect 24176 20992 24182 21004
rect 24176 20964 24716 20992
rect 24176 20952 24182 20964
rect 13596 20896 15424 20924
rect 15473 20927 15531 20933
rect 13596 20884 13602 20896
rect 15473 20893 15485 20927
rect 15519 20924 15531 20927
rect 15562 20924 15568 20936
rect 15519 20896 15568 20924
rect 15519 20893 15531 20896
rect 15473 20887 15531 20893
rect 15562 20884 15568 20896
rect 15620 20884 15626 20936
rect 17586 20924 17592 20936
rect 15672 20896 17264 20924
rect 17547 20896 17592 20924
rect 9852 20859 9910 20865
rect 9852 20825 9864 20859
rect 9898 20856 9910 20859
rect 9950 20856 9956 20868
rect 9898 20828 9956 20856
rect 9898 20825 9910 20828
rect 9852 20819 9910 20825
rect 9950 20816 9956 20828
rect 10008 20816 10014 20868
rect 13906 20816 13912 20868
rect 13964 20856 13970 20868
rect 14458 20856 14464 20868
rect 13964 20828 14464 20856
rect 13964 20816 13970 20828
rect 14458 20816 14464 20828
rect 14516 20856 14522 20868
rect 14645 20859 14703 20865
rect 14645 20856 14657 20859
rect 14516 20828 14657 20856
rect 14516 20816 14522 20828
rect 14645 20825 14657 20828
rect 14691 20856 14703 20859
rect 15672 20856 15700 20896
rect 17236 20868 17264 20896
rect 17586 20884 17592 20896
rect 17644 20884 17650 20936
rect 20530 20924 20536 20936
rect 20491 20896 20536 20924
rect 20530 20884 20536 20896
rect 20588 20884 20594 20936
rect 24486 20884 24492 20936
rect 24544 20924 24550 20936
rect 24581 20927 24639 20933
rect 24581 20924 24593 20927
rect 24544 20896 24593 20924
rect 24544 20884 24550 20896
rect 24581 20893 24593 20896
rect 24627 20893 24639 20927
rect 24688 20924 24716 20964
rect 24762 20952 24768 21004
rect 24820 20992 24826 21004
rect 24820 20964 27384 20992
rect 24820 20952 24826 20964
rect 24857 20927 24915 20933
rect 24857 20924 24869 20927
rect 24688 20896 24869 20924
rect 24581 20887 24639 20893
rect 24857 20893 24869 20896
rect 24903 20893 24915 20927
rect 24857 20887 24915 20893
rect 25041 20927 25099 20933
rect 25041 20893 25053 20927
rect 25087 20893 25099 20927
rect 25314 20924 25320 20936
rect 25275 20896 25320 20924
rect 25041 20887 25099 20893
rect 14691 20828 15700 20856
rect 14691 20825 14703 20828
rect 14645 20819 14703 20825
rect 15746 20816 15752 20868
rect 15804 20856 15810 20868
rect 15930 20856 15936 20868
rect 15804 20828 15936 20856
rect 15804 20816 15810 20828
rect 15930 20816 15936 20828
rect 15988 20816 15994 20868
rect 17218 20856 17224 20868
rect 17179 20828 17224 20856
rect 17218 20816 17224 20828
rect 17276 20816 17282 20868
rect 17497 20859 17555 20865
rect 17497 20825 17509 20859
rect 17543 20856 17555 20859
rect 17862 20856 17868 20868
rect 17543 20828 17868 20856
rect 17543 20825 17555 20828
rect 17497 20819 17555 20825
rect 17862 20816 17868 20828
rect 17920 20816 17926 20868
rect 17954 20816 17960 20868
rect 18012 20856 18018 20868
rect 18325 20859 18383 20865
rect 18012 20828 18057 20856
rect 18012 20816 18018 20828
rect 18325 20825 18337 20859
rect 18371 20856 18383 20859
rect 25056 20856 25084 20887
rect 25314 20884 25320 20896
rect 25372 20884 25378 20936
rect 25406 20884 25412 20936
rect 25464 20924 25470 20936
rect 25510 20927 25568 20933
rect 25510 20924 25522 20927
rect 25464 20896 25522 20924
rect 25464 20884 25470 20896
rect 25510 20893 25522 20896
rect 25556 20893 25568 20927
rect 26050 20924 26056 20936
rect 25510 20887 25568 20893
rect 25608 20896 26056 20924
rect 25608 20856 25636 20896
rect 26050 20884 26056 20896
rect 26108 20884 26114 20936
rect 27246 20924 27252 20936
rect 27207 20896 27252 20924
rect 27246 20884 27252 20896
rect 27304 20884 27310 20936
rect 27356 20933 27384 20964
rect 29748 20964 30788 20992
rect 27341 20927 27399 20933
rect 27341 20893 27353 20927
rect 27387 20893 27399 20927
rect 27522 20924 27528 20936
rect 27483 20896 27528 20924
rect 27341 20887 27399 20893
rect 27522 20884 27528 20896
rect 27580 20884 27586 20936
rect 27614 20884 27620 20936
rect 27672 20924 27678 20936
rect 27672 20896 27717 20924
rect 27672 20884 27678 20896
rect 27890 20884 27896 20936
rect 27948 20924 27954 20936
rect 29748 20933 29776 20964
rect 29733 20927 29791 20933
rect 29733 20924 29745 20927
rect 27948 20896 29745 20924
rect 27948 20884 27954 20896
rect 29733 20893 29745 20896
rect 29779 20893 29791 20927
rect 29914 20924 29920 20936
rect 29875 20896 29920 20924
rect 29733 20887 29791 20893
rect 29914 20884 29920 20896
rect 29972 20884 29978 20936
rect 26142 20856 26148 20868
rect 18371 20828 19334 20856
rect 25056 20828 25636 20856
rect 26103 20828 26148 20856
rect 18371 20825 18383 20828
rect 18325 20819 18383 20825
rect 6546 20748 6552 20800
rect 6604 20788 6610 20800
rect 6641 20791 6699 20797
rect 6641 20788 6653 20791
rect 6604 20760 6653 20788
rect 6604 20748 6610 20760
rect 6641 20757 6653 20760
rect 6687 20757 6699 20791
rect 6641 20751 6699 20757
rect 7009 20791 7067 20797
rect 7009 20757 7021 20791
rect 7055 20788 7067 20791
rect 7098 20788 7104 20800
rect 7055 20760 7104 20788
rect 7055 20757 7067 20760
rect 7009 20751 7067 20757
rect 7098 20748 7104 20760
rect 7156 20748 7162 20800
rect 14274 20788 14280 20800
rect 14235 20760 14280 20788
rect 14274 20748 14280 20760
rect 14332 20748 14338 20800
rect 14734 20748 14740 20800
rect 14792 20788 14798 20800
rect 14792 20760 14837 20788
rect 14792 20748 14798 20760
rect 15194 20748 15200 20800
rect 15252 20788 15258 20800
rect 15654 20788 15660 20800
rect 15252 20760 15660 20788
rect 15252 20748 15258 20760
rect 15654 20748 15660 20760
rect 15712 20748 15718 20800
rect 19306 20788 19334 20828
rect 26142 20816 26148 20828
rect 26200 20816 26206 20868
rect 30650 20856 30656 20868
rect 26896 20828 30656 20856
rect 20070 20788 20076 20800
rect 19306 20760 20076 20788
rect 20070 20748 20076 20760
rect 20128 20788 20134 20800
rect 20990 20788 20996 20800
rect 20128 20760 20996 20788
rect 20128 20748 20134 20760
rect 20990 20748 20996 20760
rect 21048 20788 21054 20800
rect 24762 20788 24768 20800
rect 21048 20760 24768 20788
rect 21048 20748 21054 20760
rect 24762 20748 24768 20760
rect 24820 20748 24826 20800
rect 25222 20748 25228 20800
rect 25280 20788 25286 20800
rect 26896 20788 26924 20828
rect 30650 20816 30656 20828
rect 30708 20816 30714 20868
rect 30760 20856 30788 20964
rect 30834 20952 30840 21004
rect 30892 20992 30898 21004
rect 31665 20995 31723 21001
rect 31665 20992 31677 20995
rect 30892 20964 31677 20992
rect 30892 20952 30898 20964
rect 31665 20961 31677 20964
rect 31711 20992 31723 20995
rect 31754 20992 31760 21004
rect 31711 20964 31760 20992
rect 31711 20961 31723 20964
rect 31665 20955 31723 20961
rect 31754 20952 31760 20964
rect 31812 20952 31818 21004
rect 34606 20992 34612 21004
rect 32508 20964 34612 20992
rect 31294 20924 31300 20936
rect 31255 20896 31300 20924
rect 31294 20884 31300 20896
rect 31352 20884 31358 20936
rect 31444 20927 31502 20933
rect 31444 20893 31456 20927
rect 31490 20924 31502 20927
rect 31570 20924 31576 20936
rect 31490 20896 31576 20924
rect 31490 20893 31502 20896
rect 31444 20887 31502 20893
rect 31570 20884 31576 20896
rect 31628 20884 31634 20936
rect 32508 20856 32536 20964
rect 34606 20952 34612 20964
rect 34664 20952 34670 21004
rect 32861 20927 32919 20933
rect 32861 20893 32873 20927
rect 32907 20924 32919 20927
rect 32950 20924 32956 20936
rect 32907 20896 32956 20924
rect 32907 20893 32919 20896
rect 32861 20887 32919 20893
rect 32950 20884 32956 20896
rect 33008 20884 33014 20936
rect 36725 20927 36783 20933
rect 36725 20893 36737 20927
rect 36771 20924 36783 20927
rect 36814 20924 36820 20936
rect 36771 20896 36820 20924
rect 36771 20893 36783 20896
rect 36725 20887 36783 20893
rect 36814 20884 36820 20896
rect 36872 20884 36878 20936
rect 30760 20828 32536 20856
rect 32585 20859 32643 20865
rect 32585 20825 32597 20859
rect 32631 20856 32643 20859
rect 33134 20856 33140 20868
rect 32631 20828 33140 20856
rect 32631 20825 32643 20828
rect 32585 20819 32643 20825
rect 33134 20816 33140 20828
rect 33192 20816 33198 20868
rect 36992 20859 37050 20865
rect 36992 20825 37004 20859
rect 37038 20856 37050 20859
rect 37458 20856 37464 20868
rect 37038 20828 37464 20856
rect 37038 20825 37050 20828
rect 36992 20819 37050 20825
rect 37458 20816 37464 20828
rect 37516 20816 37522 20868
rect 27062 20788 27068 20800
rect 25280 20760 26924 20788
rect 27023 20760 27068 20788
rect 25280 20748 25286 20760
rect 27062 20748 27068 20760
rect 27120 20748 27126 20800
rect 29822 20788 29828 20800
rect 29783 20760 29828 20788
rect 29822 20748 29828 20760
rect 29880 20748 29886 20800
rect 32766 20788 32772 20800
rect 32727 20760 32772 20788
rect 32766 20748 32772 20760
rect 32824 20788 32830 20800
rect 35894 20788 35900 20800
rect 32824 20760 35900 20788
rect 32824 20748 32830 20760
rect 35894 20748 35900 20760
rect 35952 20748 35958 20800
rect 37642 20748 37648 20800
rect 37700 20788 37706 20800
rect 38105 20791 38163 20797
rect 38105 20788 38117 20791
rect 37700 20760 38117 20788
rect 37700 20748 37706 20760
rect 38105 20757 38117 20760
rect 38151 20757 38163 20791
rect 38105 20751 38163 20757
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 4341 20587 4399 20593
rect 4341 20553 4353 20587
rect 4387 20584 4399 20587
rect 4982 20584 4988 20596
rect 4387 20556 4988 20584
rect 4387 20553 4399 20556
rect 4341 20547 4399 20553
rect 4982 20544 4988 20556
rect 5040 20544 5046 20596
rect 9950 20584 9956 20596
rect 9911 20556 9956 20584
rect 9950 20544 9956 20556
rect 10008 20544 10014 20596
rect 13541 20587 13599 20593
rect 13541 20553 13553 20587
rect 13587 20584 13599 20587
rect 13906 20584 13912 20596
rect 13587 20556 13912 20584
rect 13587 20553 13599 20556
rect 13541 20547 13599 20553
rect 13906 20544 13912 20556
rect 13964 20544 13970 20596
rect 14093 20587 14151 20593
rect 14093 20553 14105 20587
rect 14139 20584 14151 20587
rect 14734 20584 14740 20596
rect 14139 20556 14740 20584
rect 14139 20553 14151 20556
rect 14093 20547 14151 20553
rect 14734 20544 14740 20556
rect 14792 20544 14798 20596
rect 18141 20587 18199 20593
rect 15028 20556 18092 20584
rect 9214 20476 9220 20528
rect 9272 20516 9278 20528
rect 9585 20519 9643 20525
rect 9585 20516 9597 20519
rect 9272 20488 9597 20516
rect 9272 20476 9278 20488
rect 9585 20485 9597 20488
rect 9631 20485 9643 20519
rect 9585 20479 9643 20485
rect 9677 20519 9735 20525
rect 9677 20485 9689 20519
rect 9723 20516 9735 20519
rect 10962 20516 10968 20528
rect 9723 20488 10968 20516
rect 9723 20485 9735 20488
rect 9677 20479 9735 20485
rect 10962 20476 10968 20488
rect 11020 20476 11026 20528
rect 12428 20519 12486 20525
rect 12428 20485 12440 20519
rect 12474 20516 12486 20519
rect 14274 20516 14280 20528
rect 12474 20488 14280 20516
rect 12474 20485 12486 20488
rect 12428 20479 12486 20485
rect 14274 20476 14280 20488
rect 14332 20476 14338 20528
rect 4249 20451 4307 20457
rect 4249 20417 4261 20451
rect 4295 20448 4307 20451
rect 5350 20448 5356 20460
rect 4295 20420 5356 20448
rect 4295 20417 4307 20420
rect 4249 20411 4307 20417
rect 5350 20408 5356 20420
rect 5408 20408 5414 20460
rect 6816 20451 6874 20457
rect 6816 20417 6828 20451
rect 6862 20448 6874 20451
rect 7098 20448 7104 20460
rect 6862 20420 7104 20448
rect 6862 20417 6874 20420
rect 6816 20411 6874 20417
rect 7098 20408 7104 20420
rect 7156 20408 7162 20460
rect 9398 20448 9404 20460
rect 9359 20420 9404 20448
rect 9398 20408 9404 20420
rect 9456 20408 9462 20460
rect 9766 20448 9772 20460
rect 9679 20420 9772 20448
rect 9766 20408 9772 20420
rect 9824 20408 9830 20460
rect 14458 20408 14464 20460
rect 14516 20448 14522 20460
rect 14516 20420 14561 20448
rect 14516 20408 14522 20420
rect 4525 20383 4583 20389
rect 4525 20349 4537 20383
rect 4571 20380 4583 20383
rect 4614 20380 4620 20392
rect 4571 20352 4620 20380
rect 4571 20349 4583 20352
rect 4525 20343 4583 20349
rect 4614 20340 4620 20352
rect 4672 20340 4678 20392
rect 6549 20383 6607 20389
rect 6549 20349 6561 20383
rect 6595 20349 6607 20383
rect 6549 20343 6607 20349
rect 3970 20272 3976 20324
rect 4028 20312 4034 20324
rect 6564 20312 6592 20343
rect 4028 20284 6592 20312
rect 9784 20312 9812 20408
rect 11698 20340 11704 20392
rect 11756 20380 11762 20392
rect 12158 20380 12164 20392
rect 11756 20352 12164 20380
rect 11756 20340 11762 20352
rect 12158 20340 12164 20352
rect 12216 20340 12222 20392
rect 14550 20380 14556 20392
rect 14511 20352 14556 20380
rect 14550 20340 14556 20352
rect 14608 20340 14614 20392
rect 14734 20340 14740 20392
rect 14792 20380 14798 20392
rect 15028 20380 15056 20556
rect 15286 20516 15292 20528
rect 15247 20488 15292 20516
rect 15286 20476 15292 20488
rect 15344 20476 15350 20528
rect 15378 20476 15384 20528
rect 15436 20476 15442 20528
rect 15746 20476 15752 20528
rect 15804 20516 15810 20528
rect 17586 20516 17592 20528
rect 15804 20488 17592 20516
rect 15804 20476 15810 20488
rect 17586 20476 17592 20488
rect 17644 20516 17650 20528
rect 18064 20516 18092 20556
rect 18141 20553 18153 20587
rect 18187 20584 18199 20587
rect 22646 20584 22652 20596
rect 18187 20556 22652 20584
rect 18187 20553 18199 20556
rect 18141 20547 18199 20553
rect 22646 20544 22652 20556
rect 22704 20544 22710 20596
rect 22922 20544 22928 20596
rect 22980 20584 22986 20596
rect 23382 20584 23388 20596
rect 22980 20556 23388 20584
rect 22980 20544 22986 20556
rect 23382 20544 23388 20556
rect 23440 20544 23446 20596
rect 24857 20587 24915 20593
rect 24857 20553 24869 20587
rect 24903 20584 24915 20587
rect 25406 20584 25412 20596
rect 24903 20556 25412 20584
rect 24903 20553 24915 20556
rect 24857 20547 24915 20553
rect 25406 20544 25412 20556
rect 25464 20544 25470 20596
rect 25866 20544 25872 20596
rect 25924 20544 25930 20596
rect 27614 20544 27620 20596
rect 27672 20584 27678 20596
rect 27801 20587 27859 20593
rect 27801 20584 27813 20587
rect 27672 20556 27813 20584
rect 27672 20544 27678 20556
rect 27801 20553 27813 20556
rect 27847 20553 27859 20587
rect 27801 20547 27859 20553
rect 28074 20544 28080 20596
rect 28132 20584 28138 20596
rect 32766 20584 32772 20596
rect 28132 20556 32772 20584
rect 28132 20544 28138 20556
rect 32766 20544 32772 20556
rect 32824 20544 32830 20596
rect 33134 20584 33140 20596
rect 33095 20556 33140 20584
rect 33134 20544 33140 20556
rect 33192 20544 33198 20596
rect 33962 20584 33968 20596
rect 33923 20556 33968 20584
rect 33962 20544 33968 20556
rect 34020 20544 34026 20596
rect 37458 20584 37464 20596
rect 37419 20556 37464 20584
rect 37458 20544 37464 20556
rect 37516 20544 37522 20596
rect 20438 20516 20444 20528
rect 17644 20488 18000 20516
rect 18064 20488 20444 20516
rect 17644 20476 17650 20488
rect 15396 20448 15424 20476
rect 15473 20451 15531 20457
rect 15473 20448 15485 20451
rect 15396 20420 15485 20448
rect 15473 20417 15485 20420
rect 15519 20417 15531 20451
rect 15473 20411 15531 20417
rect 15565 20451 15623 20457
rect 15565 20417 15577 20451
rect 15611 20417 15623 20451
rect 15565 20411 15623 20417
rect 15841 20451 15899 20457
rect 15841 20417 15853 20451
rect 15887 20448 15899 20451
rect 16574 20448 16580 20460
rect 15887 20420 16580 20448
rect 15887 20417 15899 20420
rect 15841 20411 15899 20417
rect 14792 20352 15056 20380
rect 14792 20340 14798 20352
rect 15378 20340 15384 20392
rect 15436 20380 15442 20392
rect 15580 20380 15608 20411
rect 16574 20408 16580 20420
rect 16632 20408 16638 20460
rect 17972 20457 18000 20488
rect 20438 20476 20444 20488
rect 20496 20476 20502 20528
rect 25884 20516 25912 20544
rect 22020 20488 25912 20516
rect 17957 20451 18015 20457
rect 17957 20417 17969 20451
rect 18003 20417 18015 20451
rect 17957 20411 18015 20417
rect 18230 20408 18236 20460
rect 18288 20448 18294 20460
rect 22020 20457 22048 20488
rect 26694 20476 26700 20528
rect 26752 20516 26758 20528
rect 27338 20516 27344 20528
rect 26752 20488 27344 20516
rect 26752 20476 26758 20488
rect 27338 20476 27344 20488
rect 27396 20516 27402 20528
rect 27522 20516 27528 20528
rect 27396 20488 27528 20516
rect 27396 20476 27402 20488
rect 27522 20476 27528 20488
rect 27580 20516 27586 20528
rect 28445 20519 28503 20525
rect 28445 20516 28457 20519
rect 27580 20488 28457 20516
rect 27580 20476 27586 20488
rect 28445 20485 28457 20488
rect 28491 20485 28503 20519
rect 29270 20516 29276 20528
rect 29231 20488 29276 20516
rect 28445 20479 28503 20485
rect 29270 20476 29276 20488
rect 29328 20476 29334 20528
rect 32214 20516 32220 20528
rect 29472 20488 32220 20516
rect 19429 20451 19487 20457
rect 19429 20448 19441 20451
rect 18288 20420 19441 20448
rect 18288 20408 18294 20420
rect 19429 20417 19441 20420
rect 19475 20417 19487 20451
rect 19685 20451 19743 20457
rect 19685 20448 19697 20451
rect 19429 20411 19487 20417
rect 19536 20420 19697 20448
rect 15436 20352 15608 20380
rect 15436 20340 15442 20352
rect 15654 20340 15660 20392
rect 15712 20380 15718 20392
rect 15749 20383 15807 20389
rect 15749 20380 15761 20383
rect 15712 20352 15761 20380
rect 15712 20340 15718 20352
rect 15749 20349 15761 20352
rect 15795 20349 15807 20383
rect 15749 20343 15807 20349
rect 18417 20383 18475 20389
rect 18417 20349 18429 20383
rect 18463 20349 18475 20383
rect 18417 20343 18475 20349
rect 11882 20312 11888 20324
rect 9784 20284 11888 20312
rect 4028 20272 4034 20284
rect 11882 20272 11888 20284
rect 11940 20272 11946 20324
rect 16482 20312 16488 20324
rect 13464 20284 16488 20312
rect 3878 20244 3884 20256
rect 3839 20216 3884 20244
rect 3878 20204 3884 20216
rect 3936 20204 3942 20256
rect 6822 20204 6828 20256
rect 6880 20244 6886 20256
rect 7929 20247 7987 20253
rect 7929 20244 7941 20247
rect 6880 20216 7941 20244
rect 6880 20204 6886 20216
rect 7929 20213 7941 20216
rect 7975 20244 7987 20247
rect 13464 20244 13492 20284
rect 16482 20272 16488 20284
rect 16540 20272 16546 20324
rect 18046 20272 18052 20324
rect 18104 20312 18110 20324
rect 18432 20312 18460 20343
rect 18506 20340 18512 20392
rect 18564 20380 18570 20392
rect 18564 20352 18609 20380
rect 18564 20340 18570 20352
rect 19334 20340 19340 20392
rect 19392 20380 19398 20392
rect 19536 20380 19564 20420
rect 19685 20417 19697 20420
rect 19731 20417 19743 20451
rect 19685 20411 19743 20417
rect 22005 20451 22063 20457
rect 22005 20417 22017 20451
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 22094 20408 22100 20460
rect 22152 20448 22158 20460
rect 22272 20451 22330 20457
rect 22272 20448 22284 20451
rect 22152 20420 22284 20448
rect 22152 20408 22158 20420
rect 22272 20417 22284 20420
rect 22318 20417 22330 20451
rect 24026 20448 24032 20460
rect 23987 20420 24032 20448
rect 22272 20411 22330 20417
rect 24026 20408 24032 20420
rect 24084 20408 24090 20460
rect 25038 20448 25044 20460
rect 24999 20420 25044 20448
rect 25038 20408 25044 20420
rect 25096 20408 25102 20460
rect 25130 20408 25136 20460
rect 25188 20448 25194 20460
rect 25225 20451 25283 20457
rect 25225 20448 25237 20451
rect 25188 20420 25237 20448
rect 25188 20408 25194 20420
rect 25225 20417 25237 20420
rect 25271 20417 25283 20451
rect 25225 20411 25283 20417
rect 25317 20451 25375 20457
rect 25317 20417 25329 20451
rect 25363 20417 25375 20451
rect 25317 20411 25375 20417
rect 19392 20352 19564 20380
rect 19392 20340 19398 20352
rect 20898 20340 20904 20392
rect 20956 20380 20962 20392
rect 22112 20380 22140 20408
rect 20956 20352 22140 20380
rect 20956 20340 20962 20352
rect 23842 20340 23848 20392
rect 23900 20380 23906 20392
rect 23937 20383 23995 20389
rect 23937 20380 23949 20383
rect 23900 20352 23949 20380
rect 23900 20340 23906 20352
rect 23937 20349 23949 20352
rect 23983 20349 23995 20383
rect 23937 20343 23995 20349
rect 18104 20284 18460 20312
rect 20809 20315 20867 20321
rect 18104 20272 18110 20284
rect 20809 20281 20821 20315
rect 20855 20312 20867 20315
rect 20990 20312 20996 20324
rect 20855 20284 20996 20312
rect 20855 20281 20867 20284
rect 20809 20275 20867 20281
rect 20990 20272 20996 20284
rect 21048 20272 21054 20324
rect 24397 20315 24455 20321
rect 24397 20281 24409 20315
rect 24443 20312 24455 20315
rect 24762 20312 24768 20324
rect 24443 20284 24768 20312
rect 24443 20281 24455 20284
rect 24397 20275 24455 20281
rect 24762 20272 24768 20284
rect 24820 20312 24826 20324
rect 25332 20312 25360 20411
rect 25774 20408 25780 20460
rect 25832 20448 25838 20460
rect 25869 20451 25927 20457
rect 25869 20448 25881 20451
rect 25832 20420 25881 20448
rect 25832 20408 25838 20420
rect 25869 20417 25881 20420
rect 25915 20417 25927 20451
rect 25869 20411 25927 20417
rect 26016 20451 26074 20457
rect 26016 20417 26028 20451
rect 26062 20448 26074 20451
rect 26602 20448 26608 20460
rect 26062 20420 26608 20448
rect 26062 20417 26074 20420
rect 26016 20411 26074 20417
rect 26602 20408 26608 20420
rect 26660 20408 26666 20460
rect 28077 20451 28135 20457
rect 28077 20417 28089 20451
rect 28123 20448 28135 20451
rect 28123 20420 28488 20448
rect 28123 20417 28135 20420
rect 28077 20411 28135 20417
rect 28460 20392 28488 20420
rect 28810 20408 28816 20460
rect 28868 20448 28874 20460
rect 29362 20448 29368 20460
rect 28868 20420 29368 20448
rect 28868 20408 28874 20420
rect 29362 20408 29368 20420
rect 29420 20448 29426 20460
rect 29472 20457 29500 20488
rect 32214 20476 32220 20488
rect 32272 20476 32278 20528
rect 32861 20519 32919 20525
rect 32861 20485 32873 20519
rect 32907 20516 32919 20519
rect 33226 20516 33232 20528
rect 32907 20488 33232 20516
rect 32907 20485 32919 20488
rect 32861 20479 32919 20485
rect 33226 20476 33232 20488
rect 33284 20476 33290 20528
rect 33594 20516 33600 20528
rect 33555 20488 33600 20516
rect 33594 20476 33600 20488
rect 33652 20476 33658 20528
rect 34164 20488 35664 20516
rect 29457 20451 29515 20457
rect 29457 20448 29469 20451
rect 29420 20420 29469 20448
rect 29420 20408 29426 20420
rect 29457 20417 29469 20420
rect 29503 20417 29515 20451
rect 29638 20448 29644 20460
rect 29599 20420 29644 20448
rect 29457 20411 29515 20417
rect 29638 20408 29644 20420
rect 29696 20408 29702 20460
rect 29733 20451 29791 20457
rect 29733 20417 29745 20451
rect 29779 20448 29791 20451
rect 30098 20448 30104 20460
rect 29779 20420 30104 20448
rect 29779 20417 29791 20420
rect 29733 20411 29791 20417
rect 30098 20408 30104 20420
rect 30156 20408 30162 20460
rect 30746 20451 30804 20457
rect 30746 20448 30758 20451
rect 30208 20420 30758 20448
rect 26237 20383 26295 20389
rect 26237 20349 26249 20383
rect 26283 20380 26295 20383
rect 26418 20380 26424 20392
rect 26283 20352 26424 20380
rect 26283 20349 26295 20352
rect 26237 20343 26295 20349
rect 26418 20340 26424 20352
rect 26476 20380 26482 20392
rect 27798 20380 27804 20392
rect 26476 20352 27804 20380
rect 26476 20340 26482 20352
rect 27798 20340 27804 20352
rect 27856 20340 27862 20392
rect 27982 20380 27988 20392
rect 27943 20352 27988 20380
rect 27982 20340 27988 20352
rect 28040 20340 28046 20392
rect 28258 20340 28264 20392
rect 28316 20380 28322 20392
rect 28353 20383 28411 20389
rect 28353 20380 28365 20383
rect 28316 20352 28365 20380
rect 28316 20340 28322 20352
rect 28353 20349 28365 20352
rect 28399 20349 28411 20383
rect 28353 20343 28411 20349
rect 28442 20340 28448 20392
rect 28500 20340 28506 20392
rect 29178 20340 29184 20392
rect 29236 20380 29242 20392
rect 29914 20380 29920 20392
rect 29236 20352 29920 20380
rect 29236 20340 29242 20352
rect 29914 20340 29920 20352
rect 29972 20340 29978 20392
rect 24820 20284 25360 20312
rect 24820 20272 24826 20284
rect 25406 20272 25412 20324
rect 25464 20312 25470 20324
rect 30208 20312 30236 20420
rect 30746 20417 30758 20420
rect 30792 20417 30804 20451
rect 32490 20448 32496 20460
rect 32451 20420 32496 20448
rect 30746 20411 30804 20417
rect 32490 20408 32496 20420
rect 32548 20408 32554 20460
rect 32674 20457 32680 20460
rect 32641 20451 32680 20457
rect 32641 20417 32653 20451
rect 32641 20411 32680 20417
rect 32674 20408 32680 20411
rect 32732 20408 32738 20460
rect 32766 20408 32772 20460
rect 32824 20448 32830 20460
rect 33042 20457 33048 20460
rect 32999 20451 33048 20457
rect 32824 20420 32869 20448
rect 32824 20408 32830 20420
rect 32999 20417 33011 20451
rect 33045 20417 33048 20451
rect 32999 20411 33048 20417
rect 33042 20408 33048 20411
rect 33100 20408 33106 20460
rect 33134 20408 33140 20460
rect 33192 20448 33198 20460
rect 33781 20451 33839 20457
rect 33781 20448 33793 20451
rect 33192 20420 33793 20448
rect 33192 20408 33198 20420
rect 33781 20417 33793 20420
rect 33827 20417 33839 20451
rect 33781 20411 33839 20417
rect 30650 20340 30656 20392
rect 30708 20380 30714 20392
rect 31113 20383 31171 20389
rect 31113 20380 31125 20383
rect 30708 20352 31125 20380
rect 30708 20340 30714 20352
rect 31113 20349 31125 20352
rect 31159 20349 31171 20383
rect 31113 20343 31171 20349
rect 31205 20383 31263 20389
rect 31205 20349 31217 20383
rect 31251 20380 31263 20383
rect 31478 20380 31484 20392
rect 31251 20352 31484 20380
rect 31251 20349 31263 20352
rect 31205 20343 31263 20349
rect 25464 20284 30236 20312
rect 25464 20272 25470 20284
rect 7975 20216 13492 20244
rect 7975 20213 7987 20216
rect 7929 20207 7987 20213
rect 13998 20204 14004 20256
rect 14056 20244 14062 20256
rect 14458 20244 14464 20256
rect 14056 20216 14464 20244
rect 14056 20204 14062 20216
rect 14458 20204 14464 20216
rect 14516 20244 14522 20256
rect 20530 20244 20536 20256
rect 14516 20216 20536 20244
rect 14516 20204 14522 20216
rect 20530 20204 20536 20216
rect 20588 20204 20594 20256
rect 22278 20204 22284 20256
rect 22336 20244 22342 20256
rect 25222 20244 25228 20256
rect 22336 20216 25228 20244
rect 22336 20204 22342 20216
rect 25222 20204 25228 20216
rect 25280 20204 25286 20256
rect 26145 20247 26203 20253
rect 26145 20213 26157 20247
rect 26191 20244 26203 20247
rect 26326 20244 26332 20256
rect 26191 20216 26332 20244
rect 26191 20213 26203 20216
rect 26145 20207 26203 20213
rect 26326 20204 26332 20216
rect 26384 20204 26390 20256
rect 26513 20247 26571 20253
rect 26513 20213 26525 20247
rect 26559 20244 26571 20247
rect 26878 20244 26884 20256
rect 26559 20216 26884 20244
rect 26559 20213 26571 20216
rect 26513 20207 26571 20213
rect 26878 20204 26884 20216
rect 26936 20204 26942 20256
rect 28258 20204 28264 20256
rect 28316 20244 28322 20256
rect 29454 20244 29460 20256
rect 28316 20216 29460 20244
rect 28316 20204 28322 20216
rect 29454 20204 29460 20216
rect 29512 20204 29518 20256
rect 30650 20244 30656 20256
rect 30611 20216 30656 20244
rect 30650 20204 30656 20216
rect 30708 20204 30714 20256
rect 31128 20244 31156 20343
rect 31478 20340 31484 20352
rect 31536 20340 31542 20392
rect 31294 20272 31300 20324
rect 31352 20312 31358 20324
rect 31938 20312 31944 20324
rect 31352 20284 31944 20312
rect 31352 20272 31358 20284
rect 31938 20272 31944 20284
rect 31996 20272 32002 20324
rect 32766 20272 32772 20324
rect 32824 20312 32830 20324
rect 34164 20312 34192 20488
rect 35526 20448 35532 20460
rect 35487 20420 35532 20448
rect 35526 20408 35532 20420
rect 35584 20408 35590 20460
rect 35636 20457 35664 20488
rect 35621 20451 35679 20457
rect 35621 20417 35633 20451
rect 35667 20417 35679 20451
rect 35894 20448 35900 20460
rect 35855 20420 35900 20448
rect 35621 20411 35679 20417
rect 35894 20408 35900 20420
rect 35952 20408 35958 20460
rect 37642 20408 37648 20460
rect 37700 20448 37706 20460
rect 37829 20451 37887 20457
rect 37829 20448 37841 20451
rect 37700 20420 37841 20448
rect 37700 20408 37706 20420
rect 37829 20417 37841 20420
rect 37875 20417 37887 20451
rect 37829 20411 37887 20417
rect 35345 20383 35403 20389
rect 35345 20349 35357 20383
rect 35391 20380 35403 20383
rect 37921 20383 37979 20389
rect 37921 20380 37933 20383
rect 35391 20352 37933 20380
rect 35391 20349 35403 20352
rect 35345 20343 35403 20349
rect 37844 20324 37872 20352
rect 37921 20349 37933 20352
rect 37967 20349 37979 20383
rect 37921 20343 37979 20349
rect 38010 20340 38016 20392
rect 38068 20380 38074 20392
rect 38068 20352 38113 20380
rect 38068 20340 38074 20352
rect 32824 20284 34192 20312
rect 35805 20315 35863 20321
rect 32824 20272 32830 20284
rect 35805 20281 35817 20315
rect 35851 20312 35863 20315
rect 35986 20312 35992 20324
rect 35851 20284 35992 20312
rect 35851 20281 35863 20284
rect 35805 20275 35863 20281
rect 35986 20272 35992 20284
rect 36044 20312 36050 20324
rect 36538 20312 36544 20324
rect 36044 20284 36544 20312
rect 36044 20272 36050 20284
rect 36538 20272 36544 20284
rect 36596 20272 36602 20324
rect 37826 20272 37832 20324
rect 37884 20272 37890 20324
rect 34514 20244 34520 20256
rect 31128 20216 34520 20244
rect 34514 20204 34520 20216
rect 34572 20204 34578 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 7098 20040 7104 20052
rect 7059 20012 7104 20040
rect 7098 20000 7104 20012
rect 7156 20000 7162 20052
rect 12621 20043 12679 20049
rect 12621 20040 12633 20043
rect 10520 20012 12633 20040
rect 5350 19972 5356 19984
rect 5263 19944 5356 19972
rect 5350 19932 5356 19944
rect 5408 19972 5414 19984
rect 10410 19972 10416 19984
rect 5408 19944 10416 19972
rect 5408 19932 5414 19944
rect 10410 19932 10416 19944
rect 10468 19932 10474 19984
rect 3970 19904 3976 19916
rect 3931 19876 3976 19904
rect 3970 19864 3976 19876
rect 4028 19864 4034 19916
rect 9674 19904 9680 19916
rect 8312 19876 9680 19904
rect 3878 19796 3884 19848
rect 3936 19836 3942 19848
rect 4229 19839 4287 19845
rect 4229 19836 4241 19839
rect 3936 19808 4241 19836
rect 3936 19796 3942 19808
rect 4229 19805 4241 19808
rect 4275 19805 4287 19839
rect 6546 19836 6552 19848
rect 6507 19808 6552 19836
rect 4229 19799 4287 19805
rect 6546 19796 6552 19808
rect 6604 19796 6610 19848
rect 6822 19836 6828 19848
rect 6783 19808 6828 19836
rect 6822 19796 6828 19808
rect 6880 19796 6886 19848
rect 6914 19796 6920 19848
rect 6972 19836 6978 19848
rect 8202 19836 8208 19848
rect 6972 19808 8208 19836
rect 6972 19796 6978 19808
rect 8202 19796 8208 19808
rect 8260 19796 8266 19848
rect 8312 19845 8340 19876
rect 9674 19864 9680 19876
rect 9732 19864 9738 19916
rect 8297 19839 8355 19845
rect 8297 19805 8309 19839
rect 8343 19805 8355 19839
rect 8297 19799 8355 19805
rect 8481 19839 8539 19845
rect 8481 19805 8493 19839
rect 8527 19805 8539 19839
rect 10226 19836 10232 19848
rect 10187 19808 10232 19836
rect 8481 19799 8539 19805
rect 6730 19768 6736 19780
rect 6691 19740 6736 19768
rect 6730 19728 6736 19740
rect 6788 19728 6794 19780
rect 8220 19768 8248 19796
rect 8496 19768 8524 19799
rect 10226 19796 10232 19808
rect 10284 19796 10290 19848
rect 10520 19845 10548 20012
rect 12621 20009 12633 20012
rect 12667 20040 12679 20043
rect 13814 20040 13820 20052
rect 12667 20012 13820 20040
rect 12667 20009 12679 20012
rect 12621 20003 12679 20009
rect 13814 20000 13820 20012
rect 13872 20000 13878 20052
rect 14550 20000 14556 20052
rect 14608 20040 14614 20052
rect 14921 20043 14979 20049
rect 14921 20040 14933 20043
rect 14608 20012 14933 20040
rect 14608 20000 14614 20012
rect 14921 20009 14933 20012
rect 14967 20009 14979 20043
rect 14921 20003 14979 20009
rect 16482 20000 16488 20052
rect 16540 20040 16546 20052
rect 16577 20043 16635 20049
rect 16577 20040 16589 20043
rect 16540 20012 16589 20040
rect 16540 20000 16546 20012
rect 16577 20009 16589 20012
rect 16623 20009 16635 20043
rect 16577 20003 16635 20009
rect 19886 20000 19892 20052
rect 19944 20040 19950 20052
rect 20254 20040 20260 20052
rect 19944 20012 20260 20040
rect 19944 20000 19950 20012
rect 20254 20000 20260 20012
rect 20312 20000 20318 20052
rect 22278 20040 22284 20052
rect 22020 20012 22284 20040
rect 18506 19932 18512 19984
rect 18564 19972 18570 19984
rect 20530 19972 20536 19984
rect 18564 19944 20392 19972
rect 20491 19944 20536 19972
rect 18564 19932 18570 19944
rect 15565 19907 15623 19913
rect 15565 19873 15577 19907
rect 15611 19904 15623 19907
rect 16574 19904 16580 19916
rect 15611 19876 16580 19904
rect 15611 19873 15623 19876
rect 15565 19867 15623 19873
rect 16574 19864 16580 19876
rect 16632 19864 16638 19916
rect 16666 19864 16672 19916
rect 16724 19904 16730 19916
rect 18524 19904 18552 19932
rect 19426 19904 19432 19916
rect 16724 19876 16769 19904
rect 16868 19876 18552 19904
rect 19387 19876 19432 19904
rect 16724 19864 16730 19876
rect 10505 19839 10563 19845
rect 10505 19805 10517 19839
rect 10551 19805 10563 19839
rect 10505 19799 10563 19805
rect 10594 19796 10600 19848
rect 10652 19836 10658 19848
rect 11241 19839 11299 19845
rect 10652 19808 10697 19836
rect 10652 19796 10658 19808
rect 11241 19805 11253 19839
rect 11287 19836 11299 19839
rect 11287 19808 11744 19836
rect 11287 19805 11299 19808
rect 11241 19799 11299 19805
rect 11716 19780 11744 19808
rect 15930 19796 15936 19848
rect 15988 19836 15994 19848
rect 16868 19845 16896 19876
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 20254 19904 20260 19916
rect 19628 19876 20260 19904
rect 16853 19839 16911 19845
rect 16853 19836 16865 19839
rect 15988 19808 16865 19836
rect 15988 19796 15994 19808
rect 16853 19805 16865 19808
rect 16899 19805 16911 19839
rect 16853 19799 16911 19805
rect 17402 19796 17408 19848
rect 17460 19836 17466 19848
rect 17497 19839 17555 19845
rect 17497 19836 17509 19839
rect 17460 19808 17509 19836
rect 17460 19796 17466 19808
rect 17497 19805 17509 19808
rect 17543 19836 17555 19839
rect 18138 19836 18144 19848
rect 17543 19808 18144 19836
rect 17543 19805 17555 19808
rect 17497 19799 17555 19805
rect 18138 19796 18144 19808
rect 18196 19796 18202 19848
rect 18414 19796 18420 19848
rect 18472 19836 18478 19848
rect 19628 19845 19656 19876
rect 20254 19864 20260 19876
rect 20312 19864 20318 19916
rect 19613 19839 19671 19845
rect 19613 19836 19625 19839
rect 18472 19808 19625 19836
rect 18472 19796 18478 19808
rect 19613 19805 19625 19808
rect 19659 19805 19671 19839
rect 19886 19836 19892 19848
rect 19847 19808 19892 19836
rect 19613 19799 19671 19805
rect 19886 19796 19892 19808
rect 19944 19796 19950 19848
rect 20073 19839 20131 19845
rect 20073 19805 20085 19839
rect 20119 19836 20131 19839
rect 20364 19836 20392 19944
rect 20530 19932 20536 19944
rect 20588 19932 20594 19984
rect 20806 19864 20812 19916
rect 20864 19904 20870 19916
rect 21085 19907 21143 19913
rect 21085 19904 21097 19907
rect 20864 19876 21097 19904
rect 20864 19864 20870 19876
rect 21085 19873 21097 19876
rect 21131 19873 21143 19907
rect 21085 19867 21143 19873
rect 20898 19836 20904 19848
rect 20119 19808 20392 19836
rect 20859 19808 20904 19836
rect 20119 19805 20131 19808
rect 20073 19799 20131 19805
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 20993 19839 21051 19845
rect 20993 19805 21005 19839
rect 21039 19836 21051 19839
rect 21358 19836 21364 19848
rect 21039 19808 21364 19836
rect 21039 19805 21051 19808
rect 20993 19799 21051 19805
rect 21358 19796 21364 19808
rect 21416 19796 21422 19848
rect 22020 19845 22048 20012
rect 22278 20000 22284 20012
rect 22336 20000 22342 20052
rect 22370 20000 22376 20052
rect 22428 20040 22434 20052
rect 24765 20043 24823 20049
rect 22428 20012 23796 20040
rect 22428 20000 22434 20012
rect 22094 19932 22100 19984
rect 22152 19972 22158 19984
rect 22388 19972 22416 20000
rect 22152 19944 22416 19972
rect 22152 19932 22158 19944
rect 22738 19932 22744 19984
rect 22796 19972 22802 19984
rect 23661 19975 23719 19981
rect 23661 19972 23673 19975
rect 22796 19944 23673 19972
rect 22796 19932 22802 19944
rect 23661 19941 23673 19944
rect 23707 19941 23719 19975
rect 23661 19935 23719 19941
rect 22204 19876 23336 19904
rect 22005 19839 22063 19845
rect 22005 19805 22017 19839
rect 22051 19805 22063 19839
rect 22005 19799 22063 19805
rect 22204 19780 22232 19876
rect 22370 19796 22376 19848
rect 22428 19845 22434 19848
rect 22428 19836 22436 19845
rect 23109 19839 23167 19845
rect 22428 19808 22473 19836
rect 22428 19799 22436 19808
rect 23109 19805 23121 19839
rect 23155 19836 23167 19839
rect 23198 19836 23204 19848
rect 23155 19808 23204 19836
rect 23155 19805 23167 19808
rect 23109 19799 23167 19805
rect 22428 19796 22434 19799
rect 23198 19796 23204 19808
rect 23256 19796 23262 19848
rect 23308 19845 23336 19876
rect 23293 19839 23351 19845
rect 23293 19805 23305 19839
rect 23339 19805 23351 19839
rect 23293 19799 23351 19805
rect 23529 19839 23587 19845
rect 23529 19805 23541 19839
rect 23575 19836 23587 19839
rect 23768 19836 23796 20012
rect 24765 20009 24777 20043
rect 24811 20040 24823 20043
rect 25314 20040 25320 20052
rect 24811 20012 25320 20040
rect 24811 20009 24823 20012
rect 24765 20003 24823 20009
rect 25314 20000 25320 20012
rect 25372 20000 25378 20052
rect 29270 20000 29276 20052
rect 29328 20040 29334 20052
rect 29733 20043 29791 20049
rect 29733 20040 29745 20043
rect 29328 20012 29745 20040
rect 29328 20000 29334 20012
rect 29733 20009 29745 20012
rect 29779 20009 29791 20043
rect 29733 20003 29791 20009
rect 35894 20000 35900 20052
rect 35952 20040 35958 20052
rect 36265 20043 36323 20049
rect 36265 20040 36277 20043
rect 35952 20012 36277 20040
rect 35952 20000 35958 20012
rect 36265 20009 36277 20012
rect 36311 20009 36323 20043
rect 36265 20003 36323 20009
rect 23934 19932 23940 19984
rect 23992 19972 23998 19984
rect 25958 19972 25964 19984
rect 23992 19944 25964 19972
rect 23992 19932 23998 19944
rect 25958 19932 25964 19944
rect 26016 19932 26022 19984
rect 26326 19932 26332 19984
rect 26384 19972 26390 19984
rect 30742 19972 30748 19984
rect 26384 19944 30748 19972
rect 26384 19932 26390 19944
rect 30742 19932 30748 19944
rect 30800 19932 30806 19984
rect 30929 19975 30987 19981
rect 30929 19941 30941 19975
rect 30975 19972 30987 19975
rect 32030 19972 32036 19984
rect 30975 19944 32036 19972
rect 30975 19941 30987 19944
rect 30929 19935 30987 19941
rect 32030 19932 32036 19944
rect 32088 19932 32094 19984
rect 33594 19972 33600 19984
rect 33244 19944 33600 19972
rect 28074 19904 28080 19916
rect 23575 19808 23796 19836
rect 24228 19876 28080 19904
rect 23575 19805 23587 19808
rect 23529 19799 23587 19805
rect 9766 19768 9772 19780
rect 8220 19740 9772 19768
rect 9766 19728 9772 19740
rect 9824 19768 9830 19780
rect 10318 19768 10324 19780
rect 9824 19740 10324 19768
rect 9824 19728 9830 19740
rect 10318 19728 10324 19740
rect 10376 19728 10382 19780
rect 10413 19771 10471 19777
rect 10413 19737 10425 19771
rect 10459 19737 10471 19771
rect 11486 19771 11544 19777
rect 11486 19768 11498 19771
rect 10413 19731 10471 19737
rect 10796 19740 11498 19768
rect 8386 19700 8392 19712
rect 8347 19672 8392 19700
rect 8386 19660 8392 19672
rect 8444 19700 8450 19712
rect 10428 19700 10456 19731
rect 10796 19709 10824 19740
rect 11486 19737 11498 19740
rect 11532 19737 11544 19771
rect 11486 19731 11544 19737
rect 11698 19728 11704 19780
rect 11756 19728 11762 19780
rect 15194 19728 15200 19780
rect 15252 19768 15258 19780
rect 15381 19771 15439 19777
rect 15381 19768 15393 19771
rect 15252 19740 15393 19768
rect 15252 19728 15258 19740
rect 15381 19737 15393 19740
rect 15427 19768 15439 19771
rect 16298 19768 16304 19780
rect 15427 19740 16304 19768
rect 15427 19737 15439 19740
rect 15381 19731 15439 19737
rect 16298 19728 16304 19740
rect 16356 19728 16362 19780
rect 16574 19768 16580 19780
rect 16535 19740 16580 19768
rect 16574 19728 16580 19740
rect 16632 19728 16638 19780
rect 17770 19728 17776 19780
rect 17828 19768 17834 19780
rect 18693 19771 18751 19777
rect 18693 19768 18705 19771
rect 17828 19740 18705 19768
rect 17828 19728 17834 19740
rect 18693 19737 18705 19740
rect 18739 19768 18751 19771
rect 21910 19768 21916 19780
rect 18739 19740 21916 19768
rect 18739 19737 18751 19740
rect 18693 19731 18751 19737
rect 21910 19728 21916 19740
rect 21968 19728 21974 19780
rect 22186 19768 22192 19780
rect 22147 19740 22192 19768
rect 22186 19728 22192 19740
rect 22244 19728 22250 19780
rect 22281 19771 22339 19777
rect 22281 19737 22293 19771
rect 22327 19768 22339 19771
rect 23385 19771 23443 19777
rect 22327 19740 23336 19768
rect 22327 19737 22339 19740
rect 22281 19731 22339 19737
rect 8444 19672 10456 19700
rect 10781 19703 10839 19709
rect 8444 19660 8450 19672
rect 10781 19669 10793 19703
rect 10827 19669 10839 19703
rect 15286 19700 15292 19712
rect 15247 19672 15292 19700
rect 10781 19663 10839 19669
rect 15286 19660 15292 19672
rect 15344 19660 15350 19712
rect 17037 19703 17095 19709
rect 17037 19669 17049 19703
rect 17083 19700 17095 19703
rect 18506 19700 18512 19712
rect 17083 19672 18512 19700
rect 17083 19669 17095 19672
rect 17037 19663 17095 19669
rect 18506 19660 18512 19672
rect 18564 19660 18570 19712
rect 18782 19660 18788 19712
rect 18840 19700 18846 19712
rect 22565 19703 22623 19709
rect 22565 19700 22577 19703
rect 18840 19672 22577 19700
rect 18840 19660 18846 19672
rect 22565 19669 22577 19672
rect 22611 19669 22623 19703
rect 23308 19700 23336 19740
rect 23385 19737 23397 19771
rect 23431 19768 23443 19771
rect 24228 19768 24256 19876
rect 28074 19864 28080 19876
rect 28132 19864 28138 19916
rect 29822 19904 29828 19916
rect 29783 19876 29828 19904
rect 29822 19864 29828 19876
rect 29880 19864 29886 19916
rect 30374 19864 30380 19916
rect 30432 19904 30438 19916
rect 33244 19913 33272 19944
rect 33594 19932 33600 19944
rect 33652 19932 33658 19984
rect 31297 19907 31355 19913
rect 31297 19904 31309 19907
rect 30432 19876 31309 19904
rect 30432 19864 30438 19876
rect 31297 19873 31309 19876
rect 31343 19904 31355 19907
rect 33229 19907 33287 19913
rect 31343 19876 31754 19904
rect 31343 19873 31355 19876
rect 31297 19867 31355 19873
rect 24762 19836 24768 19848
rect 24723 19808 24768 19836
rect 24762 19796 24768 19808
rect 24820 19796 24826 19848
rect 24949 19839 25007 19845
rect 24949 19805 24961 19839
rect 24995 19836 25007 19839
rect 25130 19836 25136 19848
rect 24995 19808 25136 19836
rect 24995 19805 25007 19808
rect 24949 19799 25007 19805
rect 25130 19796 25136 19808
rect 25188 19796 25194 19848
rect 26878 19796 26884 19848
rect 26936 19836 26942 19848
rect 27249 19839 27307 19845
rect 27249 19836 27261 19839
rect 26936 19808 27261 19836
rect 26936 19796 26942 19808
rect 27249 19805 27261 19808
rect 27295 19805 27307 19839
rect 27249 19799 27307 19805
rect 27617 19839 27675 19845
rect 27617 19805 27629 19839
rect 27663 19836 27675 19839
rect 27982 19836 27988 19848
rect 27663 19808 27988 19836
rect 27663 19805 27675 19808
rect 27617 19799 27675 19805
rect 27982 19796 27988 19808
rect 28040 19836 28046 19848
rect 29178 19836 29184 19848
rect 28040 19808 29184 19836
rect 28040 19796 28046 19808
rect 29178 19796 29184 19808
rect 29236 19836 29242 19848
rect 29454 19836 29460 19848
rect 29236 19808 29460 19836
rect 29236 19796 29242 19808
rect 29454 19796 29460 19808
rect 29512 19796 29518 19848
rect 29730 19836 29736 19848
rect 29691 19808 29736 19836
rect 29730 19796 29736 19808
rect 29788 19796 29794 19848
rect 31110 19796 31116 19848
rect 31168 19836 31174 19848
rect 31478 19836 31484 19848
rect 31168 19808 31484 19836
rect 31168 19796 31174 19808
rect 31478 19796 31484 19808
rect 31536 19796 31542 19848
rect 27062 19768 27068 19780
rect 23431 19740 24256 19768
rect 27023 19740 27068 19768
rect 23431 19737 23443 19740
rect 23385 19731 23443 19737
rect 27062 19728 27068 19740
rect 27120 19728 27126 19780
rect 29270 19768 29276 19780
rect 28966 19740 29276 19768
rect 24578 19700 24584 19712
rect 23308 19672 24584 19700
rect 22565 19663 22623 19669
rect 24578 19660 24584 19672
rect 24636 19660 24642 19712
rect 28626 19660 28632 19712
rect 28684 19700 28690 19712
rect 28966 19700 28994 19740
rect 29270 19728 29276 19740
rect 29328 19768 29334 19780
rect 30282 19768 30288 19780
rect 29328 19740 30288 19768
rect 29328 19728 29334 19740
rect 30282 19728 30288 19740
rect 30340 19728 30346 19780
rect 31726 19768 31754 19876
rect 33229 19873 33241 19907
rect 33275 19873 33287 19907
rect 33229 19867 33287 19873
rect 33505 19907 33563 19913
rect 33505 19873 33517 19907
rect 33551 19873 33563 19907
rect 38102 19904 38108 19916
rect 38063 19876 38108 19904
rect 33505 19867 33563 19873
rect 33134 19836 33140 19848
rect 33095 19808 33140 19836
rect 33134 19796 33140 19808
rect 33192 19796 33198 19848
rect 33226 19768 33232 19780
rect 31726 19740 33232 19768
rect 33226 19728 33232 19740
rect 33284 19728 33290 19780
rect 33520 19768 33548 19867
rect 38102 19864 38108 19876
rect 38160 19864 38166 19916
rect 34885 19839 34943 19845
rect 34885 19805 34897 19839
rect 34931 19836 34943 19839
rect 36814 19836 36820 19848
rect 34931 19808 36820 19836
rect 34931 19805 34943 19808
rect 34885 19799 34943 19805
rect 36814 19796 36820 19808
rect 36872 19796 36878 19848
rect 37826 19836 37832 19848
rect 37787 19808 37832 19836
rect 37826 19796 37832 19808
rect 37884 19796 37890 19848
rect 35130 19771 35188 19777
rect 35130 19768 35142 19771
rect 33520 19740 35142 19768
rect 35130 19737 35142 19740
rect 35176 19737 35188 19771
rect 35130 19731 35188 19737
rect 28684 19672 28994 19700
rect 28684 19660 28690 19672
rect 29546 19660 29552 19712
rect 29604 19700 29610 19712
rect 30101 19703 30159 19709
rect 30101 19700 30113 19703
rect 29604 19672 30113 19700
rect 29604 19660 29610 19672
rect 30101 19669 30113 19672
rect 30147 19669 30159 19703
rect 30101 19663 30159 19669
rect 31018 19660 31024 19712
rect 31076 19700 31082 19712
rect 31389 19703 31447 19709
rect 31389 19700 31401 19703
rect 31076 19672 31401 19700
rect 31076 19660 31082 19672
rect 31389 19669 31401 19672
rect 31435 19700 31447 19703
rect 34974 19700 34980 19712
rect 31435 19672 34980 19700
rect 31435 19669 31447 19672
rect 31389 19663 31447 19669
rect 34974 19660 34980 19672
rect 35032 19660 35038 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 9490 19496 9496 19508
rect 8036 19468 9496 19496
rect 5445 19431 5503 19437
rect 5445 19397 5457 19431
rect 5491 19428 5503 19431
rect 5626 19428 5632 19440
rect 5491 19400 5632 19428
rect 5491 19397 5503 19400
rect 5445 19391 5503 19397
rect 5626 19388 5632 19400
rect 5684 19388 5690 19440
rect 4614 19320 4620 19372
rect 4672 19360 4678 19372
rect 4672 19332 5672 19360
rect 4672 19320 4678 19332
rect 5537 19295 5595 19301
rect 5537 19261 5549 19295
rect 5583 19261 5595 19295
rect 5644 19292 5672 19332
rect 6730 19320 6736 19372
rect 6788 19360 6794 19372
rect 8036 19369 8064 19468
rect 9490 19456 9496 19468
rect 9548 19456 9554 19508
rect 15286 19496 15292 19508
rect 15247 19468 15292 19496
rect 15286 19456 15292 19468
rect 15344 19456 15350 19508
rect 16574 19456 16580 19508
rect 16632 19496 16638 19508
rect 17405 19499 17463 19505
rect 17405 19496 17417 19499
rect 16632 19468 17417 19496
rect 16632 19456 16638 19468
rect 17405 19465 17417 19468
rect 17451 19465 17463 19499
rect 19334 19496 19340 19508
rect 19295 19468 19340 19496
rect 17405 19459 17463 19465
rect 19334 19456 19340 19468
rect 19392 19456 19398 19508
rect 19797 19499 19855 19505
rect 19797 19465 19809 19499
rect 19843 19496 19855 19499
rect 20530 19496 20536 19508
rect 19843 19468 20536 19496
rect 19843 19465 19855 19468
rect 19797 19459 19855 19465
rect 20530 19456 20536 19468
rect 20588 19456 20594 19508
rect 26878 19496 26884 19508
rect 20732 19468 22876 19496
rect 8205 19431 8263 19437
rect 8205 19397 8217 19431
rect 8251 19397 8263 19431
rect 8205 19391 8263 19397
rect 8297 19431 8355 19437
rect 8297 19397 8309 19431
rect 8343 19428 8355 19431
rect 9306 19428 9312 19440
rect 8343 19400 9312 19428
rect 8343 19397 8355 19400
rect 8297 19391 8355 19397
rect 8021 19363 8079 19369
rect 6788 19332 7972 19360
rect 6788 19320 6794 19332
rect 5721 19295 5779 19301
rect 5721 19292 5733 19295
rect 5644 19264 5733 19292
rect 5537 19255 5595 19261
rect 5721 19261 5733 19264
rect 5767 19292 5779 19295
rect 7098 19292 7104 19304
rect 5767 19264 7104 19292
rect 5767 19261 5779 19264
rect 5721 19255 5779 19261
rect 5552 19224 5580 19255
rect 7098 19252 7104 19264
rect 7156 19252 7162 19304
rect 7944 19292 7972 19332
rect 8021 19329 8033 19363
rect 8067 19329 8079 19363
rect 8021 19323 8079 19329
rect 8220 19292 8248 19391
rect 9306 19388 9312 19400
rect 9364 19388 9370 19440
rect 12342 19428 12348 19440
rect 11716 19400 12348 19428
rect 8389 19363 8447 19369
rect 8389 19360 8401 19363
rect 7944 19264 8248 19292
rect 8312 19332 8401 19360
rect 7374 19224 7380 19236
rect 5552 19196 7380 19224
rect 7374 19184 7380 19196
rect 7432 19184 7438 19236
rect 5074 19156 5080 19168
rect 5035 19128 5080 19156
rect 5074 19116 5080 19128
rect 5132 19116 5138 19168
rect 8128 19156 8156 19264
rect 8202 19184 8208 19236
rect 8260 19224 8266 19236
rect 8312 19224 8340 19332
rect 8389 19329 8401 19332
rect 8435 19329 8447 19363
rect 8389 19323 8447 19329
rect 9122 19320 9128 19372
rect 9180 19360 9186 19372
rect 9401 19363 9459 19369
rect 9401 19360 9413 19363
rect 9180 19332 9413 19360
rect 9180 19320 9186 19332
rect 9401 19329 9413 19332
rect 9447 19329 9459 19363
rect 9401 19323 9459 19329
rect 9668 19363 9726 19369
rect 9668 19329 9680 19363
rect 9714 19360 9726 19363
rect 9950 19360 9956 19372
rect 9714 19332 9956 19360
rect 9714 19329 9726 19332
rect 9668 19323 9726 19329
rect 9950 19320 9956 19332
rect 10008 19320 10014 19372
rect 10594 19320 10600 19372
rect 10652 19360 10658 19372
rect 11716 19369 11744 19400
rect 12342 19388 12348 19400
rect 12400 19428 12406 19440
rect 16666 19428 16672 19440
rect 12400 19400 16672 19428
rect 12400 19388 12406 19400
rect 16666 19388 16672 19400
rect 16724 19388 16730 19440
rect 19705 19431 19763 19437
rect 19705 19397 19717 19431
rect 19751 19428 19763 19431
rect 20070 19428 20076 19440
rect 19751 19400 20076 19428
rect 19751 19397 19763 19400
rect 19705 19391 19763 19397
rect 20070 19388 20076 19400
rect 20128 19388 20134 19440
rect 20732 19437 20760 19468
rect 20717 19431 20775 19437
rect 20717 19428 20729 19431
rect 20627 19400 20729 19428
rect 11701 19363 11759 19369
rect 10652 19332 11652 19360
rect 10652 19320 10658 19332
rect 11624 19292 11652 19332
rect 11701 19329 11713 19363
rect 11747 19329 11759 19363
rect 11977 19363 12035 19369
rect 11977 19360 11989 19363
rect 11701 19323 11759 19329
rect 11808 19332 11989 19360
rect 11808 19292 11836 19332
rect 11977 19329 11989 19332
rect 12023 19329 12035 19363
rect 15654 19360 15660 19372
rect 15615 19332 15660 19360
rect 11977 19323 12035 19329
rect 15654 19320 15660 19332
rect 15712 19320 15718 19372
rect 15746 19320 15752 19372
rect 15804 19360 15810 19372
rect 17586 19360 17592 19372
rect 15804 19332 15849 19360
rect 17547 19332 17592 19360
rect 15804 19320 15810 19332
rect 17586 19320 17592 19332
rect 17644 19320 17650 19372
rect 17770 19360 17776 19372
rect 17731 19332 17776 19360
rect 17770 19320 17776 19332
rect 17828 19320 17834 19372
rect 18506 19360 18512 19372
rect 18467 19332 18512 19360
rect 18506 19320 18512 19332
rect 18564 19320 18570 19372
rect 18598 19320 18604 19372
rect 18656 19360 18662 19372
rect 18877 19363 18935 19369
rect 18656 19332 18701 19360
rect 18656 19320 18662 19332
rect 18877 19329 18889 19363
rect 18923 19360 18935 19363
rect 19978 19360 19984 19372
rect 18923 19332 19984 19360
rect 18923 19329 18935 19332
rect 18877 19323 18935 19329
rect 19978 19320 19984 19332
rect 20036 19320 20042 19372
rect 20530 19360 20536 19372
rect 20491 19332 20536 19360
rect 20530 19320 20536 19332
rect 20588 19320 20594 19372
rect 15930 19292 15936 19304
rect 11624 19264 11836 19292
rect 15891 19264 15936 19292
rect 15930 19252 15936 19264
rect 15988 19252 15994 19304
rect 17865 19295 17923 19301
rect 17865 19261 17877 19295
rect 17911 19261 17923 19295
rect 17865 19255 17923 19261
rect 10778 19224 10784 19236
rect 8260 19196 8340 19224
rect 8404 19196 8892 19224
rect 10691 19196 10784 19224
rect 8260 19184 8266 19196
rect 8404 19156 8432 19196
rect 8570 19156 8576 19168
rect 8128 19128 8432 19156
rect 8531 19128 8576 19156
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 8864 19156 8892 19196
rect 10778 19184 10784 19196
rect 10836 19224 10842 19236
rect 14918 19224 14924 19236
rect 10836 19196 14924 19224
rect 10836 19184 10842 19196
rect 14918 19184 14924 19196
rect 14976 19184 14982 19236
rect 16758 19184 16764 19236
rect 16816 19224 16822 19236
rect 17310 19224 17316 19236
rect 16816 19196 17316 19224
rect 16816 19184 16822 19196
rect 17310 19184 17316 19196
rect 17368 19184 17374 19236
rect 17880 19224 17908 19255
rect 17954 19252 17960 19304
rect 18012 19292 18018 19304
rect 19889 19295 19947 19301
rect 19889 19292 19901 19295
rect 18012 19264 19901 19292
rect 18012 19252 18018 19264
rect 19889 19261 19901 19264
rect 19935 19261 19947 19295
rect 19889 19255 19947 19261
rect 20254 19252 20260 19304
rect 20312 19292 20318 19304
rect 20640 19292 20668 19400
rect 20717 19397 20729 19400
rect 20763 19397 20775 19431
rect 20717 19391 20775 19397
rect 20806 19388 20812 19440
rect 20864 19428 20870 19440
rect 20901 19431 20959 19437
rect 20901 19428 20913 19431
rect 20864 19400 20913 19428
rect 20864 19388 20870 19400
rect 20901 19397 20913 19400
rect 20947 19397 20959 19431
rect 20901 19391 20959 19397
rect 22097 19363 22155 19369
rect 22097 19329 22109 19363
rect 22143 19360 22155 19363
rect 22370 19360 22376 19372
rect 22143 19332 22376 19360
rect 22143 19329 22155 19332
rect 22097 19323 22155 19329
rect 22370 19320 22376 19332
rect 22428 19320 22434 19372
rect 22554 19360 22560 19372
rect 22515 19332 22560 19360
rect 22554 19320 22560 19332
rect 22612 19320 22618 19372
rect 22646 19320 22652 19372
rect 22704 19360 22710 19372
rect 22704 19332 22749 19360
rect 22704 19320 22710 19332
rect 20312 19264 20668 19292
rect 22848 19292 22876 19468
rect 22940 19468 26884 19496
rect 22940 19369 22968 19468
rect 26878 19456 26884 19468
rect 26936 19456 26942 19508
rect 27522 19456 27528 19508
rect 27580 19496 27586 19508
rect 30006 19496 30012 19508
rect 27580 19468 29040 19496
rect 27580 19456 27586 19468
rect 23474 19428 23480 19440
rect 23216 19400 23480 19428
rect 23216 19369 23244 19400
rect 23474 19388 23480 19400
rect 23532 19388 23538 19440
rect 25774 19388 25780 19440
rect 25832 19428 25838 19440
rect 29012 19437 29040 19468
rect 29104 19468 30012 19496
rect 29104 19437 29132 19468
rect 30006 19456 30012 19468
rect 30064 19456 30070 19508
rect 32674 19456 32680 19508
rect 32732 19496 32738 19508
rect 35526 19496 35532 19508
rect 32732 19468 35296 19496
rect 35487 19468 35532 19496
rect 32732 19456 32738 19468
rect 26237 19431 26295 19437
rect 26237 19428 26249 19431
rect 25832 19400 26249 19428
rect 25832 19388 25838 19400
rect 26237 19397 26249 19400
rect 26283 19397 26295 19431
rect 26237 19391 26295 19397
rect 28997 19431 29055 19437
rect 28997 19397 29009 19431
rect 29043 19397 29055 19431
rect 28997 19391 29055 19397
rect 29089 19431 29147 19437
rect 29089 19397 29101 19431
rect 29135 19397 29147 19431
rect 29089 19391 29147 19397
rect 30193 19431 30251 19437
rect 30193 19397 30205 19431
rect 30239 19428 30251 19431
rect 32306 19428 32312 19440
rect 30239 19400 32312 19428
rect 30239 19397 30251 19400
rect 30193 19391 30251 19397
rect 22925 19363 22983 19369
rect 22925 19329 22937 19363
rect 22971 19329 22983 19363
rect 22925 19323 22983 19329
rect 23201 19363 23259 19369
rect 23201 19329 23213 19363
rect 23247 19329 23259 19363
rect 23382 19360 23388 19372
rect 23343 19332 23388 19360
rect 23201 19323 23259 19329
rect 23382 19320 23388 19332
rect 23440 19320 23446 19372
rect 24302 19360 24308 19372
rect 23492 19332 24308 19360
rect 23492 19292 23520 19332
rect 24302 19320 24308 19332
rect 24360 19320 24366 19372
rect 24397 19363 24455 19369
rect 24397 19329 24409 19363
rect 24443 19360 24455 19363
rect 24946 19360 24952 19372
rect 24443 19332 24952 19360
rect 24443 19329 24455 19332
rect 24397 19323 24455 19329
rect 24946 19320 24952 19332
rect 25004 19320 25010 19372
rect 25406 19360 25412 19372
rect 25148 19332 25412 19360
rect 22848 19264 23520 19292
rect 24673 19295 24731 19301
rect 20312 19252 20318 19264
rect 24673 19261 24685 19295
rect 24719 19292 24731 19295
rect 25038 19292 25044 19304
rect 24719 19264 25044 19292
rect 24719 19261 24731 19264
rect 24673 19255 24731 19261
rect 25038 19252 25044 19264
rect 25096 19252 25102 19304
rect 22278 19224 22284 19236
rect 17880 19196 22284 19224
rect 22278 19184 22284 19196
rect 22336 19184 22342 19236
rect 22830 19184 22836 19236
rect 22888 19224 22894 19236
rect 23382 19224 23388 19236
rect 22888 19196 23388 19224
rect 22888 19184 22894 19196
rect 23382 19184 23388 19196
rect 23440 19184 23446 19236
rect 24949 19227 25007 19233
rect 24949 19193 24961 19227
rect 24995 19224 25007 19227
rect 25148 19224 25176 19332
rect 25406 19320 25412 19332
rect 25464 19320 25470 19372
rect 26050 19360 26056 19372
rect 26011 19332 26056 19360
rect 26050 19320 26056 19332
rect 26108 19320 26114 19372
rect 26326 19360 26332 19372
rect 26287 19332 26332 19360
rect 26326 19320 26332 19332
rect 26384 19320 26390 19372
rect 26418 19320 26424 19372
rect 26476 19360 26482 19372
rect 26476 19332 26521 19360
rect 26476 19320 26482 19332
rect 26878 19320 26884 19372
rect 26936 19360 26942 19372
rect 27157 19363 27215 19369
rect 27157 19360 27169 19363
rect 26936 19332 27169 19360
rect 26936 19320 26942 19332
rect 27157 19329 27169 19332
rect 27203 19329 27215 19363
rect 27617 19363 27675 19369
rect 27617 19360 27629 19363
rect 27157 19323 27215 19329
rect 27264 19332 27629 19360
rect 27062 19252 27068 19304
rect 27120 19292 27126 19304
rect 27264 19292 27292 19332
rect 27617 19329 27629 19332
rect 27663 19329 27675 19363
rect 27617 19323 27675 19329
rect 27893 19363 27951 19369
rect 27893 19329 27905 19363
rect 27939 19360 27951 19363
rect 28721 19363 28779 19369
rect 28721 19360 28733 19363
rect 27939 19332 28733 19360
rect 27939 19329 27951 19332
rect 27893 19323 27951 19329
rect 28721 19329 28733 19332
rect 28767 19329 28779 19363
rect 28721 19323 28779 19329
rect 27120 19264 27292 19292
rect 28736 19292 28764 19323
rect 28810 19320 28816 19372
rect 28868 19360 28874 19372
rect 28868 19332 28913 19360
rect 28868 19320 28874 19332
rect 28902 19292 28908 19304
rect 28736 19264 28908 19292
rect 27120 19252 27126 19264
rect 28902 19252 28908 19264
rect 28960 19252 28966 19304
rect 24995 19196 25176 19224
rect 29012 19224 29040 19391
rect 32306 19388 32312 19400
rect 32364 19388 32370 19440
rect 32861 19431 32919 19437
rect 32861 19397 32873 19431
rect 32907 19428 32919 19431
rect 33502 19428 33508 19440
rect 32907 19400 33508 19428
rect 32907 19397 32919 19400
rect 32861 19391 32919 19397
rect 33502 19388 33508 19400
rect 33560 19388 33566 19440
rect 34422 19388 34428 19440
rect 34480 19428 34486 19440
rect 35158 19428 35164 19440
rect 34480 19400 35164 19428
rect 34480 19388 34486 19400
rect 35158 19388 35164 19400
rect 35216 19388 35222 19440
rect 35268 19437 35296 19468
rect 35526 19456 35532 19468
rect 35584 19456 35590 19508
rect 35253 19431 35311 19437
rect 35253 19397 35265 19431
rect 35299 19428 35311 19431
rect 37642 19428 37648 19440
rect 35299 19400 37648 19428
rect 35299 19397 35311 19400
rect 35253 19391 35311 19397
rect 37642 19388 37648 19400
rect 37700 19388 37706 19440
rect 29270 19369 29276 19372
rect 29227 19363 29276 19369
rect 29227 19329 29239 19363
rect 29273 19329 29276 19363
rect 29227 19323 29276 19329
rect 29270 19320 29276 19323
rect 29328 19320 29334 19372
rect 29822 19360 29828 19372
rect 29880 19369 29886 19372
rect 29790 19332 29828 19360
rect 29822 19320 29828 19332
rect 29880 19323 29890 19369
rect 29918 19363 29976 19369
rect 29918 19329 29930 19363
rect 29964 19360 29976 19363
rect 30006 19360 30012 19372
rect 29964 19332 30012 19360
rect 29964 19329 29976 19332
rect 29918 19323 29976 19329
rect 29880 19320 29886 19323
rect 30006 19320 30012 19332
rect 30064 19320 30070 19372
rect 30101 19363 30159 19369
rect 30101 19329 30113 19363
rect 30147 19329 30159 19363
rect 30282 19360 30288 19372
rect 30340 19369 30346 19372
rect 30248 19332 30288 19360
rect 30101 19323 30159 19329
rect 30116 19224 30144 19323
rect 30282 19320 30288 19332
rect 30340 19323 30348 19369
rect 30340 19320 30346 19323
rect 30742 19320 30748 19372
rect 30800 19360 30806 19372
rect 32674 19360 32680 19372
rect 30800 19332 32680 19360
rect 30800 19320 30806 19332
rect 32674 19320 32680 19332
rect 32732 19360 32738 19372
rect 33045 19363 33103 19369
rect 33045 19360 33057 19363
rect 32732 19332 33057 19360
rect 32732 19320 32738 19332
rect 33045 19329 33057 19332
rect 33091 19329 33103 19363
rect 33045 19323 33103 19329
rect 33137 19363 33195 19369
rect 33137 19329 33149 19363
rect 33183 19334 33195 19363
rect 33183 19329 33217 19334
rect 33137 19323 33217 19329
rect 33152 19306 33217 19323
rect 33318 19320 33324 19372
rect 33376 19360 33382 19372
rect 33376 19332 34836 19360
rect 33376 19320 33382 19332
rect 32950 19252 32956 19304
rect 33008 19292 33014 19304
rect 33152 19292 33180 19306
rect 33008 19264 33180 19292
rect 34808 19292 34836 19332
rect 34882 19320 34888 19372
rect 34940 19360 34946 19372
rect 35066 19369 35072 19372
rect 35033 19363 35072 19369
rect 34940 19332 34985 19360
rect 34940 19320 34946 19332
rect 35033 19329 35045 19363
rect 35033 19323 35072 19329
rect 35066 19320 35072 19323
rect 35124 19320 35130 19372
rect 35391 19363 35449 19369
rect 35391 19360 35403 19363
rect 35176 19332 35403 19360
rect 35176 19304 35204 19332
rect 35391 19329 35403 19332
rect 35437 19360 35449 19363
rect 35526 19360 35532 19372
rect 35437 19332 35532 19360
rect 35437 19329 35449 19332
rect 35391 19323 35449 19329
rect 35526 19320 35532 19332
rect 35584 19320 35590 19372
rect 37734 19320 37740 19372
rect 37792 19360 37798 19372
rect 37829 19363 37887 19369
rect 37829 19360 37841 19363
rect 37792 19332 37841 19360
rect 37792 19320 37798 19332
rect 37829 19329 37841 19332
rect 37875 19329 37887 19363
rect 38102 19360 38108 19372
rect 38063 19332 38108 19360
rect 37829 19323 37887 19329
rect 38102 19320 38108 19332
rect 38160 19320 38166 19372
rect 34808 19264 35112 19292
rect 33008 19252 33014 19264
rect 29012 19196 30144 19224
rect 24995 19193 25007 19196
rect 24949 19187 25007 19193
rect 31754 19184 31760 19236
rect 31812 19224 31818 19236
rect 34974 19224 34980 19236
rect 31812 19196 34980 19224
rect 31812 19184 31818 19196
rect 34974 19184 34980 19196
rect 35032 19184 35038 19236
rect 35084 19224 35112 19264
rect 35158 19252 35164 19304
rect 35216 19252 35222 19304
rect 36354 19224 36360 19236
rect 35084 19196 36360 19224
rect 36354 19184 36360 19196
rect 36412 19184 36418 19236
rect 9674 19156 9680 19168
rect 8864 19128 9680 19156
rect 9674 19116 9680 19128
rect 9732 19116 9738 19168
rect 12250 19116 12256 19168
rect 12308 19156 12314 19168
rect 18138 19156 18144 19168
rect 12308 19128 18144 19156
rect 12308 19116 12314 19128
rect 18138 19116 18144 19128
rect 18196 19116 18202 19168
rect 18325 19159 18383 19165
rect 18325 19125 18337 19159
rect 18371 19156 18383 19159
rect 18690 19156 18696 19168
rect 18371 19128 18696 19156
rect 18371 19125 18383 19128
rect 18325 19119 18383 19125
rect 18690 19116 18696 19128
rect 18748 19116 18754 19168
rect 18785 19159 18843 19165
rect 18785 19125 18797 19159
rect 18831 19156 18843 19159
rect 20806 19156 20812 19168
rect 18831 19128 20812 19156
rect 18831 19125 18843 19128
rect 18785 19119 18843 19125
rect 20806 19116 20812 19128
rect 20864 19116 20870 19168
rect 24486 19156 24492 19168
rect 24447 19128 24492 19156
rect 24486 19116 24492 19128
rect 24544 19116 24550 19168
rect 26602 19156 26608 19168
rect 26563 19128 26608 19156
rect 26602 19116 26608 19128
rect 26660 19116 26666 19168
rect 28534 19116 28540 19168
rect 28592 19156 28598 19168
rect 29178 19156 29184 19168
rect 28592 19128 29184 19156
rect 28592 19116 28598 19128
rect 29178 19116 29184 19128
rect 29236 19116 29242 19168
rect 29365 19159 29423 19165
rect 29365 19125 29377 19159
rect 29411 19156 29423 19159
rect 29730 19156 29736 19168
rect 29411 19128 29736 19156
rect 29411 19125 29423 19128
rect 29365 19119 29423 19125
rect 29730 19116 29736 19128
rect 29788 19116 29794 19168
rect 30282 19116 30288 19168
rect 30340 19156 30346 19168
rect 30469 19159 30527 19165
rect 30469 19156 30481 19159
rect 30340 19128 30481 19156
rect 30340 19116 30346 19128
rect 30469 19125 30481 19128
rect 30515 19125 30527 19159
rect 30469 19119 30527 19125
rect 32861 19159 32919 19165
rect 32861 19125 32873 19159
rect 32907 19156 32919 19159
rect 33318 19156 33324 19168
rect 32907 19128 33324 19156
rect 32907 19125 32919 19128
rect 32861 19119 32919 19125
rect 33318 19116 33324 19128
rect 33376 19116 33382 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 9950 18952 9956 18964
rect 9911 18924 9956 18952
rect 9950 18912 9956 18924
rect 10008 18912 10014 18964
rect 13265 18955 13323 18961
rect 13265 18952 13277 18955
rect 10060 18924 13277 18952
rect 5626 18884 5632 18896
rect 5539 18856 5632 18884
rect 5626 18844 5632 18856
rect 5684 18884 5690 18896
rect 5684 18856 9260 18884
rect 5684 18844 5690 18856
rect 3970 18776 3976 18828
rect 4028 18816 4034 18828
rect 4249 18819 4307 18825
rect 4249 18816 4261 18819
rect 4028 18788 4261 18816
rect 4028 18776 4034 18788
rect 4249 18785 4261 18788
rect 4295 18785 4307 18819
rect 8113 18819 8171 18825
rect 8113 18816 8125 18819
rect 4249 18779 4307 18785
rect 5828 18788 8125 18816
rect 4264 18748 4292 18779
rect 5828 18760 5856 18788
rect 8113 18785 8125 18788
rect 8159 18816 8171 18819
rect 9122 18816 9128 18828
rect 8159 18788 9128 18816
rect 8159 18785 8171 18788
rect 8113 18779 8171 18785
rect 9122 18776 9128 18788
rect 9180 18776 9186 18828
rect 9232 18816 9260 18856
rect 9306 18844 9312 18896
rect 9364 18884 9370 18896
rect 10060 18884 10088 18924
rect 13265 18921 13277 18924
rect 13311 18952 13323 18955
rect 15381 18955 15439 18961
rect 13311 18924 14320 18952
rect 13311 18921 13323 18924
rect 13265 18915 13323 18921
rect 9364 18856 10088 18884
rect 10152 18856 14228 18884
rect 9364 18844 9370 18856
rect 10152 18816 10180 18856
rect 9232 18788 10180 18816
rect 11422 18776 11428 18828
rect 11480 18816 11486 18828
rect 13081 18819 13139 18825
rect 13081 18816 13093 18819
rect 11480 18788 13093 18816
rect 11480 18776 11486 18788
rect 13081 18785 13093 18788
rect 13127 18785 13139 18819
rect 13081 18779 13139 18785
rect 5810 18748 5816 18760
rect 4264 18720 5816 18748
rect 5810 18708 5816 18720
rect 5868 18708 5874 18760
rect 6454 18748 6460 18760
rect 6415 18720 6460 18748
rect 6454 18708 6460 18720
rect 6512 18708 6518 18760
rect 6549 18751 6607 18757
rect 6549 18717 6561 18751
rect 6595 18748 6607 18751
rect 7558 18748 7564 18760
rect 6595 18720 7564 18748
rect 6595 18717 6607 18720
rect 6549 18711 6607 18717
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 9401 18751 9459 18757
rect 9401 18717 9413 18751
rect 9447 18748 9459 18751
rect 9490 18748 9496 18760
rect 9447 18720 9496 18748
rect 9447 18717 9459 18720
rect 9401 18711 9459 18717
rect 9490 18708 9496 18720
rect 9548 18708 9554 18760
rect 9766 18748 9772 18760
rect 9727 18720 9772 18748
rect 9766 18708 9772 18720
rect 9824 18748 9830 18760
rect 10410 18748 10416 18760
rect 9824 18720 10416 18748
rect 9824 18708 9830 18720
rect 10410 18708 10416 18720
rect 10468 18708 10474 18760
rect 13265 18751 13323 18757
rect 13265 18717 13277 18751
rect 13311 18748 13323 18751
rect 13354 18748 13360 18760
rect 13311 18720 13360 18748
rect 13311 18717 13323 18720
rect 13265 18711 13323 18717
rect 13354 18708 13360 18720
rect 13412 18708 13418 18760
rect 4516 18683 4574 18689
rect 4516 18649 4528 18683
rect 4562 18680 4574 18683
rect 5074 18680 5080 18692
rect 4562 18652 5080 18680
rect 4562 18649 4574 18652
rect 4516 18643 4574 18649
rect 5074 18640 5080 18652
rect 5132 18640 5138 18692
rect 6822 18680 6828 18692
rect 6783 18652 6828 18680
rect 6822 18640 6828 18652
rect 6880 18640 6886 18692
rect 6917 18683 6975 18689
rect 6917 18649 6929 18683
rect 6963 18680 6975 18683
rect 7190 18680 7196 18692
rect 6963 18652 7196 18680
rect 6963 18649 6975 18652
rect 6917 18643 6975 18649
rect 7190 18640 7196 18652
rect 7248 18640 7254 18692
rect 7374 18680 7380 18692
rect 7335 18652 7380 18680
rect 7374 18640 7380 18652
rect 7432 18640 7438 18692
rect 8386 18640 8392 18692
rect 8444 18680 8450 18692
rect 9585 18683 9643 18689
rect 9585 18680 9597 18683
rect 8444 18652 9597 18680
rect 8444 18640 8450 18652
rect 9585 18649 9597 18652
rect 9631 18649 9643 18683
rect 9585 18643 9643 18649
rect 9677 18683 9735 18689
rect 9677 18649 9689 18683
rect 9723 18680 9735 18683
rect 10778 18680 10784 18692
rect 9723 18652 10784 18680
rect 9723 18649 9735 18652
rect 9677 18643 9735 18649
rect 10778 18640 10784 18652
rect 10836 18640 10842 18692
rect 12434 18640 12440 18692
rect 12492 18680 12498 18692
rect 12989 18683 13047 18689
rect 12989 18680 13001 18683
rect 12492 18652 13001 18680
rect 12492 18640 12498 18652
rect 12989 18649 13001 18652
rect 13035 18680 13047 18683
rect 13078 18680 13084 18692
rect 13035 18652 13084 18680
rect 13035 18649 13047 18652
rect 12989 18643 13047 18649
rect 13078 18640 13084 18652
rect 13136 18640 13142 18692
rect 14200 18680 14228 18856
rect 14292 18757 14320 18924
rect 15381 18921 15393 18955
rect 15427 18952 15439 18955
rect 15654 18952 15660 18964
rect 15427 18924 15660 18952
rect 15427 18921 15439 18924
rect 15381 18915 15439 18921
rect 15654 18912 15660 18924
rect 15712 18912 15718 18964
rect 17954 18952 17960 18964
rect 15764 18924 17540 18952
rect 17915 18924 17960 18952
rect 15470 18844 15476 18896
rect 15528 18884 15534 18896
rect 15764 18884 15792 18924
rect 15528 18856 15792 18884
rect 15528 18844 15534 18856
rect 15838 18844 15844 18896
rect 15896 18884 15902 18896
rect 17512 18884 17540 18924
rect 17954 18912 17960 18924
rect 18012 18912 18018 18964
rect 18138 18912 18144 18964
rect 18196 18952 18202 18964
rect 19150 18952 19156 18964
rect 18196 18924 19156 18952
rect 18196 18912 18202 18924
rect 19150 18912 19156 18924
rect 19208 18912 19214 18964
rect 20622 18912 20628 18964
rect 20680 18952 20686 18964
rect 21545 18955 21603 18961
rect 21545 18952 21557 18955
rect 20680 18924 21557 18952
rect 20680 18912 20686 18924
rect 21545 18921 21557 18924
rect 21591 18952 21603 18955
rect 23477 18955 23535 18961
rect 21591 18924 22094 18952
rect 21591 18921 21603 18924
rect 21545 18915 21603 18921
rect 22066 18884 22094 18924
rect 23477 18921 23489 18955
rect 23523 18952 23535 18955
rect 24026 18952 24032 18964
rect 23523 18924 24032 18952
rect 23523 18921 23535 18924
rect 23477 18915 23535 18921
rect 24026 18912 24032 18924
rect 24084 18952 24090 18964
rect 24486 18952 24492 18964
rect 24084 18924 24492 18952
rect 24084 18912 24090 18924
rect 24486 18912 24492 18924
rect 24544 18912 24550 18964
rect 24581 18955 24639 18961
rect 24581 18921 24593 18955
rect 24627 18921 24639 18955
rect 24946 18952 24952 18964
rect 24907 18924 24952 18952
rect 24581 18915 24639 18921
rect 15896 18856 17448 18884
rect 15896 18844 15902 18856
rect 16945 18819 17003 18825
rect 16945 18785 16957 18819
rect 16991 18816 17003 18819
rect 17034 18816 17040 18828
rect 16991 18788 17040 18816
rect 16991 18785 17003 18788
rect 16945 18779 17003 18785
rect 17034 18776 17040 18788
rect 17092 18816 17098 18828
rect 17092 18788 17356 18816
rect 17092 18776 17098 18788
rect 14277 18751 14335 18757
rect 14277 18717 14289 18751
rect 14323 18717 14335 18751
rect 14277 18711 14335 18717
rect 14918 18708 14924 18760
rect 14976 18748 14982 18760
rect 15289 18751 15347 18757
rect 15289 18748 15301 18751
rect 14976 18720 15301 18748
rect 14976 18708 14982 18720
rect 15289 18717 15301 18720
rect 15335 18717 15347 18751
rect 17126 18748 17132 18760
rect 17087 18720 17132 18748
rect 15289 18711 15347 18717
rect 17126 18708 17132 18720
rect 17184 18708 17190 18760
rect 17221 18751 17279 18757
rect 17221 18717 17233 18751
rect 17267 18717 17279 18751
rect 17221 18711 17279 18717
rect 17236 18680 17264 18711
rect 14200 18652 17264 18680
rect 17328 18680 17356 18788
rect 17420 18757 17448 18856
rect 17512 18856 20024 18884
rect 22066 18856 23704 18884
rect 17512 18757 17540 18856
rect 19996 18828 20024 18856
rect 18325 18819 18383 18825
rect 18325 18816 18337 18819
rect 17604 18788 18337 18816
rect 17405 18751 17463 18757
rect 17405 18717 17417 18751
rect 17451 18717 17463 18751
rect 17405 18711 17463 18717
rect 17497 18751 17555 18757
rect 17497 18717 17509 18751
rect 17543 18717 17555 18751
rect 17497 18711 17555 18717
rect 17604 18680 17632 18788
rect 18325 18785 18337 18788
rect 18371 18785 18383 18819
rect 18325 18779 18383 18785
rect 18414 18776 18420 18828
rect 18472 18816 18478 18828
rect 18472 18788 18517 18816
rect 18472 18776 18478 18788
rect 19978 18776 19984 18828
rect 20036 18816 20042 18828
rect 20349 18819 20407 18825
rect 20349 18816 20361 18819
rect 20036 18788 20361 18816
rect 20036 18776 20042 18788
rect 20349 18785 20361 18788
rect 20395 18785 20407 18819
rect 20349 18779 20407 18785
rect 21542 18776 21548 18828
rect 21600 18816 21606 18828
rect 21637 18819 21695 18825
rect 21637 18816 21649 18819
rect 21600 18788 21649 18816
rect 21600 18776 21606 18788
rect 21637 18785 21649 18788
rect 21683 18816 21695 18819
rect 23474 18816 23480 18828
rect 21683 18788 23480 18816
rect 21683 18785 21695 18788
rect 21637 18779 21695 18785
rect 23474 18776 23480 18788
rect 23532 18776 23538 18828
rect 18141 18751 18199 18757
rect 18141 18717 18153 18751
rect 18187 18717 18199 18751
rect 18141 18711 18199 18717
rect 21821 18751 21879 18757
rect 21821 18717 21833 18751
rect 21867 18748 21879 18751
rect 21910 18748 21916 18760
rect 21867 18720 21916 18748
rect 21867 18717 21879 18720
rect 21821 18711 21879 18717
rect 17328 18652 17632 18680
rect 18156 18680 18184 18711
rect 21910 18708 21916 18720
rect 21968 18708 21974 18760
rect 22462 18748 22468 18760
rect 22423 18720 22468 18748
rect 22462 18708 22468 18720
rect 22520 18708 22526 18760
rect 23676 18757 23704 18856
rect 23934 18816 23940 18828
rect 23847 18788 23940 18816
rect 23934 18776 23940 18788
rect 23992 18816 23998 18828
rect 24596 18816 24624 18915
rect 24946 18912 24952 18924
rect 25004 18912 25010 18964
rect 29178 18912 29184 18964
rect 29236 18952 29242 18964
rect 29730 18952 29736 18964
rect 29236 18924 29736 18952
rect 29236 18912 29242 18924
rect 29730 18912 29736 18924
rect 29788 18912 29794 18964
rect 33413 18955 33471 18961
rect 33413 18921 33425 18955
rect 33459 18952 33471 18955
rect 33502 18952 33508 18964
rect 33459 18924 33508 18952
rect 33459 18921 33471 18924
rect 33413 18915 33471 18921
rect 33502 18912 33508 18924
rect 33560 18912 33566 18964
rect 28902 18844 28908 18896
rect 28960 18884 28966 18896
rect 29822 18884 29828 18896
rect 28960 18856 29828 18884
rect 28960 18844 28966 18856
rect 29822 18844 29828 18856
rect 29880 18844 29886 18896
rect 30466 18844 30472 18896
rect 30524 18884 30530 18896
rect 31294 18884 31300 18896
rect 30524 18856 31300 18884
rect 30524 18844 30530 18856
rect 31294 18844 31300 18856
rect 31352 18844 31358 18896
rect 32217 18887 32275 18893
rect 32217 18853 32229 18887
rect 32263 18884 32275 18887
rect 32306 18884 32312 18896
rect 32263 18856 32312 18884
rect 32263 18853 32275 18856
rect 32217 18847 32275 18853
rect 32306 18844 32312 18856
rect 32364 18884 32370 18896
rect 32950 18884 32956 18896
rect 32364 18856 32956 18884
rect 32364 18844 32370 18856
rect 32950 18844 32956 18856
rect 33008 18844 33014 18896
rect 33042 18844 33048 18896
rect 33100 18884 33106 18896
rect 33226 18884 33232 18896
rect 33100 18856 33232 18884
rect 33100 18844 33106 18856
rect 33226 18844 33232 18856
rect 33284 18844 33290 18896
rect 34882 18844 34888 18896
rect 34940 18884 34946 18896
rect 36078 18884 36084 18896
rect 34940 18856 36084 18884
rect 34940 18844 34946 18856
rect 36078 18844 36084 18856
rect 36136 18844 36142 18896
rect 25866 18816 25872 18828
rect 23992 18788 24624 18816
rect 25827 18788 25872 18816
rect 23992 18776 23998 18788
rect 25866 18776 25872 18788
rect 25924 18776 25930 18828
rect 27890 18776 27896 18828
rect 27948 18816 27954 18828
rect 30006 18816 30012 18828
rect 27948 18788 30012 18816
rect 27948 18776 27954 18788
rect 30006 18776 30012 18788
rect 30064 18776 30070 18828
rect 33152 18788 35480 18816
rect 22649 18751 22707 18757
rect 22649 18717 22661 18751
rect 22695 18717 22707 18751
rect 22649 18711 22707 18717
rect 23661 18751 23719 18757
rect 23661 18717 23673 18751
rect 23707 18717 23719 18751
rect 23842 18748 23848 18760
rect 23803 18720 23848 18748
rect 23661 18711 23719 18717
rect 18506 18680 18512 18692
rect 18156 18652 18512 18680
rect 6086 18572 6092 18624
rect 6144 18612 6150 18624
rect 6273 18615 6331 18621
rect 6273 18612 6285 18615
rect 6144 18584 6285 18612
rect 6144 18572 6150 18584
rect 6273 18581 6285 18584
rect 6319 18581 6331 18615
rect 13446 18612 13452 18624
rect 13407 18584 13452 18612
rect 6273 18575 6331 18581
rect 13446 18572 13452 18584
rect 13504 18572 13510 18624
rect 14274 18572 14280 18624
rect 14332 18612 14338 18624
rect 14369 18615 14427 18621
rect 14369 18612 14381 18615
rect 14332 18584 14381 18612
rect 14332 18572 14338 18584
rect 14369 18581 14381 18584
rect 14415 18581 14427 18615
rect 17236 18612 17264 18652
rect 18506 18640 18512 18652
rect 18564 18640 18570 18692
rect 21358 18640 21364 18692
rect 21416 18680 21422 18692
rect 21545 18683 21603 18689
rect 21545 18680 21557 18683
rect 21416 18652 21557 18680
rect 21416 18640 21422 18652
rect 21545 18649 21557 18652
rect 21591 18649 21603 18683
rect 22664 18680 22692 18711
rect 21545 18643 21603 18649
rect 22020 18652 22692 18680
rect 18598 18612 18604 18624
rect 17236 18584 18604 18612
rect 14369 18575 14427 18581
rect 18598 18572 18604 18584
rect 18656 18572 18662 18624
rect 19797 18615 19855 18621
rect 19797 18581 19809 18615
rect 19843 18612 19855 18615
rect 19978 18612 19984 18624
rect 19843 18584 19984 18612
rect 19843 18581 19855 18584
rect 19797 18575 19855 18581
rect 19978 18572 19984 18584
rect 20036 18572 20042 18624
rect 20162 18612 20168 18624
rect 20123 18584 20168 18612
rect 20162 18572 20168 18584
rect 20220 18572 20226 18624
rect 20257 18615 20315 18621
rect 20257 18581 20269 18615
rect 20303 18612 20315 18615
rect 20346 18612 20352 18624
rect 20303 18584 20352 18612
rect 20303 18581 20315 18584
rect 20257 18575 20315 18581
rect 20346 18572 20352 18584
rect 20404 18572 20410 18624
rect 22020 18621 22048 18652
rect 22005 18615 22063 18621
rect 22005 18581 22017 18615
rect 22051 18581 22063 18615
rect 22554 18612 22560 18624
rect 22515 18584 22560 18612
rect 22005 18575 22063 18581
rect 22554 18572 22560 18584
rect 22612 18572 22618 18624
rect 23676 18612 23704 18711
rect 23842 18708 23848 18720
rect 23900 18708 23906 18760
rect 24581 18751 24639 18757
rect 24581 18717 24593 18751
rect 24627 18717 24639 18751
rect 24581 18711 24639 18717
rect 24673 18751 24731 18757
rect 24673 18717 24685 18751
rect 24719 18748 24731 18751
rect 29362 18748 29368 18760
rect 24719 18720 29368 18748
rect 24719 18717 24731 18720
rect 24673 18711 24731 18717
rect 23860 18680 23888 18708
rect 24596 18680 24624 18711
rect 23860 18652 24624 18680
rect 24688 18612 24716 18711
rect 29362 18708 29368 18720
rect 29420 18708 29426 18760
rect 30834 18748 30840 18760
rect 30795 18720 30840 18748
rect 30834 18708 30840 18720
rect 30892 18708 30898 18760
rect 31297 18751 31355 18757
rect 31297 18717 31309 18751
rect 31343 18748 31355 18751
rect 31386 18748 31392 18760
rect 31343 18720 31392 18748
rect 31343 18717 31355 18720
rect 31297 18711 31355 18717
rect 26136 18683 26194 18689
rect 26136 18649 26148 18683
rect 26182 18680 26194 18683
rect 28718 18680 28724 18692
rect 26182 18652 28724 18680
rect 26182 18649 26194 18652
rect 26136 18643 26194 18649
rect 28718 18640 28724 18652
rect 28776 18640 28782 18692
rect 30006 18640 30012 18692
rect 30064 18680 30070 18692
rect 31312 18680 31340 18711
rect 31386 18708 31392 18720
rect 31444 18708 31450 18760
rect 31570 18708 31576 18760
rect 31628 18748 31634 18760
rect 31757 18751 31815 18757
rect 31757 18748 31769 18751
rect 31628 18720 31769 18748
rect 31628 18708 31634 18720
rect 31757 18717 31769 18720
rect 31803 18717 31815 18751
rect 31757 18711 31815 18717
rect 31938 18708 31944 18760
rect 31996 18748 32002 18760
rect 32033 18751 32091 18757
rect 32033 18748 32045 18751
rect 31996 18720 32045 18748
rect 31996 18708 32002 18720
rect 32033 18717 32045 18720
rect 32079 18717 32091 18751
rect 32033 18711 32091 18717
rect 32490 18708 32496 18760
rect 32548 18748 32554 18760
rect 32769 18751 32827 18757
rect 32769 18748 32781 18751
rect 32548 18720 32781 18748
rect 32548 18708 32554 18720
rect 32769 18717 32781 18720
rect 32815 18717 32827 18751
rect 32769 18711 32827 18717
rect 32917 18751 32975 18757
rect 32917 18717 32929 18751
rect 32963 18748 32975 18751
rect 33152 18748 33180 18788
rect 32963 18720 33180 18748
rect 32963 18717 32975 18720
rect 32917 18711 32975 18717
rect 33226 18708 33232 18760
rect 33284 18757 33290 18760
rect 33284 18748 33292 18757
rect 33284 18720 33329 18748
rect 33284 18711 33292 18720
rect 33284 18708 33290 18711
rect 34790 18708 34796 18760
rect 34848 18748 34854 18760
rect 35058 18751 35116 18757
rect 35058 18748 35070 18751
rect 34848 18720 35070 18748
rect 34848 18708 34854 18720
rect 35058 18717 35070 18720
rect 35104 18717 35116 18751
rect 35058 18711 35116 18717
rect 35158 18708 35164 18760
rect 35216 18748 35222 18760
rect 35342 18748 35348 18760
rect 35216 18720 35261 18748
rect 35303 18720 35348 18748
rect 35216 18708 35222 18720
rect 35342 18708 35348 18720
rect 35400 18708 35406 18760
rect 35452 18757 35480 18788
rect 35437 18751 35495 18757
rect 35437 18717 35449 18751
rect 35483 18717 35495 18751
rect 35437 18711 35495 18717
rect 33045 18683 33103 18689
rect 33045 18680 33057 18683
rect 30064 18652 31340 18680
rect 32876 18652 33057 18680
rect 30064 18640 30070 18652
rect 32876 18624 32904 18652
rect 33045 18649 33057 18652
rect 33091 18649 33103 18683
rect 33045 18643 33103 18649
rect 33137 18683 33195 18689
rect 33137 18649 33149 18683
rect 33183 18680 33195 18683
rect 33318 18680 33324 18692
rect 33183 18652 33324 18680
rect 33183 18649 33195 18652
rect 33137 18643 33195 18649
rect 33318 18640 33324 18652
rect 33376 18680 33382 18692
rect 33594 18680 33600 18692
rect 33376 18652 33600 18680
rect 33376 18640 33382 18652
rect 33594 18640 33600 18652
rect 33652 18640 33658 18692
rect 33778 18640 33784 18692
rect 33836 18680 33842 18692
rect 35176 18680 35204 18708
rect 33836 18652 35204 18680
rect 35452 18680 35480 18711
rect 35526 18708 35532 18760
rect 35584 18757 35590 18760
rect 35584 18748 35592 18757
rect 36725 18751 36783 18757
rect 35584 18720 35629 18748
rect 35584 18711 35592 18720
rect 36725 18717 36737 18751
rect 36771 18748 36783 18751
rect 36814 18748 36820 18760
rect 36771 18720 36820 18748
rect 36771 18717 36783 18720
rect 36725 18711 36783 18717
rect 35584 18708 35590 18711
rect 36814 18708 36820 18720
rect 36872 18708 36878 18760
rect 36992 18683 37050 18689
rect 35452 18652 36952 18680
rect 33836 18640 33842 18652
rect 23676 18584 24716 18612
rect 26786 18572 26792 18624
rect 26844 18612 26850 18624
rect 27249 18615 27307 18621
rect 27249 18612 27261 18615
rect 26844 18584 27261 18612
rect 26844 18572 26850 18584
rect 27249 18581 27261 18584
rect 27295 18612 27307 18615
rect 30742 18612 30748 18624
rect 27295 18584 30748 18612
rect 27295 18581 27307 18584
rect 27249 18575 27307 18581
rect 30742 18572 30748 18584
rect 30800 18572 30806 18624
rect 32858 18572 32864 18624
rect 32916 18572 32922 18624
rect 32950 18572 32956 18624
rect 33008 18612 33014 18624
rect 34882 18612 34888 18624
rect 33008 18584 34888 18612
rect 33008 18572 33014 18584
rect 34882 18572 34888 18584
rect 34940 18572 34946 18624
rect 35710 18612 35716 18624
rect 35671 18584 35716 18612
rect 35710 18572 35716 18584
rect 35768 18572 35774 18624
rect 36924 18612 36952 18652
rect 36992 18649 37004 18683
rect 37038 18680 37050 18683
rect 37458 18680 37464 18692
rect 37038 18652 37464 18680
rect 37038 18649 37050 18652
rect 36992 18643 37050 18649
rect 37458 18640 37464 18652
rect 37516 18640 37522 18692
rect 37826 18612 37832 18624
rect 36924 18584 37832 18612
rect 37826 18572 37832 18584
rect 37884 18612 37890 18624
rect 38105 18615 38163 18621
rect 38105 18612 38117 18615
rect 37884 18584 38117 18612
rect 37884 18572 37890 18584
rect 38105 18581 38117 18584
rect 38151 18581 38163 18615
rect 38105 18575 38163 18581
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 6454 18368 6460 18420
rect 6512 18408 6518 18420
rect 6917 18411 6975 18417
rect 6917 18408 6929 18411
rect 6512 18380 6929 18408
rect 6512 18368 6518 18380
rect 6917 18377 6929 18380
rect 6963 18377 6975 18411
rect 8754 18408 8760 18420
rect 6917 18371 6975 18377
rect 8128 18380 8760 18408
rect 8128 18340 8156 18380
rect 8754 18368 8760 18380
rect 8812 18368 8818 18420
rect 9306 18408 9312 18420
rect 9267 18380 9312 18408
rect 9306 18368 9312 18380
rect 9364 18368 9370 18420
rect 10226 18368 10232 18420
rect 10284 18368 10290 18420
rect 12250 18368 12256 18420
rect 12308 18408 12314 18420
rect 13081 18411 13139 18417
rect 13081 18408 13093 18411
rect 12308 18380 13093 18408
rect 12308 18368 12314 18380
rect 13081 18377 13093 18380
rect 13127 18377 13139 18411
rect 13081 18371 13139 18377
rect 13173 18411 13231 18417
rect 13173 18377 13185 18411
rect 13219 18408 13231 18411
rect 13909 18411 13967 18417
rect 13909 18408 13921 18411
rect 13219 18380 13921 18408
rect 13219 18377 13231 18380
rect 13173 18371 13231 18377
rect 13909 18377 13921 18380
rect 13955 18377 13967 18411
rect 14274 18408 14280 18420
rect 14235 18380 14280 18408
rect 13909 18371 13967 18377
rect 14274 18368 14280 18380
rect 14332 18368 14338 18420
rect 14369 18411 14427 18417
rect 14369 18377 14381 18411
rect 14415 18408 14427 18411
rect 14415 18380 17908 18408
rect 14415 18377 14427 18380
rect 14369 18371 14427 18377
rect 6840 18312 8156 18340
rect 8196 18343 8254 18349
rect 6840 18281 6868 18312
rect 8196 18309 8208 18343
rect 8242 18340 8254 18343
rect 8570 18340 8576 18352
rect 8242 18312 8576 18340
rect 8242 18309 8254 18312
rect 8196 18303 8254 18309
rect 8570 18300 8576 18312
rect 8628 18300 8634 18352
rect 10244 18340 10272 18368
rect 10060 18312 10272 18340
rect 10321 18343 10379 18349
rect 6825 18275 6883 18281
rect 6825 18241 6837 18275
rect 6871 18241 6883 18275
rect 6825 18235 6883 18241
rect 7009 18275 7067 18281
rect 7009 18241 7021 18275
rect 7055 18272 7067 18275
rect 7098 18272 7104 18284
rect 7055 18244 7104 18272
rect 7055 18241 7067 18244
rect 7009 18235 7067 18241
rect 7098 18232 7104 18244
rect 7156 18232 7162 18284
rect 10060 18281 10088 18312
rect 10321 18309 10333 18343
rect 10367 18340 10379 18343
rect 11422 18340 11428 18352
rect 10367 18312 11428 18340
rect 10367 18309 10379 18312
rect 10321 18303 10379 18309
rect 11422 18300 11428 18312
rect 11480 18300 11486 18352
rect 14734 18340 14740 18352
rect 13280 18312 14740 18340
rect 10045 18275 10103 18281
rect 10045 18241 10057 18275
rect 10091 18241 10103 18275
rect 10045 18235 10103 18241
rect 10229 18275 10287 18281
rect 10229 18241 10241 18275
rect 10275 18241 10287 18275
rect 10410 18272 10416 18284
rect 10371 18244 10416 18272
rect 10229 18235 10287 18241
rect 7926 18204 7932 18216
rect 7887 18176 7932 18204
rect 7926 18164 7932 18176
rect 7984 18164 7990 18216
rect 9674 18164 9680 18216
rect 9732 18204 9738 18216
rect 10244 18204 10272 18235
rect 10410 18232 10416 18244
rect 10468 18232 10474 18284
rect 13280 18213 13308 18312
rect 14734 18300 14740 18312
rect 14792 18300 14798 18352
rect 15930 18300 15936 18352
rect 15988 18340 15994 18352
rect 15988 18312 17632 18340
rect 15988 18300 15994 18312
rect 13446 18232 13452 18284
rect 13504 18272 13510 18284
rect 15289 18275 15347 18281
rect 15289 18272 15301 18275
rect 13504 18244 15301 18272
rect 13504 18232 13510 18244
rect 15289 18241 15301 18244
rect 15335 18241 15347 18275
rect 15289 18235 15347 18241
rect 15378 18232 15384 18284
rect 15436 18272 15442 18284
rect 15473 18275 15531 18281
rect 15473 18272 15485 18275
rect 15436 18244 15485 18272
rect 15436 18232 15442 18244
rect 15473 18241 15485 18244
rect 15519 18241 15531 18275
rect 15473 18235 15531 18241
rect 15565 18275 15623 18281
rect 15565 18241 15577 18275
rect 15611 18272 15623 18275
rect 15838 18272 15844 18284
rect 15611 18244 15844 18272
rect 15611 18241 15623 18244
rect 15565 18235 15623 18241
rect 15838 18232 15844 18244
rect 15896 18232 15902 18284
rect 9732 18176 10272 18204
rect 13265 18207 13323 18213
rect 9732 18164 9738 18176
rect 13265 18173 13277 18207
rect 13311 18173 13323 18207
rect 13265 18167 13323 18173
rect 14553 18207 14611 18213
rect 14553 18173 14565 18207
rect 14599 18204 14611 18207
rect 15194 18204 15200 18216
rect 14599 18176 15200 18204
rect 14599 18173 14611 18176
rect 14553 18167 14611 18173
rect 13354 18096 13360 18148
rect 13412 18136 13418 18148
rect 14568 18136 14596 18167
rect 15194 18164 15200 18176
rect 15252 18204 15258 18216
rect 15948 18204 15976 18300
rect 17034 18232 17040 18284
rect 17092 18272 17098 18284
rect 17129 18275 17187 18281
rect 17129 18272 17141 18275
rect 17092 18244 17141 18272
rect 17092 18232 17098 18244
rect 17129 18241 17141 18244
rect 17175 18241 17187 18275
rect 17129 18235 17187 18241
rect 17310 18232 17316 18284
rect 17368 18272 17374 18284
rect 17405 18275 17463 18281
rect 17405 18272 17417 18275
rect 17368 18244 17417 18272
rect 17368 18232 17374 18244
rect 17405 18241 17417 18244
rect 17451 18272 17463 18275
rect 17494 18272 17500 18284
rect 17451 18244 17500 18272
rect 17451 18241 17463 18244
rect 17405 18235 17463 18241
rect 17494 18232 17500 18244
rect 17552 18232 17558 18284
rect 17604 18281 17632 18312
rect 17589 18275 17647 18281
rect 17589 18241 17601 18275
rect 17635 18241 17647 18275
rect 17589 18235 17647 18241
rect 15252 18176 15976 18204
rect 15252 18164 15258 18176
rect 16666 18164 16672 18216
rect 16724 18204 16730 18216
rect 17221 18207 17279 18213
rect 17221 18204 17233 18207
rect 16724 18176 17233 18204
rect 16724 18164 16730 18176
rect 17221 18173 17233 18176
rect 17267 18173 17279 18207
rect 17880 18204 17908 18380
rect 17954 18368 17960 18420
rect 18012 18408 18018 18420
rect 18509 18411 18567 18417
rect 18509 18408 18521 18411
rect 18012 18380 18521 18408
rect 18012 18368 18018 18380
rect 18432 18272 18460 18380
rect 18509 18377 18521 18380
rect 18555 18377 18567 18411
rect 18509 18371 18567 18377
rect 18601 18411 18659 18417
rect 18601 18377 18613 18411
rect 18647 18408 18659 18411
rect 19337 18411 19395 18417
rect 19337 18408 19349 18411
rect 18647 18380 19349 18408
rect 18647 18377 18659 18380
rect 18601 18371 18659 18377
rect 19337 18377 19349 18380
rect 19383 18377 19395 18411
rect 19337 18371 19395 18377
rect 19797 18411 19855 18417
rect 19797 18377 19809 18411
rect 19843 18408 19855 18411
rect 19978 18408 19984 18420
rect 19843 18380 19984 18408
rect 19843 18377 19855 18380
rect 19797 18371 19855 18377
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 23382 18408 23388 18420
rect 22296 18380 23388 18408
rect 19705 18343 19763 18349
rect 19705 18309 19717 18343
rect 19751 18340 19763 18343
rect 20070 18340 20076 18352
rect 19751 18312 20076 18340
rect 19751 18309 19763 18312
rect 19705 18303 19763 18309
rect 20070 18300 20076 18312
rect 20128 18300 20134 18352
rect 22296 18340 22324 18380
rect 23382 18368 23388 18380
rect 23440 18368 23446 18420
rect 24305 18411 24363 18417
rect 24305 18377 24317 18411
rect 24351 18408 24363 18411
rect 25130 18408 25136 18420
rect 24351 18380 25136 18408
rect 24351 18377 24363 18380
rect 24305 18371 24363 18377
rect 25130 18368 25136 18380
rect 25188 18368 25194 18420
rect 30745 18411 30803 18417
rect 30745 18408 30757 18411
rect 29380 18380 30757 18408
rect 23934 18340 23940 18352
rect 22112 18312 22324 18340
rect 23032 18312 23940 18340
rect 19334 18272 19340 18284
rect 18432 18244 19340 18272
rect 19334 18232 19340 18244
rect 19392 18232 19398 18284
rect 19518 18232 19524 18284
rect 19576 18272 19582 18284
rect 22002 18272 22008 18284
rect 19576 18244 22008 18272
rect 19576 18232 19582 18244
rect 22002 18232 22008 18244
rect 22060 18232 22066 18284
rect 18690 18204 18696 18216
rect 17880 18176 18552 18204
rect 18651 18176 18696 18204
rect 17221 18167 17279 18173
rect 13412 18108 14596 18136
rect 13412 18096 13418 18108
rect 15746 18096 15752 18148
rect 15804 18136 15810 18148
rect 18414 18136 18420 18148
rect 15804 18108 18420 18136
rect 15804 18096 15810 18108
rect 18414 18096 18420 18108
rect 18472 18096 18478 18148
rect 10594 18068 10600 18080
rect 10555 18040 10600 18068
rect 10594 18028 10600 18040
rect 10652 18028 10658 18080
rect 12710 18068 12716 18080
rect 12671 18040 12716 18068
rect 12710 18028 12716 18040
rect 12768 18028 12774 18080
rect 13998 18028 14004 18080
rect 14056 18068 14062 18080
rect 15105 18071 15163 18077
rect 15105 18068 15117 18071
rect 14056 18040 15117 18068
rect 14056 18028 14062 18040
rect 15105 18037 15117 18040
rect 15151 18037 15163 18071
rect 16850 18068 16856 18080
rect 16811 18040 16856 18068
rect 15105 18031 15163 18037
rect 16850 18028 16856 18040
rect 16908 18028 16914 18080
rect 17310 18028 17316 18080
rect 17368 18068 17374 18080
rect 18138 18068 18144 18080
rect 17368 18040 17413 18068
rect 18099 18040 18144 18068
rect 17368 18028 17374 18040
rect 18138 18028 18144 18040
rect 18196 18028 18202 18080
rect 18524 18068 18552 18176
rect 18690 18164 18696 18176
rect 18748 18164 18754 18216
rect 19426 18164 19432 18216
rect 19484 18204 19490 18216
rect 22112 18213 22140 18312
rect 22281 18275 22339 18281
rect 22281 18272 22293 18275
rect 22204 18244 22293 18272
rect 19889 18207 19947 18213
rect 19889 18204 19901 18207
rect 19484 18176 19901 18204
rect 19484 18164 19490 18176
rect 19889 18173 19901 18176
rect 19935 18173 19947 18207
rect 19889 18167 19947 18173
rect 22097 18207 22155 18213
rect 22097 18173 22109 18207
rect 22143 18173 22155 18207
rect 22097 18167 22155 18173
rect 18598 18096 18604 18148
rect 18656 18136 18662 18148
rect 22204 18136 22232 18244
rect 22281 18241 22293 18244
rect 22327 18272 22339 18275
rect 22554 18272 22560 18284
rect 22327 18244 22560 18272
rect 22327 18241 22339 18244
rect 22281 18235 22339 18241
rect 22554 18232 22560 18244
rect 22612 18232 22618 18284
rect 23032 18281 23060 18312
rect 23934 18300 23940 18312
rect 23992 18300 23998 18352
rect 24670 18300 24676 18352
rect 24728 18340 24734 18352
rect 29380 18349 29408 18380
rect 30745 18377 30757 18380
rect 30791 18377 30803 18411
rect 30745 18371 30803 18377
rect 33134 18368 33140 18420
rect 33192 18408 33198 18420
rect 33689 18411 33747 18417
rect 33689 18408 33701 18411
rect 33192 18380 33701 18408
rect 33192 18368 33198 18380
rect 33689 18377 33701 18380
rect 33735 18377 33747 18411
rect 37458 18408 37464 18420
rect 37419 18380 37464 18408
rect 33689 18371 33747 18377
rect 37458 18368 37464 18380
rect 37516 18368 37522 18420
rect 37826 18408 37832 18420
rect 37787 18380 37832 18408
rect 37826 18368 37832 18380
rect 37884 18368 37890 18420
rect 24765 18343 24823 18349
rect 24765 18340 24777 18343
rect 24728 18312 24777 18340
rect 24728 18300 24734 18312
rect 24765 18309 24777 18312
rect 24811 18309 24823 18343
rect 29365 18343 29423 18349
rect 29365 18340 29377 18343
rect 24765 18303 24823 18309
rect 28368 18312 29377 18340
rect 23017 18275 23075 18281
rect 23017 18241 23029 18275
rect 23063 18241 23075 18275
rect 23017 18235 23075 18241
rect 23201 18275 23259 18281
rect 23201 18241 23213 18275
rect 23247 18272 23259 18275
rect 23474 18272 23480 18284
rect 23247 18244 23480 18272
rect 23247 18241 23259 18244
rect 23201 18235 23259 18241
rect 23474 18232 23480 18244
rect 23532 18272 23538 18284
rect 24026 18272 24032 18284
rect 23532 18244 23796 18272
rect 23987 18244 24032 18272
rect 23532 18232 23538 18244
rect 23566 18164 23572 18216
rect 23624 18204 23630 18216
rect 23661 18207 23719 18213
rect 23661 18204 23673 18207
rect 23624 18176 23673 18204
rect 23624 18164 23630 18176
rect 23661 18173 23673 18176
rect 23707 18173 23719 18207
rect 23661 18167 23719 18173
rect 23768 18148 23796 18244
rect 24026 18232 24032 18244
rect 24084 18232 24090 18284
rect 26970 18232 26976 18284
rect 27028 18272 27034 18284
rect 27706 18272 27712 18284
rect 27028 18244 27712 18272
rect 27028 18232 27034 18244
rect 27706 18232 27712 18244
rect 27764 18232 27770 18284
rect 28368 18281 28396 18312
rect 29365 18309 29377 18312
rect 29411 18309 29423 18343
rect 29365 18303 29423 18309
rect 30650 18300 30656 18352
rect 30708 18340 30714 18352
rect 34422 18340 34428 18352
rect 30708 18312 34428 18340
rect 30708 18300 30714 18312
rect 34422 18300 34428 18312
rect 34480 18300 34486 18352
rect 35529 18343 35587 18349
rect 35529 18309 35541 18343
rect 35575 18340 35587 18343
rect 37734 18340 37740 18352
rect 35575 18312 37740 18340
rect 35575 18309 35587 18312
rect 35529 18303 35587 18309
rect 37734 18300 37740 18312
rect 37792 18340 37798 18352
rect 37921 18343 37979 18349
rect 37921 18340 37933 18343
rect 37792 18312 37933 18340
rect 37792 18300 37798 18312
rect 37921 18309 37933 18312
rect 37967 18309 37979 18343
rect 37921 18303 37979 18309
rect 28353 18275 28411 18281
rect 28353 18241 28365 18275
rect 28399 18241 28411 18275
rect 29181 18275 29239 18281
rect 29181 18272 29193 18275
rect 28353 18235 28411 18241
rect 28460 18244 29193 18272
rect 24118 18164 24124 18216
rect 24176 18204 24182 18216
rect 25593 18207 25651 18213
rect 24176 18176 24221 18204
rect 24176 18164 24182 18176
rect 25593 18173 25605 18207
rect 25639 18204 25651 18207
rect 25774 18204 25780 18216
rect 25639 18176 25780 18204
rect 25639 18173 25651 18176
rect 25593 18167 25651 18173
rect 25774 18164 25780 18176
rect 25832 18164 25838 18216
rect 27154 18164 27160 18216
rect 27212 18204 27218 18216
rect 28261 18207 28319 18213
rect 28261 18204 28273 18207
rect 27212 18176 28273 18204
rect 27212 18164 27218 18176
rect 28261 18173 28273 18176
rect 28307 18204 28319 18207
rect 28460 18204 28488 18244
rect 29181 18241 29193 18244
rect 29227 18241 29239 18275
rect 30558 18272 30564 18284
rect 30519 18244 30564 18272
rect 29181 18235 29239 18241
rect 30558 18232 30564 18244
rect 30616 18232 30622 18284
rect 30745 18275 30803 18281
rect 30745 18272 30757 18275
rect 30668 18244 30757 18272
rect 30668 18216 30696 18244
rect 30745 18241 30757 18244
rect 30791 18241 30803 18275
rect 30745 18235 30803 18241
rect 33321 18275 33379 18281
rect 33321 18241 33333 18275
rect 33367 18272 33379 18275
rect 33410 18272 33416 18284
rect 33367 18244 33416 18272
rect 33367 18241 33379 18244
rect 33321 18235 33379 18241
rect 33410 18232 33416 18244
rect 33468 18232 33474 18284
rect 33505 18275 33563 18281
rect 33505 18241 33517 18275
rect 33551 18272 33563 18275
rect 33686 18272 33692 18284
rect 33551 18244 33692 18272
rect 33551 18241 33563 18244
rect 33505 18235 33563 18241
rect 33686 18232 33692 18244
rect 33744 18232 33750 18284
rect 35710 18272 35716 18284
rect 35671 18244 35716 18272
rect 35710 18232 35716 18244
rect 35768 18232 35774 18284
rect 35802 18232 35808 18284
rect 35860 18272 35866 18284
rect 36081 18275 36139 18281
rect 35860 18244 35905 18272
rect 35860 18232 35866 18244
rect 36081 18241 36093 18275
rect 36127 18272 36139 18275
rect 36354 18272 36360 18284
rect 36127 18244 36360 18272
rect 36127 18241 36139 18244
rect 36081 18235 36139 18241
rect 36354 18232 36360 18244
rect 36412 18232 36418 18284
rect 28718 18204 28724 18216
rect 28307 18176 28488 18204
rect 28679 18176 28724 18204
rect 28307 18173 28319 18176
rect 28261 18167 28319 18173
rect 28718 18164 28724 18176
rect 28776 18164 28782 18216
rect 30650 18164 30656 18216
rect 30708 18164 30714 18216
rect 31110 18204 31116 18216
rect 31071 18176 31116 18204
rect 31110 18164 31116 18176
rect 31168 18164 31174 18216
rect 33594 18164 33600 18216
rect 33652 18204 33658 18216
rect 36170 18204 36176 18216
rect 33652 18176 36176 18204
rect 33652 18164 33658 18176
rect 36170 18164 36176 18176
rect 36228 18164 36234 18216
rect 38010 18204 38016 18216
rect 37971 18176 38016 18204
rect 38010 18164 38016 18176
rect 38068 18164 38074 18216
rect 18656 18108 22232 18136
rect 22296 18108 23704 18136
rect 18656 18096 18662 18108
rect 19426 18068 19432 18080
rect 18524 18040 19432 18068
rect 19426 18028 19432 18040
rect 19484 18028 19490 18080
rect 20162 18028 20168 18080
rect 20220 18068 20226 18080
rect 22296 18077 22324 18108
rect 23676 18080 23704 18108
rect 23750 18096 23756 18148
rect 23808 18136 23814 18148
rect 27890 18136 27896 18148
rect 23808 18108 27896 18136
rect 23808 18096 23814 18108
rect 27890 18096 27896 18108
rect 27948 18096 27954 18148
rect 29086 18096 29092 18148
rect 29144 18136 29150 18148
rect 35434 18136 35440 18148
rect 29144 18108 35440 18136
rect 29144 18096 29150 18108
rect 35434 18096 35440 18108
rect 35492 18096 35498 18148
rect 35986 18136 35992 18148
rect 35947 18108 35992 18136
rect 35986 18096 35992 18108
rect 36044 18136 36050 18148
rect 36630 18136 36636 18148
rect 36044 18108 36636 18136
rect 36044 18096 36050 18108
rect 36630 18096 36636 18108
rect 36688 18096 36694 18148
rect 22281 18071 22339 18077
rect 22281 18068 22293 18071
rect 20220 18040 22293 18068
rect 20220 18028 20226 18040
rect 22281 18037 22293 18040
rect 22327 18037 22339 18071
rect 22462 18068 22468 18080
rect 22423 18040 22468 18068
rect 22281 18031 22339 18037
rect 22462 18028 22468 18040
rect 22520 18028 22526 18080
rect 23109 18071 23167 18077
rect 23109 18037 23121 18071
rect 23155 18068 23167 18071
rect 23198 18068 23204 18080
rect 23155 18040 23204 18068
rect 23155 18037 23167 18040
rect 23109 18031 23167 18037
rect 23198 18028 23204 18040
rect 23256 18028 23262 18080
rect 23658 18028 23664 18080
rect 23716 18028 23722 18080
rect 29549 18071 29607 18077
rect 29549 18037 29561 18071
rect 29595 18068 29607 18071
rect 33502 18068 33508 18080
rect 29595 18040 33508 18068
rect 29595 18037 29607 18040
rect 29549 18031 29607 18037
rect 33502 18028 33508 18040
rect 33560 18028 33566 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 11422 17864 11428 17876
rect 11383 17836 11428 17864
rect 11422 17824 11428 17836
rect 11480 17824 11486 17876
rect 15102 17824 15108 17876
rect 15160 17864 15166 17876
rect 21542 17864 21548 17876
rect 15160 17836 21548 17864
rect 15160 17824 15166 17836
rect 21542 17824 21548 17836
rect 21600 17824 21606 17876
rect 24026 17864 24032 17876
rect 22848 17836 24032 17864
rect 15194 17756 15200 17808
rect 15252 17756 15258 17808
rect 17494 17756 17500 17808
rect 17552 17796 17558 17808
rect 17552 17768 19748 17796
rect 17552 17756 17558 17768
rect 5810 17728 5816 17740
rect 5771 17700 5816 17728
rect 5810 17688 5816 17700
rect 5868 17688 5874 17740
rect 9122 17688 9128 17740
rect 9180 17728 9186 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9180 17700 10057 17728
rect 9180 17688 9186 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 12710 17688 12716 17740
rect 12768 17728 12774 17740
rect 12805 17731 12863 17737
rect 12805 17728 12817 17731
rect 12768 17700 12817 17728
rect 12768 17688 12774 17700
rect 12805 17697 12817 17700
rect 12851 17697 12863 17731
rect 12805 17691 12863 17697
rect 12989 17731 13047 17737
rect 12989 17697 13001 17731
rect 13035 17728 13047 17731
rect 13998 17728 14004 17740
rect 13035 17700 14004 17728
rect 13035 17697 13047 17700
rect 12989 17691 13047 17697
rect 13998 17688 14004 17700
rect 14056 17688 14062 17740
rect 15212 17728 15240 17756
rect 15028 17700 15240 17728
rect 16761 17731 16819 17737
rect 6086 17669 6092 17672
rect 6080 17660 6092 17669
rect 6047 17632 6092 17660
rect 6080 17623 6092 17632
rect 6086 17620 6092 17623
rect 6144 17620 6150 17672
rect 10312 17663 10370 17669
rect 10312 17629 10324 17663
rect 10358 17660 10370 17663
rect 10594 17660 10600 17672
rect 10358 17632 10600 17660
rect 10358 17629 10370 17632
rect 10312 17623 10370 17629
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 13078 17620 13084 17672
rect 13136 17660 13142 17672
rect 15028 17669 15056 17700
rect 16761 17697 16773 17731
rect 16807 17728 16819 17731
rect 16850 17728 16856 17740
rect 16807 17700 16856 17728
rect 16807 17697 16819 17700
rect 16761 17691 16819 17697
rect 16850 17688 16856 17700
rect 16908 17688 16914 17740
rect 14645 17663 14703 17669
rect 14645 17660 14657 17663
rect 13136 17632 14657 17660
rect 13136 17620 13142 17632
rect 14645 17629 14657 17632
rect 14691 17629 14703 17663
rect 14645 17623 14703 17629
rect 14738 17663 14796 17669
rect 14738 17629 14750 17663
rect 14784 17629 14796 17663
rect 14738 17623 14796 17629
rect 15013 17663 15071 17669
rect 15013 17629 15025 17663
rect 15059 17629 15071 17663
rect 15013 17623 15071 17629
rect 13814 17552 13820 17604
rect 13872 17592 13878 17604
rect 14752 17592 14780 17623
rect 15102 17620 15108 17672
rect 15160 17669 15166 17672
rect 15160 17660 15168 17669
rect 19518 17660 19524 17672
rect 15160 17632 15205 17660
rect 15304 17632 19524 17660
rect 15160 17623 15168 17632
rect 15160 17620 15166 17623
rect 14918 17592 14924 17604
rect 13872 17564 14780 17592
rect 14879 17564 14924 17592
rect 13872 17552 13878 17564
rect 14918 17552 14924 17564
rect 14976 17552 14982 17604
rect 15304 17592 15332 17632
rect 19518 17620 19524 17632
rect 19576 17620 19582 17672
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17660 19671 17663
rect 19720 17660 19748 17768
rect 20162 17756 20168 17808
rect 20220 17796 20226 17808
rect 21821 17799 21879 17805
rect 21821 17796 21833 17799
rect 20220 17768 21833 17796
rect 20220 17756 20226 17768
rect 21821 17765 21833 17768
rect 21867 17765 21879 17799
rect 21821 17759 21879 17765
rect 22646 17728 22652 17740
rect 21560 17700 22652 17728
rect 21266 17660 21272 17672
rect 19659 17632 19748 17660
rect 21227 17632 21272 17660
rect 19659 17629 19671 17632
rect 19613 17623 19671 17629
rect 21266 17620 21272 17632
rect 21324 17620 21330 17672
rect 21560 17669 21588 17700
rect 22646 17688 22652 17700
rect 22704 17688 22710 17740
rect 21545 17663 21603 17669
rect 21545 17629 21557 17663
rect 21591 17629 21603 17663
rect 21545 17623 21603 17629
rect 21689 17663 21747 17669
rect 21689 17629 21701 17663
rect 21735 17660 21747 17663
rect 22094 17660 22100 17672
rect 21735 17632 22100 17660
rect 21735 17629 21747 17632
rect 21689 17623 21747 17629
rect 22094 17620 22100 17632
rect 22152 17620 22158 17672
rect 22848 17660 22876 17836
rect 24026 17824 24032 17836
rect 24084 17824 24090 17876
rect 25590 17864 25596 17876
rect 24688 17836 25596 17864
rect 22925 17799 22983 17805
rect 22925 17765 22937 17799
rect 22971 17796 22983 17799
rect 22971 17768 24256 17796
rect 22971 17765 22983 17768
rect 22925 17759 22983 17765
rect 23106 17688 23112 17740
rect 23164 17728 23170 17740
rect 24118 17728 24124 17740
rect 23164 17700 24124 17728
rect 23164 17688 23170 17700
rect 24118 17688 24124 17700
rect 24176 17688 24182 17740
rect 22925 17663 22983 17669
rect 22925 17660 22937 17663
rect 22848 17632 22937 17660
rect 22925 17629 22937 17632
rect 22971 17629 22983 17663
rect 23198 17660 23204 17672
rect 23159 17632 23204 17660
rect 22925 17623 22983 17629
rect 23198 17620 23204 17632
rect 23256 17660 23262 17672
rect 23566 17660 23572 17672
rect 23256 17632 23572 17660
rect 23256 17620 23262 17632
rect 23566 17620 23572 17632
rect 23624 17620 23630 17672
rect 23661 17663 23719 17669
rect 23661 17629 23673 17663
rect 23707 17660 23719 17663
rect 23934 17660 23940 17672
rect 23707 17632 23940 17660
rect 23707 17629 23719 17632
rect 23661 17623 23719 17629
rect 23934 17620 23940 17632
rect 23992 17620 23998 17672
rect 15028 17564 15332 17592
rect 7190 17524 7196 17536
rect 7151 17496 7196 17524
rect 7190 17484 7196 17496
rect 7248 17484 7254 17536
rect 12342 17524 12348 17536
rect 12303 17496 12348 17524
rect 12342 17484 12348 17496
rect 12400 17484 12406 17536
rect 12713 17527 12771 17533
rect 12713 17493 12725 17527
rect 12759 17524 12771 17527
rect 13078 17524 13084 17536
rect 12759 17496 13084 17524
rect 12759 17493 12771 17496
rect 12713 17487 12771 17493
rect 13078 17484 13084 17496
rect 13136 17524 13142 17536
rect 15028 17524 15056 17564
rect 15470 17552 15476 17604
rect 15528 17592 15534 17604
rect 16577 17595 16635 17601
rect 16577 17592 16589 17595
rect 15528 17564 16589 17592
rect 15528 17552 15534 17564
rect 16577 17561 16589 17564
rect 16623 17561 16635 17595
rect 16577 17555 16635 17561
rect 18046 17552 18052 17604
rect 18104 17592 18110 17604
rect 21284 17592 21312 17620
rect 18104 17564 21312 17592
rect 18104 17552 18110 17564
rect 21450 17552 21456 17604
rect 21508 17592 21514 17604
rect 22186 17592 22192 17604
rect 21508 17564 22192 17592
rect 21508 17552 21514 17564
rect 22186 17552 22192 17564
rect 22244 17552 22250 17604
rect 23750 17552 23756 17604
rect 23808 17592 23814 17604
rect 23845 17595 23903 17601
rect 23845 17592 23857 17595
rect 23808 17564 23857 17592
rect 23808 17552 23814 17564
rect 23845 17561 23857 17564
rect 23891 17561 23903 17595
rect 24228 17592 24256 17768
rect 24688 17740 24716 17836
rect 25590 17824 25596 17836
rect 25648 17824 25654 17876
rect 29086 17864 29092 17876
rect 26436 17836 29092 17864
rect 24670 17728 24676 17740
rect 24583 17700 24676 17728
rect 24670 17688 24676 17700
rect 24728 17688 24734 17740
rect 24762 17660 24768 17672
rect 24723 17632 24768 17660
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 25225 17663 25283 17669
rect 25225 17629 25237 17663
rect 25271 17629 25283 17663
rect 25225 17623 25283 17629
rect 25240 17592 25268 17623
rect 25314 17620 25320 17672
rect 25372 17660 25378 17672
rect 25372 17632 25417 17660
rect 25372 17620 25378 17632
rect 26326 17620 26332 17672
rect 26384 17660 26390 17672
rect 26436 17660 26464 17836
rect 29086 17824 29092 17836
rect 29144 17824 29150 17876
rect 30282 17864 30288 17876
rect 30243 17836 30288 17864
rect 30282 17824 30288 17836
rect 30340 17824 30346 17876
rect 31110 17824 31116 17876
rect 31168 17864 31174 17876
rect 31389 17867 31447 17873
rect 31389 17864 31401 17867
rect 31168 17836 31401 17864
rect 31168 17824 31174 17836
rect 31389 17833 31401 17836
rect 31435 17833 31447 17867
rect 33502 17864 33508 17876
rect 33463 17836 33508 17864
rect 31389 17827 31447 17833
rect 33502 17824 33508 17836
rect 33560 17824 33566 17876
rect 28718 17756 28724 17808
rect 28776 17796 28782 17808
rect 36722 17796 36728 17808
rect 28776 17768 36728 17796
rect 28776 17756 28782 17768
rect 27338 17688 27344 17740
rect 27396 17688 27402 17740
rect 30558 17688 30564 17740
rect 30616 17728 30622 17740
rect 30616 17700 31616 17728
rect 30616 17688 30622 17700
rect 26384 17632 26464 17660
rect 26384 17620 26390 17632
rect 26602 17620 26608 17672
rect 26660 17660 26666 17672
rect 27065 17663 27123 17669
rect 27065 17660 27077 17663
rect 26660 17632 27077 17660
rect 26660 17620 26666 17632
rect 27065 17629 27077 17632
rect 27111 17629 27123 17663
rect 27065 17623 27123 17629
rect 27154 17620 27160 17672
rect 27212 17660 27218 17672
rect 27356 17660 27384 17688
rect 27530 17663 27588 17669
rect 27530 17660 27542 17663
rect 27212 17632 27257 17660
rect 27356 17632 27542 17660
rect 27212 17620 27218 17632
rect 27530 17629 27542 17632
rect 27576 17660 27588 17663
rect 28074 17660 28080 17672
rect 27576 17632 28080 17660
rect 27576 17629 27588 17632
rect 27530 17623 27588 17629
rect 28074 17620 28080 17632
rect 28132 17620 28138 17672
rect 29822 17620 29828 17672
rect 29880 17669 29886 17672
rect 29880 17663 29916 17669
rect 29904 17629 29916 17663
rect 30374 17660 30380 17672
rect 30335 17632 30380 17660
rect 29880 17623 29916 17629
rect 29880 17620 29886 17623
rect 30374 17620 30380 17632
rect 30432 17620 30438 17672
rect 30837 17663 30895 17669
rect 30837 17629 30849 17663
rect 30883 17660 30895 17663
rect 30926 17660 30932 17672
rect 30883 17632 30932 17660
rect 30883 17629 30895 17632
rect 30837 17623 30895 17629
rect 30926 17620 30932 17632
rect 30984 17620 30990 17672
rect 31205 17663 31263 17669
rect 31205 17629 31217 17663
rect 31251 17660 31263 17663
rect 31251 17632 31524 17660
rect 31251 17629 31263 17632
rect 31205 17623 31263 17629
rect 24228 17564 25268 17592
rect 23845 17555 23903 17561
rect 26694 17552 26700 17604
rect 26752 17592 26758 17604
rect 27341 17595 27399 17601
rect 27341 17592 27353 17595
rect 26752 17564 27353 17592
rect 26752 17552 26758 17564
rect 27341 17561 27353 17564
rect 27387 17561 27399 17595
rect 27341 17555 27399 17561
rect 27430 17552 27436 17604
rect 27488 17592 27494 17604
rect 31018 17592 31024 17604
rect 27488 17564 27533 17592
rect 30979 17564 31024 17592
rect 27488 17552 27494 17564
rect 31018 17552 31024 17564
rect 31076 17552 31082 17604
rect 31113 17595 31171 17601
rect 31113 17561 31125 17595
rect 31159 17592 31171 17595
rect 31294 17592 31300 17604
rect 31159 17564 31300 17592
rect 31159 17561 31171 17564
rect 31113 17555 31171 17561
rect 31294 17552 31300 17564
rect 31352 17552 31358 17604
rect 13136 17496 15056 17524
rect 15289 17527 15347 17533
rect 13136 17484 13142 17496
rect 15289 17493 15301 17527
rect 15335 17524 15347 17527
rect 15654 17524 15660 17536
rect 15335 17496 15660 17524
rect 15335 17493 15347 17496
rect 15289 17487 15347 17493
rect 15654 17484 15660 17496
rect 15712 17484 15718 17536
rect 16114 17524 16120 17536
rect 16075 17496 16120 17524
rect 16114 17484 16120 17496
rect 16172 17484 16178 17536
rect 16485 17527 16543 17533
rect 16485 17493 16497 17527
rect 16531 17524 16543 17527
rect 17954 17524 17960 17536
rect 16531 17496 17960 17524
rect 16531 17493 16543 17496
rect 16485 17487 16543 17493
rect 17954 17484 17960 17496
rect 18012 17484 18018 17536
rect 19797 17527 19855 17533
rect 19797 17493 19809 17527
rect 19843 17524 19855 17527
rect 20070 17524 20076 17536
rect 19843 17496 20076 17524
rect 19843 17493 19855 17496
rect 19797 17487 19855 17493
rect 20070 17484 20076 17496
rect 20128 17484 20134 17536
rect 23106 17524 23112 17536
rect 23067 17496 23112 17524
rect 23106 17484 23112 17496
rect 23164 17484 23170 17536
rect 24029 17527 24087 17533
rect 24029 17493 24041 17527
rect 24075 17524 24087 17527
rect 24118 17524 24124 17536
rect 24075 17496 24124 17524
rect 24075 17493 24087 17496
rect 24029 17487 24087 17493
rect 24118 17484 24124 17496
rect 24176 17524 24182 17536
rect 24578 17524 24584 17536
rect 24176 17496 24584 17524
rect 24176 17484 24182 17496
rect 24578 17484 24584 17496
rect 24636 17484 24642 17536
rect 25682 17484 25688 17536
rect 25740 17524 25746 17536
rect 25777 17527 25835 17533
rect 25777 17524 25789 17527
rect 25740 17496 25789 17524
rect 25740 17484 25746 17496
rect 25777 17493 25789 17496
rect 25823 17493 25835 17527
rect 25777 17487 25835 17493
rect 27709 17527 27767 17533
rect 27709 17493 27721 17527
rect 27755 17524 27767 17527
rect 27982 17524 27988 17536
rect 27755 17496 27988 17524
rect 27755 17493 27767 17496
rect 27709 17487 27767 17493
rect 27982 17484 27988 17496
rect 28040 17484 28046 17536
rect 29730 17524 29736 17536
rect 29691 17496 29736 17524
rect 29730 17484 29736 17496
rect 29788 17484 29794 17536
rect 29914 17524 29920 17536
rect 29875 17496 29920 17524
rect 29914 17484 29920 17496
rect 29972 17484 29978 17536
rect 31496 17524 31524 17632
rect 31588 17592 31616 17700
rect 31864 17669 31892 17768
rect 36722 17756 36728 17768
rect 36780 17756 36786 17808
rect 33042 17728 33048 17740
rect 32232 17700 33048 17728
rect 32232 17669 32260 17700
rect 33042 17688 33048 17700
rect 33100 17688 33106 17740
rect 38102 17728 38108 17740
rect 38063 17700 38108 17728
rect 38102 17688 38108 17700
rect 38160 17688 38166 17740
rect 31849 17663 31907 17669
rect 31849 17629 31861 17663
rect 31895 17629 31907 17663
rect 32033 17663 32091 17669
rect 32033 17660 32045 17663
rect 31849 17623 31907 17629
rect 31956 17632 32045 17660
rect 31956 17604 31984 17632
rect 32033 17629 32045 17632
rect 32079 17629 32091 17663
rect 32033 17623 32091 17629
rect 32217 17663 32275 17669
rect 32217 17629 32229 17663
rect 32263 17629 32275 17663
rect 33134 17660 33140 17672
rect 33095 17632 33140 17660
rect 32217 17623 32275 17629
rect 31938 17592 31944 17604
rect 31588 17564 31944 17592
rect 31938 17552 31944 17564
rect 31996 17552 32002 17604
rect 32122 17592 32128 17604
rect 32083 17564 32128 17592
rect 32122 17552 32128 17564
rect 32180 17552 32186 17604
rect 32232 17524 32260 17623
rect 33134 17620 33140 17632
rect 33192 17620 33198 17672
rect 33318 17620 33324 17672
rect 33376 17660 33382 17672
rect 33505 17663 33563 17669
rect 33505 17660 33517 17663
rect 33376 17632 33517 17660
rect 33376 17620 33382 17632
rect 33505 17629 33517 17632
rect 33551 17629 33563 17663
rect 37826 17660 37832 17672
rect 37787 17632 37832 17660
rect 33505 17623 33563 17629
rect 37826 17620 37832 17632
rect 37884 17620 37890 17672
rect 31496 17496 32260 17524
rect 32401 17527 32459 17533
rect 32401 17493 32413 17527
rect 32447 17524 32459 17527
rect 33226 17524 33232 17536
rect 32447 17496 33232 17524
rect 32447 17493 32459 17496
rect 32401 17487 32459 17493
rect 33226 17484 33232 17496
rect 33284 17484 33290 17536
rect 33321 17527 33379 17533
rect 33321 17493 33333 17527
rect 33367 17524 33379 17527
rect 33686 17524 33692 17536
rect 33367 17496 33692 17524
rect 33367 17493 33379 17496
rect 33321 17487 33379 17493
rect 33686 17484 33692 17496
rect 33744 17484 33750 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 7190 17280 7196 17332
rect 7248 17320 7254 17332
rect 14829 17323 14887 17329
rect 7248 17292 14780 17320
rect 7248 17280 7254 17292
rect 7650 17212 7656 17264
rect 7708 17252 7714 17264
rect 8297 17255 8355 17261
rect 8297 17252 8309 17255
rect 7708 17224 8309 17252
rect 7708 17212 7714 17224
rect 8297 17221 8309 17224
rect 8343 17221 8355 17255
rect 8297 17215 8355 17221
rect 8389 17255 8447 17261
rect 8389 17221 8401 17255
rect 8435 17252 8447 17255
rect 10502 17252 10508 17264
rect 8435 17224 10508 17252
rect 8435 17221 8447 17224
rect 8389 17215 8447 17221
rect 10502 17212 10508 17224
rect 10560 17212 10566 17264
rect 11968 17255 12026 17261
rect 11968 17221 11980 17255
rect 12014 17252 12026 17255
rect 12342 17252 12348 17264
rect 12014 17224 12348 17252
rect 12014 17221 12026 17224
rect 11968 17215 12026 17221
rect 12342 17212 12348 17224
rect 12400 17212 12406 17264
rect 14752 17252 14780 17292
rect 14829 17289 14841 17323
rect 14875 17320 14887 17323
rect 14918 17320 14924 17332
rect 14875 17292 14924 17320
rect 14875 17289 14887 17292
rect 14829 17283 14887 17289
rect 14918 17280 14924 17292
rect 14976 17280 14982 17332
rect 15470 17320 15476 17332
rect 15431 17292 15476 17320
rect 15470 17280 15476 17292
rect 15528 17280 15534 17332
rect 19334 17280 19340 17332
rect 19392 17320 19398 17332
rect 19613 17323 19671 17329
rect 19613 17320 19625 17323
rect 19392 17292 19625 17320
rect 19392 17280 19398 17292
rect 19613 17289 19625 17292
rect 19659 17320 19671 17323
rect 23106 17320 23112 17332
rect 19659 17292 23112 17320
rect 19659 17289 19671 17292
rect 19613 17283 19671 17289
rect 23106 17280 23112 17292
rect 23164 17280 23170 17332
rect 23661 17323 23719 17329
rect 23661 17289 23673 17323
rect 23707 17320 23719 17323
rect 23842 17320 23848 17332
rect 23707 17292 23848 17320
rect 23707 17289 23719 17292
rect 23661 17283 23719 17289
rect 23842 17280 23848 17292
rect 23900 17280 23906 17332
rect 24305 17323 24363 17329
rect 24305 17289 24317 17323
rect 24351 17320 24363 17323
rect 25314 17320 25320 17332
rect 24351 17292 25320 17320
rect 24351 17289 24363 17292
rect 24305 17283 24363 17289
rect 25314 17280 25320 17292
rect 25372 17280 25378 17332
rect 26605 17323 26663 17329
rect 26605 17289 26617 17323
rect 26651 17320 26663 17323
rect 30374 17320 30380 17332
rect 26651 17292 30380 17320
rect 26651 17289 26663 17292
rect 26605 17283 26663 17289
rect 30374 17280 30380 17292
rect 30432 17280 30438 17332
rect 37734 17320 37740 17332
rect 35452 17292 37740 17320
rect 17310 17252 17316 17264
rect 14752 17224 17316 17252
rect 8018 17144 8024 17196
rect 8076 17184 8082 17196
rect 8113 17187 8171 17193
rect 8113 17184 8125 17187
rect 8076 17156 8125 17184
rect 8076 17144 8082 17156
rect 8113 17153 8125 17156
rect 8159 17153 8171 17187
rect 8113 17147 8171 17153
rect 8202 17144 8208 17196
rect 8260 17184 8266 17196
rect 14752 17193 14780 17224
rect 17310 17212 17316 17224
rect 17368 17212 17374 17264
rect 18138 17212 18144 17264
rect 18196 17252 18202 17264
rect 18478 17255 18536 17261
rect 18478 17252 18490 17255
rect 18196 17224 18490 17252
rect 18196 17212 18202 17224
rect 18478 17221 18490 17224
rect 18524 17221 18536 17255
rect 18478 17215 18536 17221
rect 22557 17255 22615 17261
rect 22557 17221 22569 17255
rect 22603 17221 22615 17255
rect 22557 17215 22615 17221
rect 22773 17255 22831 17261
rect 22773 17221 22785 17255
rect 22819 17252 22831 17255
rect 22922 17252 22928 17264
rect 22819 17224 22928 17252
rect 22819 17221 22831 17224
rect 22773 17215 22831 17221
rect 8481 17187 8539 17193
rect 8481 17184 8493 17187
rect 8260 17156 8493 17184
rect 8260 17144 8266 17156
rect 8481 17153 8493 17156
rect 8527 17153 8539 17187
rect 8481 17147 8539 17153
rect 14737 17187 14795 17193
rect 14737 17153 14749 17187
rect 14783 17153 14795 17187
rect 14737 17147 14795 17153
rect 14921 17187 14979 17193
rect 14921 17153 14933 17187
rect 14967 17184 14979 17187
rect 15194 17184 15200 17196
rect 14967 17156 15200 17184
rect 14967 17153 14979 17156
rect 14921 17147 14979 17153
rect 15194 17144 15200 17156
rect 15252 17144 15258 17196
rect 15654 17184 15660 17196
rect 15615 17156 15660 17184
rect 15654 17144 15660 17156
rect 15712 17144 15718 17196
rect 15838 17184 15844 17196
rect 15799 17156 15844 17184
rect 15838 17144 15844 17156
rect 15896 17144 15902 17196
rect 15933 17187 15991 17193
rect 15933 17153 15945 17187
rect 15979 17184 15991 17187
rect 18046 17184 18052 17196
rect 15979 17156 18052 17184
rect 15979 17153 15991 17156
rect 15933 17147 15991 17153
rect 18046 17144 18052 17156
rect 18104 17144 18110 17196
rect 18230 17184 18236 17196
rect 18191 17156 18236 17184
rect 18230 17144 18236 17156
rect 18288 17144 18294 17196
rect 22572 17184 22600 17215
rect 22922 17212 22928 17224
rect 22980 17212 22986 17264
rect 23198 17212 23204 17264
rect 23256 17252 23262 17264
rect 26237 17255 26295 17261
rect 23256 17224 24532 17252
rect 23256 17212 23262 17224
rect 23014 17184 23020 17196
rect 22572 17156 23020 17184
rect 23014 17144 23020 17156
rect 23072 17184 23078 17196
rect 24504 17193 24532 17224
rect 26237 17221 26249 17255
rect 26283 17252 26295 17255
rect 27338 17252 27344 17264
rect 26283 17224 27344 17252
rect 26283 17221 26295 17224
rect 26237 17215 26295 17221
rect 27338 17212 27344 17224
rect 27396 17212 27402 17264
rect 27706 17212 27712 17264
rect 27764 17252 27770 17264
rect 28445 17255 28503 17261
rect 27764 17224 28212 17252
rect 27764 17212 27770 17224
rect 23385 17187 23443 17193
rect 23385 17184 23397 17187
rect 23072 17156 23397 17184
rect 23072 17144 23078 17156
rect 23385 17153 23397 17156
rect 23431 17153 23443 17187
rect 23385 17147 23443 17153
rect 23569 17187 23627 17193
rect 23569 17153 23581 17187
rect 23615 17153 23627 17187
rect 23569 17147 23627 17153
rect 24489 17187 24547 17193
rect 24489 17153 24501 17187
rect 24535 17153 24547 17187
rect 24489 17147 24547 17153
rect 7834 17076 7840 17128
rect 7892 17116 7898 17128
rect 8220 17116 8248 17144
rect 11698 17116 11704 17128
rect 7892 17088 8248 17116
rect 11659 17088 11704 17116
rect 7892 17076 7898 17088
rect 11698 17076 11704 17088
rect 11756 17076 11762 17128
rect 15562 17076 15568 17128
rect 15620 17116 15626 17128
rect 17126 17116 17132 17128
rect 15620 17088 17132 17116
rect 15620 17076 15626 17088
rect 17126 17076 17132 17088
rect 17184 17076 17190 17128
rect 22830 17076 22836 17128
rect 22888 17116 22894 17128
rect 23584 17116 23612 17147
rect 24578 17144 24584 17196
rect 24636 17184 24642 17196
rect 26050 17184 26056 17196
rect 24636 17156 24681 17184
rect 26011 17156 26056 17184
rect 24636 17144 24642 17156
rect 26050 17144 26056 17156
rect 26108 17144 26114 17196
rect 26326 17184 26332 17196
rect 26287 17156 26332 17184
rect 26326 17144 26332 17156
rect 26384 17144 26390 17196
rect 26418 17144 26424 17196
rect 26476 17184 26482 17196
rect 27157 17187 27215 17193
rect 26476 17156 26521 17184
rect 26476 17144 26482 17156
rect 27157 17153 27169 17187
rect 27203 17153 27215 17187
rect 27430 17184 27436 17196
rect 27391 17156 27436 17184
rect 27157 17147 27215 17153
rect 22888 17088 23612 17116
rect 22888 17076 22894 17088
rect 24026 17076 24032 17128
rect 24084 17116 24090 17128
rect 24673 17119 24731 17125
rect 24673 17116 24685 17119
rect 24084 17088 24685 17116
rect 24084 17076 24090 17088
rect 24673 17085 24685 17088
rect 24719 17085 24731 17119
rect 24673 17079 24731 17085
rect 24762 17076 24768 17128
rect 24820 17116 24826 17128
rect 25774 17116 25780 17128
rect 24820 17088 25780 17116
rect 24820 17076 24826 17088
rect 25774 17076 25780 17088
rect 25832 17076 25838 17128
rect 13078 17048 13084 17060
rect 13039 17020 13084 17048
rect 13078 17008 13084 17020
rect 13136 17008 13142 17060
rect 13538 17008 13544 17060
rect 13596 17048 13602 17060
rect 15378 17048 15384 17060
rect 13596 17020 15384 17048
rect 13596 17008 13602 17020
rect 15378 17008 15384 17020
rect 15436 17048 15442 17060
rect 22462 17048 22468 17060
rect 15436 17020 15976 17048
rect 15436 17008 15442 17020
rect 8662 16980 8668 16992
rect 8623 16952 8668 16980
rect 8662 16940 8668 16952
rect 8720 16940 8726 16992
rect 14734 16940 14740 16992
rect 14792 16980 14798 16992
rect 15102 16980 15108 16992
rect 14792 16952 15108 16980
rect 14792 16940 14798 16952
rect 15102 16940 15108 16952
rect 15160 16940 15166 16992
rect 15948 16980 15976 17020
rect 19168 17020 22468 17048
rect 19168 16980 19196 17020
rect 22462 17008 22468 17020
rect 22520 17008 22526 17060
rect 22925 17051 22983 17057
rect 22925 17017 22937 17051
rect 22971 17048 22983 17051
rect 23934 17048 23940 17060
rect 22971 17020 23940 17048
rect 22971 17017 22983 17020
rect 22925 17011 22983 17017
rect 23934 17008 23940 17020
rect 23992 17008 23998 17060
rect 27172 17048 27200 17147
rect 27430 17144 27436 17156
rect 27488 17144 27494 17196
rect 28184 17193 28212 17224
rect 28445 17221 28457 17255
rect 28491 17252 28503 17255
rect 28718 17252 28724 17264
rect 28491 17224 28724 17252
rect 28491 17221 28503 17224
rect 28445 17215 28503 17221
rect 28718 17212 28724 17224
rect 28776 17212 28782 17264
rect 29178 17212 29184 17264
rect 29236 17252 29242 17264
rect 30101 17255 30159 17261
rect 30101 17252 30113 17255
rect 29236 17224 30113 17252
rect 29236 17212 29242 17224
rect 30101 17221 30113 17224
rect 30147 17221 30159 17255
rect 30101 17215 30159 17221
rect 30650 17212 30656 17264
rect 30708 17252 30714 17264
rect 31294 17252 31300 17264
rect 30708 17224 31300 17252
rect 30708 17212 30714 17224
rect 31294 17212 31300 17224
rect 31352 17252 31358 17264
rect 32582 17252 32588 17264
rect 31352 17224 32588 17252
rect 31352 17212 31358 17224
rect 32582 17212 32588 17224
rect 32640 17212 32646 17264
rect 35452 17261 35480 17292
rect 37734 17280 37740 17292
rect 37792 17280 37798 17332
rect 37826 17280 37832 17332
rect 37884 17280 37890 17332
rect 35437 17255 35495 17261
rect 35437 17252 35449 17255
rect 32968 17224 35449 17252
rect 27525 17187 27583 17193
rect 27525 17153 27537 17187
rect 27571 17153 27583 17187
rect 27525 17147 27583 17153
rect 28169 17187 28227 17193
rect 28169 17153 28181 17187
rect 28215 17153 28227 17187
rect 28169 17147 28227 17153
rect 28353 17187 28411 17193
rect 28353 17153 28365 17187
rect 28399 17153 28411 17187
rect 28353 17147 28411 17153
rect 28537 17187 28595 17193
rect 28537 17153 28549 17187
rect 28583 17153 28595 17187
rect 29825 17187 29883 17193
rect 29825 17184 29837 17187
rect 28537 17147 28595 17153
rect 28966 17156 29837 17184
rect 27338 17076 27344 17128
rect 27396 17116 27402 17128
rect 27540 17116 27568 17147
rect 27396 17088 27568 17116
rect 27396 17076 27402 17088
rect 24044 17020 27200 17048
rect 27540 17048 27568 17088
rect 28074 17076 28080 17128
rect 28132 17116 28138 17128
rect 28368 17116 28396 17147
rect 28132 17088 28396 17116
rect 28132 17076 28138 17088
rect 28552 17048 28580 17147
rect 28718 17076 28724 17128
rect 28776 17116 28782 17128
rect 28966 17116 28994 17156
rect 29825 17153 29837 17156
rect 29871 17153 29883 17187
rect 30006 17184 30012 17196
rect 29967 17156 30012 17184
rect 29825 17147 29883 17153
rect 30006 17144 30012 17156
rect 30064 17144 30070 17196
rect 30193 17187 30251 17193
rect 30193 17153 30205 17187
rect 30239 17184 30251 17187
rect 30834 17184 30840 17196
rect 30239 17156 30840 17184
rect 30239 17153 30251 17156
rect 30193 17147 30251 17153
rect 30834 17144 30840 17156
rect 30892 17144 30898 17196
rect 32968 17193 32996 17224
rect 35437 17221 35449 17224
rect 35483 17221 35495 17255
rect 35437 17215 35495 17221
rect 36173 17255 36231 17261
rect 36173 17221 36185 17255
rect 36219 17252 36231 17255
rect 37844 17252 37872 17280
rect 37921 17255 37979 17261
rect 37921 17252 37933 17255
rect 36219 17224 37933 17252
rect 36219 17221 36231 17224
rect 36173 17215 36231 17221
rect 37921 17221 37933 17224
rect 37967 17221 37979 17255
rect 37921 17215 37979 17221
rect 32953 17187 33011 17193
rect 32953 17153 32965 17187
rect 32999 17153 33011 17187
rect 32953 17147 33011 17153
rect 33226 17144 33232 17196
rect 33284 17184 33290 17196
rect 33413 17187 33471 17193
rect 33413 17184 33425 17187
rect 33284 17156 33425 17184
rect 33284 17144 33290 17156
rect 33413 17153 33425 17156
rect 33459 17153 33471 17187
rect 34238 17184 34244 17196
rect 33413 17147 33471 17153
rect 33704 17156 34244 17184
rect 28776 17088 28994 17116
rect 28776 17076 28782 17088
rect 31938 17076 31944 17128
rect 31996 17116 32002 17128
rect 32398 17116 32404 17128
rect 31996 17088 32404 17116
rect 31996 17076 32002 17088
rect 32398 17076 32404 17088
rect 32456 17076 32462 17128
rect 32858 17116 32864 17128
rect 32819 17088 32864 17116
rect 32858 17076 32864 17088
rect 32916 17076 32922 17128
rect 33704 17102 33732 17156
rect 34238 17144 34244 17156
rect 34296 17144 34302 17196
rect 34790 17144 34796 17196
rect 34848 17184 34854 17196
rect 35069 17187 35127 17193
rect 35069 17184 35081 17187
rect 34848 17156 35081 17184
rect 34848 17144 34854 17156
rect 35069 17153 35081 17156
rect 35115 17153 35127 17187
rect 35069 17147 35127 17153
rect 35158 17144 35164 17196
rect 35216 17184 35222 17196
rect 35342 17184 35348 17196
rect 35216 17156 35261 17184
rect 35303 17156 35348 17184
rect 35216 17144 35222 17156
rect 35342 17144 35348 17156
rect 35400 17144 35406 17196
rect 35526 17144 35532 17196
rect 35584 17193 35590 17196
rect 35584 17184 35592 17193
rect 36357 17187 36415 17193
rect 36357 17184 36369 17187
rect 35584 17156 35629 17184
rect 35728 17156 36369 17184
rect 35584 17147 35592 17156
rect 35584 17144 35590 17147
rect 27540 17020 28580 17048
rect 15948 16952 19196 16980
rect 22480 16980 22508 17008
rect 22701 16983 22759 16989
rect 22701 16980 22713 16983
rect 22480 16952 22713 16980
rect 22701 16949 22713 16952
rect 22747 16949 22759 16983
rect 22701 16943 22759 16949
rect 23106 16940 23112 16992
rect 23164 16980 23170 16992
rect 24044 16980 24072 17020
rect 31018 17008 31024 17060
rect 31076 17048 31082 17060
rect 32876 17048 32904 17076
rect 31076 17020 32904 17048
rect 31076 17008 31082 17020
rect 33318 17008 33324 17060
rect 33376 17048 33382 17060
rect 35728 17057 35756 17156
rect 36357 17153 36369 17156
rect 36403 17153 36415 17187
rect 36357 17147 36415 17153
rect 36449 17187 36507 17193
rect 36449 17153 36461 17187
rect 36495 17153 36507 17187
rect 36722 17184 36728 17196
rect 36683 17156 36728 17184
rect 36449 17147 36507 17153
rect 33781 17051 33839 17057
rect 33781 17048 33793 17051
rect 33376 17020 33793 17048
rect 33376 17008 33382 17020
rect 33781 17017 33793 17020
rect 33827 17017 33839 17051
rect 33781 17011 33839 17017
rect 35713 17051 35771 17057
rect 35713 17017 35725 17051
rect 35759 17017 35771 17051
rect 35713 17011 35771 17017
rect 27706 16980 27712 16992
rect 23164 16952 24072 16980
rect 27667 16952 27712 16980
rect 23164 16940 23170 16952
rect 27706 16940 27712 16952
rect 27764 16940 27770 16992
rect 28721 16983 28779 16989
rect 28721 16949 28733 16983
rect 28767 16980 28779 16983
rect 29270 16980 29276 16992
rect 28767 16952 29276 16980
rect 28767 16949 28779 16952
rect 28721 16943 28779 16949
rect 29270 16940 29276 16952
rect 29328 16940 29334 16992
rect 30377 16983 30435 16989
rect 30377 16949 30389 16983
rect 30423 16980 30435 16983
rect 32950 16980 32956 16992
rect 30423 16952 32956 16980
rect 30423 16949 30435 16952
rect 30377 16943 30435 16949
rect 32950 16940 32956 16952
rect 33008 16940 33014 16992
rect 35342 16940 35348 16992
rect 35400 16980 35406 16992
rect 36464 16980 36492 17147
rect 36722 17144 36728 17156
rect 36780 17144 36786 17196
rect 37734 17144 37740 17196
rect 37792 17184 37798 17196
rect 37829 17187 37887 17193
rect 37829 17184 37841 17187
rect 37792 17156 37841 17184
rect 37792 17144 37798 17156
rect 37829 17153 37841 17156
rect 37875 17153 37887 17187
rect 37829 17147 37887 17153
rect 36630 17116 36636 17128
rect 36591 17088 36636 17116
rect 36630 17076 36636 17088
rect 36688 17076 36694 17128
rect 38010 17116 38016 17128
rect 37971 17088 38016 17116
rect 38010 17076 38016 17088
rect 38068 17076 38074 17128
rect 35400 16952 36492 16980
rect 35400 16940 35406 16952
rect 37090 16940 37096 16992
rect 37148 16980 37154 16992
rect 37461 16983 37519 16989
rect 37461 16980 37473 16983
rect 37148 16952 37473 16980
rect 37148 16940 37154 16952
rect 37461 16949 37473 16952
rect 37507 16949 37519 16983
rect 37461 16943 37519 16949
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 8018 16776 8024 16788
rect 7979 16748 8024 16776
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 8202 16736 8208 16788
rect 8260 16776 8266 16788
rect 10502 16776 10508 16788
rect 8260 16748 10364 16776
rect 10463 16748 10508 16776
rect 8260 16736 8266 16748
rect 7926 16708 7932 16720
rect 6932 16680 7932 16708
rect 6932 16584 6960 16680
rect 7926 16668 7932 16680
rect 7984 16708 7990 16720
rect 10336 16708 10364 16748
rect 10502 16736 10508 16748
rect 10560 16736 10566 16788
rect 18230 16776 18236 16788
rect 16224 16748 18236 16776
rect 10870 16708 10876 16720
rect 7984 16680 9168 16708
rect 10336 16680 10876 16708
rect 7984 16668 7990 16680
rect 7834 16600 7840 16652
rect 7892 16640 7898 16652
rect 9140 16649 9168 16680
rect 10870 16668 10876 16680
rect 10928 16668 10934 16720
rect 13078 16708 13084 16720
rect 11624 16680 13084 16708
rect 9125 16643 9183 16649
rect 7892 16612 8064 16640
rect 7892 16600 7898 16612
rect 5629 16575 5687 16581
rect 5629 16541 5641 16575
rect 5675 16572 5687 16575
rect 6914 16572 6920 16584
rect 5675 16544 6920 16572
rect 5675 16541 5687 16544
rect 5629 16535 5687 16541
rect 6914 16532 6920 16544
rect 6972 16532 6978 16584
rect 8036 16581 8064 16612
rect 9125 16609 9137 16643
rect 9171 16609 9183 16643
rect 9125 16603 9183 16609
rect 8021 16575 8079 16581
rect 8021 16541 8033 16575
rect 8067 16541 8079 16575
rect 8202 16572 8208 16584
rect 8163 16544 8208 16572
rect 8021 16535 8079 16541
rect 8202 16532 8208 16544
rect 8260 16532 8266 16584
rect 8662 16532 8668 16584
rect 8720 16572 8726 16584
rect 9381 16575 9439 16581
rect 9381 16572 9393 16575
rect 8720 16544 9393 16572
rect 8720 16532 8726 16544
rect 9381 16541 9393 16544
rect 9427 16541 9439 16575
rect 9381 16535 9439 16541
rect 11517 16575 11575 16581
rect 11517 16541 11529 16575
rect 11563 16572 11575 16575
rect 11624 16572 11652 16680
rect 13078 16668 13084 16680
rect 13136 16668 13142 16720
rect 15470 16668 15476 16720
rect 15528 16708 15534 16720
rect 15657 16711 15715 16717
rect 15657 16708 15669 16711
rect 15528 16680 15669 16708
rect 15528 16668 15534 16680
rect 15657 16677 15669 16680
rect 15703 16677 15715 16711
rect 15657 16671 15715 16677
rect 11698 16600 11704 16652
rect 11756 16640 11762 16652
rect 13357 16643 13415 16649
rect 13357 16640 13369 16643
rect 11756 16612 13369 16640
rect 11756 16600 11762 16612
rect 13357 16609 13369 16612
rect 13403 16640 13415 16643
rect 14182 16640 14188 16652
rect 13403 16612 14188 16640
rect 13403 16609 13415 16612
rect 13357 16603 13415 16609
rect 14182 16600 14188 16612
rect 14240 16640 14246 16652
rect 16224 16649 16252 16748
rect 18230 16736 18236 16748
rect 18288 16736 18294 16788
rect 22002 16776 22008 16788
rect 19996 16748 22008 16776
rect 17589 16711 17647 16717
rect 17589 16677 17601 16711
rect 17635 16708 17647 16711
rect 17954 16708 17960 16720
rect 17635 16680 17960 16708
rect 17635 16677 17647 16680
rect 17589 16671 17647 16677
rect 17954 16668 17960 16680
rect 18012 16668 18018 16720
rect 19996 16649 20024 16748
rect 22002 16736 22008 16748
rect 22060 16736 22066 16788
rect 22830 16776 22836 16788
rect 22791 16748 22836 16776
rect 22830 16736 22836 16748
rect 22888 16736 22894 16788
rect 23934 16736 23940 16788
rect 23992 16776 23998 16788
rect 23992 16748 26464 16776
rect 23992 16736 23998 16748
rect 22646 16668 22652 16720
rect 22704 16708 22710 16720
rect 26326 16708 26332 16720
rect 22704 16680 26332 16708
rect 22704 16668 22710 16680
rect 26326 16668 26332 16680
rect 26384 16668 26390 16720
rect 26436 16708 26464 16748
rect 27706 16736 27712 16788
rect 27764 16776 27770 16788
rect 27764 16748 28856 16776
rect 27764 16736 27770 16748
rect 27890 16708 27896 16720
rect 26436 16680 27896 16708
rect 27890 16668 27896 16680
rect 27948 16668 27954 16720
rect 16209 16643 16267 16649
rect 16209 16640 16221 16643
rect 14240 16612 16221 16640
rect 14240 16600 14246 16612
rect 16209 16609 16221 16612
rect 16255 16609 16267 16643
rect 16209 16603 16267 16609
rect 19981 16643 20039 16649
rect 19981 16609 19993 16643
rect 20027 16609 20039 16643
rect 19981 16603 20039 16609
rect 26418 16600 26424 16652
rect 26476 16640 26482 16652
rect 27338 16640 27344 16652
rect 26476 16612 27344 16640
rect 26476 16600 26482 16612
rect 11882 16572 11888 16584
rect 11563 16544 11652 16572
rect 11843 16544 11888 16572
rect 11563 16541 11575 16544
rect 11517 16535 11575 16541
rect 11882 16532 11888 16544
rect 11940 16532 11946 16584
rect 12434 16532 12440 16584
rect 12492 16572 12498 16584
rect 12529 16575 12587 16581
rect 12529 16572 12541 16575
rect 12492 16544 12541 16572
rect 12492 16532 12498 16544
rect 12529 16541 12541 16544
rect 12575 16572 12587 16575
rect 13630 16572 13636 16584
rect 12575 16544 13636 16572
rect 12575 16541 12587 16544
rect 12529 16535 12587 16541
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 15378 16572 15384 16584
rect 15339 16544 15384 16572
rect 15378 16532 15384 16544
rect 15436 16532 15442 16584
rect 15473 16575 15531 16581
rect 15473 16541 15485 16575
rect 15519 16572 15531 16575
rect 15562 16572 15568 16584
rect 15519 16544 15568 16572
rect 15519 16541 15531 16544
rect 15473 16535 15531 16541
rect 15562 16532 15568 16544
rect 15620 16532 15626 16584
rect 16114 16532 16120 16584
rect 16172 16572 16178 16584
rect 16465 16575 16523 16581
rect 16465 16572 16477 16575
rect 16172 16544 16477 16572
rect 16172 16532 16178 16544
rect 16465 16541 16477 16544
rect 16511 16541 16523 16575
rect 16465 16535 16523 16541
rect 20070 16532 20076 16584
rect 20128 16572 20134 16584
rect 20237 16575 20295 16581
rect 20237 16572 20249 16575
rect 20128 16544 20249 16572
rect 20128 16532 20134 16544
rect 20237 16541 20249 16544
rect 20283 16541 20295 16575
rect 20237 16535 20295 16541
rect 21818 16532 21824 16584
rect 21876 16572 21882 16584
rect 22094 16572 22100 16584
rect 21876 16544 22100 16572
rect 21876 16532 21882 16544
rect 22094 16532 22100 16544
rect 22152 16532 22158 16584
rect 22462 16572 22468 16584
rect 22423 16544 22468 16572
rect 22462 16532 22468 16544
rect 22520 16532 22526 16584
rect 22922 16572 22928 16584
rect 22883 16544 22928 16572
rect 22922 16532 22928 16544
rect 22980 16532 22986 16584
rect 23106 16532 23112 16584
rect 23164 16572 23170 16584
rect 26234 16572 26240 16584
rect 23164 16544 26240 16572
rect 23164 16532 23170 16544
rect 26234 16532 26240 16544
rect 26292 16532 26298 16584
rect 26510 16572 26516 16584
rect 26471 16544 26516 16572
rect 26510 16532 26516 16544
rect 26568 16532 26574 16584
rect 26694 16572 26700 16584
rect 26655 16544 26700 16572
rect 26694 16532 26700 16544
rect 26752 16532 26758 16584
rect 26896 16581 26924 16612
rect 27338 16600 27344 16612
rect 27396 16600 27402 16652
rect 28828 16581 28856 16748
rect 28902 16736 28908 16788
rect 28960 16776 28966 16788
rect 32214 16776 32220 16788
rect 28960 16748 32220 16776
rect 28960 16736 28966 16748
rect 32214 16736 32220 16748
rect 32272 16736 32278 16788
rect 32493 16779 32551 16785
rect 32493 16745 32505 16779
rect 32539 16776 32551 16779
rect 33134 16776 33140 16788
rect 32539 16748 33140 16776
rect 32539 16745 32551 16748
rect 32493 16739 32551 16745
rect 33134 16736 33140 16748
rect 33192 16736 33198 16788
rect 37734 16736 37740 16788
rect 37792 16776 37798 16788
rect 38197 16779 38255 16785
rect 38197 16776 38209 16779
rect 37792 16748 38209 16776
rect 37792 16736 37798 16748
rect 38197 16745 38209 16748
rect 38243 16745 38255 16779
rect 38197 16739 38255 16745
rect 29086 16600 29092 16652
rect 29144 16640 29150 16652
rect 29454 16640 29460 16652
rect 29144 16612 29189 16640
rect 29288 16612 29460 16640
rect 29144 16600 29150 16612
rect 26881 16575 26939 16581
rect 26881 16541 26893 16575
rect 26927 16541 26939 16575
rect 26881 16535 26939 16541
rect 28813 16575 28871 16581
rect 28813 16541 28825 16575
rect 28859 16541 28871 16575
rect 28813 16535 28871 16541
rect 28902 16532 28908 16584
rect 28960 16572 28966 16584
rect 29178 16572 29184 16584
rect 28960 16544 29005 16572
rect 29139 16544 29184 16572
rect 28960 16532 28966 16544
rect 29178 16532 29184 16544
rect 29236 16572 29242 16584
rect 29288 16572 29316 16612
rect 29454 16600 29460 16612
rect 29512 16600 29518 16652
rect 31570 16640 31576 16652
rect 31036 16612 31576 16640
rect 31036 16581 31064 16612
rect 31570 16600 31576 16612
rect 31628 16600 31634 16652
rect 33410 16600 33416 16652
rect 33468 16640 33474 16652
rect 33597 16643 33655 16649
rect 33597 16640 33609 16643
rect 33468 16612 33609 16640
rect 33468 16600 33474 16612
rect 33597 16609 33609 16612
rect 33643 16609 33655 16643
rect 33597 16603 33655 16609
rect 34057 16643 34115 16649
rect 34057 16609 34069 16643
rect 34103 16640 34115 16643
rect 34698 16640 34704 16652
rect 34103 16612 34704 16640
rect 34103 16609 34115 16612
rect 34057 16603 34115 16609
rect 34698 16600 34704 16612
rect 34756 16600 34762 16652
rect 35434 16640 35440 16652
rect 35360 16612 35440 16640
rect 29236 16544 29316 16572
rect 31021 16575 31079 16581
rect 29236 16532 29242 16544
rect 31021 16541 31033 16575
rect 31067 16541 31079 16575
rect 31021 16535 31079 16541
rect 31113 16575 31171 16581
rect 31113 16541 31125 16575
rect 31159 16541 31171 16575
rect 31294 16572 31300 16584
rect 31255 16544 31300 16572
rect 31113 16535 31171 16541
rect 5896 16507 5954 16513
rect 5896 16473 5908 16507
rect 5942 16504 5954 16507
rect 6546 16504 6552 16516
rect 5942 16476 6552 16504
rect 5942 16473 5954 16476
rect 5896 16467 5954 16473
rect 6546 16464 6552 16476
rect 6604 16464 6610 16516
rect 10686 16464 10692 16516
rect 10744 16504 10750 16516
rect 11701 16507 11759 16513
rect 11701 16504 11713 16507
rect 10744 16476 11713 16504
rect 10744 16464 10750 16476
rect 11701 16473 11713 16476
rect 11747 16473 11759 16507
rect 11701 16467 11759 16473
rect 11793 16507 11851 16513
rect 11793 16473 11805 16507
rect 11839 16504 11851 16507
rect 13538 16504 13544 16516
rect 11839 16476 13544 16504
rect 11839 16473 11851 16476
rect 11793 16467 11851 16473
rect 13538 16464 13544 16476
rect 13596 16464 13602 16516
rect 17954 16464 17960 16516
rect 18012 16504 18018 16516
rect 26050 16504 26056 16516
rect 18012 16476 26056 16504
rect 18012 16464 18018 16476
rect 26050 16464 26056 16476
rect 26108 16464 26114 16516
rect 26786 16504 26792 16516
rect 26747 16476 26792 16504
rect 26786 16464 26792 16476
rect 26844 16464 26850 16516
rect 30926 16464 30932 16516
rect 30984 16504 30990 16516
rect 31128 16504 31156 16535
rect 31294 16532 31300 16544
rect 31352 16532 31358 16584
rect 31386 16532 31392 16584
rect 31444 16572 31450 16584
rect 31846 16572 31852 16584
rect 31444 16544 31489 16572
rect 31807 16544 31852 16572
rect 31444 16532 31450 16544
rect 31846 16532 31852 16544
rect 31904 16532 31910 16584
rect 31942 16575 32000 16581
rect 31942 16541 31954 16575
rect 31988 16541 32000 16575
rect 31942 16535 32000 16541
rect 31662 16504 31668 16516
rect 30984 16476 31668 16504
rect 30984 16464 30990 16476
rect 31662 16464 31668 16476
rect 31720 16464 31726 16516
rect 7006 16436 7012 16448
rect 6967 16408 7012 16436
rect 7006 16396 7012 16408
rect 7064 16396 7070 16448
rect 12066 16436 12072 16448
rect 12027 16408 12072 16436
rect 12066 16396 12072 16408
rect 12124 16396 12130 16448
rect 21361 16439 21419 16445
rect 21361 16405 21373 16439
rect 21407 16436 21419 16439
rect 22922 16436 22928 16448
rect 21407 16408 22928 16436
rect 21407 16405 21419 16408
rect 21361 16399 21419 16405
rect 22922 16396 22928 16408
rect 22980 16396 22986 16448
rect 27065 16439 27123 16445
rect 27065 16405 27077 16439
rect 27111 16436 27123 16439
rect 27614 16436 27620 16448
rect 27111 16408 27620 16436
rect 27111 16405 27123 16408
rect 27065 16399 27123 16405
rect 27614 16396 27620 16408
rect 27672 16396 27678 16448
rect 27798 16396 27804 16448
rect 27856 16436 27862 16448
rect 28629 16439 28687 16445
rect 28629 16436 28641 16439
rect 27856 16408 28641 16436
rect 27856 16396 27862 16408
rect 28629 16405 28641 16408
rect 28675 16405 28687 16439
rect 28629 16399 28687 16405
rect 28902 16396 28908 16448
rect 28960 16436 28966 16448
rect 30650 16436 30656 16448
rect 28960 16408 30656 16436
rect 28960 16396 28966 16408
rect 30650 16396 30656 16408
rect 30708 16396 30714 16448
rect 30834 16436 30840 16448
rect 30795 16408 30840 16436
rect 30834 16396 30840 16408
rect 30892 16396 30898 16448
rect 31956 16436 31984 16535
rect 32214 16532 32220 16584
rect 32272 16572 32278 16584
rect 32398 16581 32404 16584
rect 32355 16575 32404 16581
rect 32272 16544 32317 16572
rect 32272 16532 32278 16544
rect 32355 16541 32367 16575
rect 32401 16541 32404 16575
rect 32355 16535 32404 16541
rect 32398 16532 32404 16535
rect 32456 16532 32462 16584
rect 33686 16572 33692 16584
rect 33647 16544 33692 16572
rect 33686 16532 33692 16544
rect 33744 16532 33750 16584
rect 34790 16532 34796 16584
rect 34848 16572 34854 16584
rect 35066 16572 35072 16584
rect 34848 16544 35072 16572
rect 34848 16532 34854 16544
rect 35066 16532 35072 16544
rect 35124 16532 35130 16584
rect 35158 16532 35164 16584
rect 35216 16572 35222 16584
rect 35360 16581 35388 16612
rect 35434 16600 35440 16612
rect 35492 16600 35498 16652
rect 36814 16640 36820 16652
rect 36775 16612 36820 16640
rect 36814 16600 36820 16612
rect 36872 16600 36878 16652
rect 35345 16575 35403 16581
rect 35216 16544 35261 16572
rect 35216 16532 35222 16544
rect 35345 16541 35357 16575
rect 35391 16541 35403 16575
rect 35345 16535 35403 16541
rect 35526 16532 35532 16584
rect 35584 16581 35590 16584
rect 37090 16581 37096 16584
rect 35584 16572 35592 16581
rect 37084 16572 37096 16581
rect 35584 16544 35629 16572
rect 37051 16544 37096 16572
rect 35584 16535 35592 16544
rect 37084 16535 37096 16544
rect 35584 16532 35590 16535
rect 37090 16532 37096 16535
rect 37148 16532 37154 16584
rect 32125 16507 32183 16513
rect 32125 16473 32137 16507
rect 32171 16504 32183 16507
rect 32858 16504 32864 16516
rect 32171 16476 32864 16504
rect 32171 16473 32183 16476
rect 32125 16467 32183 16473
rect 32858 16464 32864 16476
rect 32916 16464 32922 16516
rect 35437 16507 35495 16513
rect 35437 16473 35449 16507
rect 35483 16504 35495 16507
rect 37826 16504 37832 16516
rect 35483 16476 37832 16504
rect 35483 16473 35495 16476
rect 35437 16467 35495 16473
rect 35452 16436 35480 16467
rect 37826 16464 37832 16476
rect 37884 16464 37890 16516
rect 35710 16436 35716 16448
rect 31956 16408 35480 16436
rect 35671 16408 35716 16436
rect 35710 16396 35716 16408
rect 35768 16396 35774 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 6546 16232 6552 16244
rect 6507 16204 6552 16232
rect 6546 16192 6552 16204
rect 6604 16192 6610 16244
rect 7929 16235 7987 16241
rect 7929 16201 7941 16235
rect 7975 16232 7987 16235
rect 8386 16232 8392 16244
rect 7975 16204 8392 16232
rect 7975 16201 7987 16204
rect 7929 16195 7987 16201
rect 8386 16192 8392 16204
rect 8444 16192 8450 16244
rect 13538 16232 13544 16244
rect 8772 16204 13400 16232
rect 13499 16204 13544 16232
rect 6917 16167 6975 16173
rect 6917 16133 6929 16167
rect 6963 16164 6975 16167
rect 7006 16164 7012 16176
rect 6963 16136 7012 16164
rect 6963 16133 6975 16136
rect 6917 16127 6975 16133
rect 7006 16124 7012 16136
rect 7064 16164 7070 16176
rect 8772 16164 8800 16204
rect 7064 16136 8800 16164
rect 7064 16124 7070 16136
rect 12066 16124 12072 16176
rect 12124 16164 12130 16176
rect 12406 16167 12464 16173
rect 12406 16164 12418 16167
rect 12124 16136 12418 16164
rect 12124 16124 12130 16136
rect 12406 16133 12418 16136
rect 12452 16133 12464 16167
rect 13372 16164 13400 16204
rect 13538 16192 13544 16204
rect 13596 16192 13602 16244
rect 17218 16232 17224 16244
rect 13648 16204 17224 16232
rect 13648 16164 13676 16204
rect 17218 16192 17224 16204
rect 17276 16192 17282 16244
rect 18877 16235 18935 16241
rect 18877 16201 18889 16235
rect 18923 16201 18935 16235
rect 25314 16232 25320 16244
rect 25227 16204 25320 16232
rect 18877 16195 18935 16201
rect 13372 16136 13676 16164
rect 12406 16127 12464 16133
rect 15746 16124 15752 16176
rect 15804 16164 15810 16176
rect 15841 16167 15899 16173
rect 15841 16164 15853 16167
rect 15804 16136 15853 16164
rect 15804 16124 15810 16136
rect 15841 16133 15853 16136
rect 15887 16133 15899 16167
rect 18892 16164 18920 16195
rect 25314 16192 25320 16204
rect 25372 16232 25378 16244
rect 30469 16235 30527 16241
rect 25372 16204 30420 16232
rect 25372 16192 25378 16204
rect 21634 16164 21640 16176
rect 15841 16127 15899 16133
rect 17604 16136 18920 16164
rect 19076 16136 21640 16164
rect 17604 16108 17632 16136
rect 7926 16099 7984 16105
rect 7926 16096 7938 16099
rect 7024 16068 7938 16096
rect 7024 16037 7052 16068
rect 7926 16065 7938 16068
rect 7972 16096 7984 16099
rect 8110 16096 8116 16108
rect 7972 16068 8116 16096
rect 7972 16065 7984 16068
rect 7926 16059 7984 16065
rect 8110 16056 8116 16068
rect 8168 16056 8174 16108
rect 14182 16096 14188 16108
rect 14143 16068 14188 16096
rect 14182 16056 14188 16068
rect 14240 16056 14246 16108
rect 17586 16096 17592 16108
rect 17499 16068 17592 16096
rect 17586 16056 17592 16068
rect 17644 16056 17650 16108
rect 17770 16096 17776 16108
rect 17731 16068 17776 16096
rect 17770 16056 17776 16068
rect 17828 16056 17834 16108
rect 17862 16056 17868 16108
rect 17920 16096 17926 16108
rect 19076 16105 19104 16136
rect 21634 16124 21640 16136
rect 21692 16124 21698 16176
rect 22462 16124 22468 16176
rect 22520 16164 22526 16176
rect 23014 16173 23020 16176
rect 22741 16167 22799 16173
rect 22741 16164 22753 16167
rect 22520 16136 22753 16164
rect 22520 16124 22526 16136
rect 22741 16133 22753 16136
rect 22787 16133 22799 16167
rect 22741 16127 22799 16133
rect 22957 16167 23020 16173
rect 22957 16133 22969 16167
rect 23003 16133 23020 16167
rect 22957 16127 23020 16133
rect 23014 16124 23020 16127
rect 23072 16124 23078 16176
rect 29822 16164 29828 16176
rect 27448 16136 29828 16164
rect 19061 16099 19119 16105
rect 17920 16068 17965 16096
rect 17920 16056 17926 16068
rect 19061 16065 19073 16099
rect 19107 16065 19119 16099
rect 19061 16059 19119 16065
rect 19245 16099 19303 16105
rect 19245 16065 19257 16099
rect 19291 16065 19303 16099
rect 19245 16059 19303 16065
rect 19613 16099 19671 16105
rect 19613 16065 19625 16099
rect 19659 16096 19671 16099
rect 20530 16096 20536 16108
rect 19659 16068 20536 16096
rect 19659 16065 19671 16068
rect 19613 16059 19671 16065
rect 7009 16031 7067 16037
rect 7009 15997 7021 16031
rect 7055 15997 7067 16031
rect 7009 15991 7067 15997
rect 7098 15988 7104 16040
rect 7156 16028 7162 16040
rect 7193 16031 7251 16037
rect 7193 16028 7205 16031
rect 7156 16000 7205 16028
rect 7156 15988 7162 16000
rect 7193 15997 7205 16000
rect 7239 15997 7251 16031
rect 8386 16028 8392 16040
rect 8347 16000 8392 16028
rect 7193 15991 7251 15997
rect 7208 15960 7236 15991
rect 8386 15988 8392 16000
rect 8444 15988 8450 16040
rect 12158 16028 12164 16040
rect 12119 16000 12164 16028
rect 12158 15988 12164 16000
rect 12216 15988 12222 16040
rect 14458 16028 14464 16040
rect 14419 16000 14464 16028
rect 14458 15988 14464 16000
rect 14516 15988 14522 16040
rect 17880 16028 17908 16056
rect 19260 16028 19288 16059
rect 20530 16056 20536 16068
rect 20588 16056 20594 16108
rect 22554 16056 22560 16108
rect 22612 16096 22618 16108
rect 25133 16099 25191 16105
rect 25133 16096 25145 16099
rect 22612 16068 25145 16096
rect 22612 16056 22618 16068
rect 25133 16065 25145 16068
rect 25179 16096 25191 16099
rect 26510 16096 26516 16108
rect 25179 16068 26516 16096
rect 25179 16065 25191 16068
rect 25133 16059 25191 16065
rect 26510 16056 26516 16068
rect 26568 16056 26574 16108
rect 27154 16056 27160 16108
rect 27212 16096 27218 16108
rect 27448 16105 27476 16136
rect 27433 16099 27491 16105
rect 27433 16096 27445 16099
rect 27212 16068 27445 16096
rect 27212 16056 27218 16068
rect 27433 16065 27445 16068
rect 27479 16065 27491 16099
rect 27433 16059 27491 16065
rect 27614 16056 27620 16108
rect 27672 16096 27678 16108
rect 27745 16099 27803 16105
rect 27672 16068 27717 16096
rect 27672 16056 27678 16068
rect 27745 16065 27757 16099
rect 27791 16096 27803 16099
rect 27890 16096 27896 16108
rect 27791 16068 27896 16096
rect 27791 16065 27803 16068
rect 27745 16059 27803 16065
rect 27890 16056 27896 16068
rect 27948 16056 27954 16108
rect 29196 16105 29224 16136
rect 29822 16124 29828 16136
rect 29880 16124 29886 16176
rect 29181 16099 29239 16105
rect 29181 16065 29193 16099
rect 29227 16065 29239 16099
rect 29181 16059 29239 16065
rect 29270 16056 29276 16108
rect 29328 16096 29334 16108
rect 29454 16096 29460 16108
rect 29328 16068 29373 16096
rect 29415 16068 29460 16096
rect 29328 16056 29334 16068
rect 29454 16056 29460 16068
rect 29512 16056 29518 16108
rect 17880 16000 19288 16028
rect 25409 16031 25467 16037
rect 25409 15997 25421 16031
rect 25455 16028 25467 16031
rect 25774 16028 25780 16040
rect 25455 16000 25780 16028
rect 25455 15997 25467 16000
rect 25409 15991 25467 15997
rect 25774 15988 25780 16000
rect 25832 16028 25838 16040
rect 26050 16028 26056 16040
rect 25832 16000 26056 16028
rect 25832 15988 25838 16000
rect 26050 15988 26056 16000
rect 26108 15988 26114 16040
rect 27522 15988 27528 16040
rect 27580 16037 27586 16040
rect 27580 16028 27587 16037
rect 27580 16000 27625 16028
rect 27580 15991 27587 16000
rect 27580 15988 27586 15991
rect 28994 15988 29000 16040
rect 29052 16028 29058 16040
rect 29365 16031 29423 16037
rect 29365 16028 29377 16031
rect 29052 16000 29377 16028
rect 29052 15988 29058 16000
rect 29365 15997 29377 16000
rect 29411 15997 29423 16031
rect 30392 16028 30420 16204
rect 30469 16201 30481 16235
rect 30515 16232 30527 16235
rect 31386 16232 31392 16244
rect 30515 16204 31392 16232
rect 30515 16201 30527 16204
rect 30469 16195 30527 16201
rect 31386 16192 31392 16204
rect 31444 16192 31450 16244
rect 32214 16192 32220 16244
rect 32272 16232 32278 16244
rect 35526 16232 35532 16244
rect 32272 16204 35532 16232
rect 32272 16192 32278 16204
rect 35526 16192 35532 16204
rect 35584 16232 35590 16244
rect 37826 16232 37832 16244
rect 35584 16204 36124 16232
rect 37787 16204 37832 16232
rect 35584 16192 35590 16204
rect 30558 16124 30564 16176
rect 30616 16164 30622 16176
rect 31021 16167 31079 16173
rect 31021 16164 31033 16167
rect 30616 16136 31033 16164
rect 30616 16124 30622 16136
rect 31021 16133 31033 16136
rect 31067 16133 31079 16167
rect 31021 16127 31079 16133
rect 31113 16167 31171 16173
rect 31113 16133 31125 16167
rect 31159 16164 31171 16167
rect 31478 16164 31484 16176
rect 31159 16136 31484 16164
rect 31159 16133 31171 16136
rect 31113 16127 31171 16133
rect 31478 16124 31484 16136
rect 31536 16124 31542 16176
rect 31938 16124 31944 16176
rect 31996 16164 32002 16176
rect 32582 16164 32588 16176
rect 31996 16136 32444 16164
rect 32543 16136 32588 16164
rect 31996 16124 32002 16136
rect 30466 16056 30472 16108
rect 30524 16096 30530 16108
rect 30653 16099 30711 16105
rect 30653 16096 30665 16099
rect 30524 16068 30665 16096
rect 30524 16056 30530 16068
rect 30653 16065 30665 16068
rect 30699 16065 30711 16099
rect 30653 16059 30711 16065
rect 30746 16100 30804 16106
rect 30746 16066 30758 16100
rect 30792 16097 30804 16100
rect 30792 16096 30880 16097
rect 31202 16096 31208 16108
rect 30792 16069 31208 16096
rect 30792 16066 30804 16069
rect 30852 16068 31208 16069
rect 30746 16060 30804 16066
rect 31202 16056 31208 16068
rect 31260 16056 31266 16108
rect 32309 16099 32367 16105
rect 32309 16065 32321 16099
rect 32355 16065 32367 16099
rect 32416 16096 32444 16136
rect 32582 16124 32588 16136
rect 32640 16124 32646 16176
rect 32950 16124 32956 16176
rect 33008 16164 33014 16176
rect 33008 16136 35848 16164
rect 33008 16124 33014 16136
rect 32493 16099 32551 16105
rect 32493 16096 32505 16099
rect 32416 16068 32505 16096
rect 32309 16059 32367 16065
rect 32493 16065 32505 16068
rect 32539 16065 32551 16099
rect 32674 16096 32680 16108
rect 32635 16068 32680 16096
rect 32493 16059 32551 16065
rect 32324 16028 32352 16059
rect 32674 16056 32680 16068
rect 32732 16056 32738 16108
rect 35710 16096 35716 16108
rect 35671 16068 35716 16096
rect 35710 16056 35716 16068
rect 35768 16056 35774 16108
rect 35820 16105 35848 16136
rect 36096 16105 36124 16204
rect 37826 16192 37832 16204
rect 37884 16192 37890 16244
rect 35805 16099 35863 16105
rect 35805 16065 35817 16099
rect 35851 16065 35863 16099
rect 35805 16059 35863 16065
rect 36081 16099 36139 16105
rect 36081 16065 36093 16099
rect 36127 16065 36139 16099
rect 36081 16059 36139 16065
rect 30392 16000 32352 16028
rect 35529 16031 35587 16037
rect 29365 15991 29423 15997
rect 35529 15997 35541 16031
rect 35575 16028 35587 16031
rect 37921 16031 37979 16037
rect 37921 16028 37933 16031
rect 35575 16000 37933 16028
rect 35575 15997 35587 16000
rect 35529 15991 35587 15997
rect 37844 15972 37872 16000
rect 37921 15997 37933 16000
rect 37967 15997 37979 16031
rect 37921 15991 37979 15997
rect 38010 15988 38016 16040
rect 38068 16028 38074 16040
rect 38068 16000 38113 16028
rect 38068 15988 38074 16000
rect 23109 15963 23167 15969
rect 7208 15932 8340 15960
rect 8312 15904 8340 15932
rect 23109 15929 23121 15963
rect 23155 15960 23167 15963
rect 24946 15960 24952 15972
rect 23155 15932 24952 15960
rect 23155 15929 23167 15932
rect 23109 15923 23167 15929
rect 24946 15920 24952 15932
rect 25004 15920 25010 15972
rect 26970 15920 26976 15972
rect 27028 15960 27034 15972
rect 30466 15960 30472 15972
rect 27028 15932 30472 15960
rect 27028 15920 27034 15932
rect 30466 15920 30472 15932
rect 30524 15920 30530 15972
rect 31294 15920 31300 15972
rect 31352 15960 31358 15972
rect 32861 15963 32919 15969
rect 32861 15960 32873 15963
rect 31352 15932 32873 15960
rect 31352 15920 31358 15932
rect 32861 15929 32873 15932
rect 32907 15929 32919 15963
rect 32861 15923 32919 15929
rect 35989 15963 36047 15969
rect 35989 15929 36001 15963
rect 36035 15960 36047 15963
rect 36630 15960 36636 15972
rect 36035 15932 36636 15960
rect 36035 15929 36047 15932
rect 35989 15923 36047 15929
rect 36630 15920 36636 15932
rect 36688 15920 36694 15972
rect 37826 15920 37832 15972
rect 37884 15920 37890 15972
rect 7742 15892 7748 15904
rect 7703 15864 7748 15892
rect 7742 15852 7748 15864
rect 7800 15852 7806 15904
rect 8294 15892 8300 15904
rect 8255 15864 8300 15892
rect 8294 15852 8300 15864
rect 8352 15852 8358 15904
rect 17405 15895 17463 15901
rect 17405 15861 17417 15895
rect 17451 15892 17463 15895
rect 17494 15892 17500 15904
rect 17451 15864 17500 15892
rect 17451 15861 17463 15864
rect 17405 15855 17463 15861
rect 17494 15852 17500 15864
rect 17552 15852 17558 15904
rect 22922 15892 22928 15904
rect 22883 15864 22928 15892
rect 22922 15852 22928 15864
rect 22980 15852 22986 15904
rect 24857 15895 24915 15901
rect 24857 15861 24869 15895
rect 24903 15892 24915 15895
rect 25222 15892 25228 15904
rect 24903 15864 25228 15892
rect 24903 15861 24915 15864
rect 24857 15855 24915 15861
rect 25222 15852 25228 15864
rect 25280 15852 25286 15904
rect 27249 15895 27307 15901
rect 27249 15861 27261 15895
rect 27295 15892 27307 15895
rect 27338 15892 27344 15904
rect 27295 15864 27344 15892
rect 27295 15861 27307 15864
rect 27249 15855 27307 15861
rect 27338 15852 27344 15864
rect 27396 15852 27402 15904
rect 28997 15895 29055 15901
rect 28997 15861 29009 15895
rect 29043 15892 29055 15895
rect 29270 15892 29276 15904
rect 29043 15864 29276 15892
rect 29043 15861 29055 15864
rect 28997 15855 29055 15861
rect 29270 15852 29276 15864
rect 29328 15852 29334 15904
rect 30006 15852 30012 15904
rect 30064 15892 30070 15904
rect 32674 15892 32680 15904
rect 30064 15864 32680 15892
rect 30064 15852 30070 15864
rect 32674 15852 32680 15864
rect 32732 15852 32738 15904
rect 37182 15852 37188 15904
rect 37240 15892 37246 15904
rect 37461 15895 37519 15901
rect 37461 15892 37473 15895
rect 37240 15864 37473 15892
rect 37240 15852 37246 15864
rect 37461 15861 37473 15864
rect 37507 15861 37519 15895
rect 37461 15855 37519 15861
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 6914 15688 6920 15700
rect 6748 15660 6920 15688
rect 6748 15561 6776 15660
rect 6914 15648 6920 15660
rect 6972 15648 6978 15700
rect 8113 15691 8171 15697
rect 8113 15657 8125 15691
rect 8159 15688 8171 15691
rect 8386 15688 8392 15700
rect 8159 15660 8392 15688
rect 8159 15657 8171 15660
rect 8113 15651 8171 15657
rect 8386 15648 8392 15660
rect 8444 15688 8450 15700
rect 17770 15688 17776 15700
rect 8444 15660 17776 15688
rect 8444 15648 8450 15660
rect 17770 15648 17776 15660
rect 17828 15648 17834 15700
rect 24946 15688 24952 15700
rect 24907 15660 24952 15688
rect 24946 15648 24952 15660
rect 25004 15648 25010 15700
rect 26786 15688 26792 15700
rect 25700 15660 26792 15688
rect 11146 15620 11152 15632
rect 11059 15592 11152 15620
rect 11146 15580 11152 15592
rect 11204 15620 11210 15632
rect 17862 15620 17868 15632
rect 11204 15592 15792 15620
rect 11204 15580 11210 15592
rect 6733 15555 6791 15561
rect 6733 15521 6745 15555
rect 6779 15521 6791 15555
rect 6733 15515 6791 15521
rect 7000 15487 7058 15493
rect 7000 15453 7012 15487
rect 7046 15484 7058 15487
rect 7742 15484 7748 15496
rect 7046 15456 7748 15484
rect 7046 15453 7058 15456
rect 7000 15447 7058 15453
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 9769 15487 9827 15493
rect 9769 15453 9781 15487
rect 9815 15484 9827 15487
rect 12158 15484 12164 15496
rect 9815 15456 12164 15484
rect 9815 15453 9827 15456
rect 9769 15447 9827 15453
rect 12158 15444 12164 15456
rect 12216 15444 12222 15496
rect 15764 15493 15792 15592
rect 16040 15592 17868 15620
rect 16040 15496 16068 15592
rect 17862 15580 17868 15592
rect 17920 15620 17926 15632
rect 20162 15620 20168 15632
rect 17920 15592 18460 15620
rect 20123 15592 20168 15620
rect 17920 15580 17926 15592
rect 17770 15512 17776 15564
rect 17828 15552 17834 15564
rect 18432 15561 18460 15592
rect 20162 15580 20168 15592
rect 20220 15580 20226 15632
rect 25700 15620 25728 15660
rect 26786 15648 26792 15660
rect 26844 15648 26850 15700
rect 27065 15691 27123 15697
rect 27065 15657 27077 15691
rect 27111 15688 27123 15691
rect 27890 15688 27896 15700
rect 27111 15660 27896 15688
rect 27111 15657 27123 15660
rect 27065 15651 27123 15657
rect 27890 15648 27896 15660
rect 27948 15648 27954 15700
rect 29454 15648 29460 15700
rect 29512 15688 29518 15700
rect 29825 15691 29883 15697
rect 29825 15688 29837 15691
rect 29512 15660 29837 15688
rect 29512 15648 29518 15660
rect 29825 15657 29837 15660
rect 29871 15657 29883 15691
rect 31110 15688 31116 15700
rect 29825 15651 29883 15657
rect 29932 15660 31116 15688
rect 25866 15620 25872 15632
rect 21928 15592 25728 15620
rect 25827 15592 25872 15620
rect 18417 15555 18475 15561
rect 17828 15524 18184 15552
rect 17828 15512 17834 15524
rect 15381 15487 15439 15493
rect 15381 15453 15393 15487
rect 15427 15453 15439 15487
rect 15381 15447 15439 15453
rect 15749 15487 15807 15493
rect 15749 15453 15761 15487
rect 15795 15453 15807 15487
rect 16022 15484 16028 15496
rect 15983 15456 16028 15484
rect 15749 15447 15807 15453
rect 10042 15425 10048 15428
rect 10036 15379 10048 15425
rect 10100 15416 10106 15428
rect 15396 15416 15424 15447
rect 16022 15444 16028 15456
rect 16080 15444 16086 15496
rect 17586 15484 17592 15496
rect 17547 15456 17592 15484
rect 17586 15444 17592 15456
rect 17644 15444 17650 15496
rect 18156 15493 18184 15524
rect 18417 15521 18429 15555
rect 18463 15521 18475 15555
rect 18417 15515 18475 15521
rect 19797 15555 19855 15561
rect 19797 15521 19809 15555
rect 19843 15552 19855 15555
rect 20254 15552 20260 15564
rect 19843 15524 20260 15552
rect 19843 15521 19855 15524
rect 19797 15515 19855 15521
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 21085 15555 21143 15561
rect 21085 15521 21097 15555
rect 21131 15521 21143 15555
rect 21085 15515 21143 15521
rect 18141 15487 18199 15493
rect 18141 15453 18153 15487
rect 18187 15453 18199 15487
rect 18141 15447 18199 15453
rect 17604 15416 17632 15444
rect 10100 15388 10136 15416
rect 15396 15388 17632 15416
rect 10042 15376 10048 15379
rect 10100 15376 10106 15388
rect 17770 15376 17776 15428
rect 17828 15416 17834 15428
rect 21100 15416 21128 15515
rect 21269 15487 21327 15493
rect 21269 15453 21281 15487
rect 21315 15453 21327 15487
rect 21269 15447 21327 15453
rect 17828 15388 21128 15416
rect 21284 15416 21312 15447
rect 21450 15444 21456 15496
rect 21508 15484 21514 15496
rect 21928 15493 21956 15592
rect 25866 15580 25872 15592
rect 25924 15580 25930 15632
rect 26050 15580 26056 15632
rect 26108 15620 26114 15632
rect 29932 15620 29960 15660
rect 31110 15648 31116 15660
rect 31168 15648 31174 15700
rect 34514 15688 34520 15700
rect 33060 15660 34520 15688
rect 33060 15620 33088 15660
rect 34514 15648 34520 15660
rect 34572 15648 34578 15700
rect 36354 15688 36360 15700
rect 36315 15660 36360 15688
rect 36354 15648 36360 15660
rect 36412 15648 36418 15700
rect 26108 15592 29960 15620
rect 30024 15592 33088 15620
rect 26108 15580 26114 15592
rect 22830 15512 22836 15564
rect 22888 15552 22894 15564
rect 22888 15524 23336 15552
rect 22888 15512 22894 15524
rect 21545 15487 21603 15493
rect 21545 15484 21557 15487
rect 21508 15456 21557 15484
rect 21508 15444 21514 15456
rect 21545 15453 21557 15456
rect 21591 15453 21603 15487
rect 21545 15447 21603 15453
rect 21913 15487 21971 15493
rect 21913 15453 21925 15487
rect 21959 15453 21971 15487
rect 21913 15447 21971 15453
rect 22186 15444 22192 15496
rect 22244 15484 22250 15496
rect 22462 15484 22468 15496
rect 22244 15456 22468 15484
rect 22244 15444 22250 15456
rect 22462 15444 22468 15456
rect 22520 15444 22526 15496
rect 23014 15444 23020 15496
rect 23072 15484 23078 15496
rect 23308 15493 23336 15524
rect 24210 15512 24216 15564
rect 24268 15552 24274 15564
rect 24857 15555 24915 15561
rect 24857 15552 24869 15555
rect 24268 15524 24869 15552
rect 24268 15512 24274 15524
rect 24857 15521 24869 15524
rect 24903 15552 24915 15555
rect 26510 15552 26516 15564
rect 24903 15524 26004 15552
rect 24903 15521 24915 15524
rect 24857 15515 24915 15521
rect 23109 15487 23167 15493
rect 23109 15484 23121 15487
rect 23072 15456 23121 15484
rect 23072 15444 23078 15456
rect 23109 15453 23121 15456
rect 23155 15453 23167 15487
rect 23109 15447 23167 15453
rect 23293 15487 23351 15493
rect 23293 15453 23305 15487
rect 23339 15453 23351 15487
rect 23293 15447 23351 15453
rect 23477 15487 23535 15493
rect 23477 15453 23489 15487
rect 23523 15484 23535 15487
rect 24394 15484 24400 15496
rect 23523 15456 24400 15484
rect 23523 15453 23535 15456
rect 23477 15447 23535 15453
rect 24394 15444 24400 15456
rect 24452 15484 24458 15496
rect 24765 15487 24823 15493
rect 24765 15484 24777 15487
rect 24452 15456 24777 15484
rect 24452 15444 24458 15456
rect 24765 15453 24777 15456
rect 24811 15453 24823 15487
rect 24765 15447 24823 15453
rect 25498 15444 25504 15496
rect 25556 15484 25562 15496
rect 25869 15487 25927 15493
rect 25869 15484 25881 15487
rect 25556 15456 25881 15484
rect 25556 15444 25562 15456
rect 25869 15453 25881 15456
rect 25915 15453 25927 15487
rect 25869 15447 25927 15453
rect 25314 15416 25320 15428
rect 21284 15388 25320 15416
rect 17828 15376 17834 15388
rect 25314 15376 25320 15388
rect 25372 15376 25378 15428
rect 15289 15351 15347 15357
rect 15289 15317 15301 15351
rect 15335 15348 15347 15351
rect 15930 15348 15936 15360
rect 15335 15320 15936 15348
rect 15335 15317 15347 15320
rect 15289 15311 15347 15317
rect 15930 15308 15936 15320
rect 15988 15308 15994 15360
rect 17678 15348 17684 15360
rect 17639 15320 17684 15348
rect 17678 15308 17684 15320
rect 17736 15308 17742 15360
rect 20162 15308 20168 15360
rect 20220 15348 20226 15360
rect 20257 15351 20315 15357
rect 20257 15348 20269 15351
rect 20220 15320 20269 15348
rect 20220 15308 20226 15320
rect 20257 15317 20269 15320
rect 20303 15317 20315 15351
rect 25130 15348 25136 15360
rect 25091 15320 25136 15348
rect 20257 15311 20315 15317
rect 25130 15308 25136 15320
rect 25188 15308 25194 15360
rect 25976 15348 26004 15524
rect 26068 15524 26516 15552
rect 26068 15493 26096 15524
rect 26510 15512 26516 15524
rect 26568 15512 26574 15564
rect 30024 15552 30052 15592
rect 33134 15580 33140 15632
rect 33192 15620 33198 15632
rect 33321 15623 33379 15629
rect 33321 15620 33333 15623
rect 33192 15592 33333 15620
rect 33192 15580 33198 15592
rect 33321 15589 33333 15592
rect 33367 15589 33379 15623
rect 33321 15583 33379 15589
rect 29748 15524 30052 15552
rect 29748 15496 29776 15524
rect 30834 15512 30840 15564
rect 30892 15552 30898 15564
rect 31570 15552 31576 15564
rect 30892 15524 31576 15552
rect 30892 15512 30898 15524
rect 31570 15512 31576 15524
rect 31628 15512 31634 15564
rect 31665 15555 31723 15561
rect 31665 15521 31677 15555
rect 31711 15521 31723 15555
rect 33336 15552 33364 15583
rect 33502 15580 33508 15632
rect 33560 15620 33566 15632
rect 34149 15623 34207 15629
rect 34149 15620 34161 15623
rect 33560 15592 34161 15620
rect 33560 15580 33566 15592
rect 34149 15589 34161 15592
rect 34195 15589 34207 15623
rect 34149 15583 34207 15589
rect 33873 15555 33931 15561
rect 33873 15552 33885 15555
rect 33336 15524 33885 15552
rect 31665 15515 31723 15521
rect 33873 15521 33885 15524
rect 33919 15521 33931 15555
rect 38102 15552 38108 15564
rect 38063 15524 38108 15552
rect 33873 15515 33931 15521
rect 26053 15487 26111 15493
rect 26053 15453 26065 15487
rect 26099 15453 26111 15487
rect 26053 15447 26111 15453
rect 26145 15487 26203 15493
rect 26145 15453 26157 15487
rect 26191 15453 26203 15487
rect 26970 15484 26976 15496
rect 26931 15456 26976 15484
rect 26145 15447 26203 15453
rect 26160 15416 26188 15447
rect 26970 15444 26976 15456
rect 27028 15444 27034 15496
rect 27154 15484 27160 15496
rect 27115 15456 27160 15484
rect 27154 15444 27160 15456
rect 27212 15444 27218 15496
rect 28074 15484 28080 15496
rect 28035 15456 28080 15484
rect 28074 15444 28080 15456
rect 28132 15444 28138 15496
rect 28166 15444 28172 15496
rect 28224 15484 28230 15496
rect 28261 15487 28319 15493
rect 28261 15484 28273 15487
rect 28224 15456 28273 15484
rect 28224 15444 28230 15456
rect 28261 15453 28273 15456
rect 28307 15453 28319 15487
rect 28261 15447 28319 15453
rect 28537 15487 28595 15493
rect 28537 15453 28549 15487
rect 28583 15484 28595 15487
rect 28626 15484 28632 15496
rect 28583 15456 28632 15484
rect 28583 15453 28595 15456
rect 28537 15447 28595 15453
rect 28552 15416 28580 15447
rect 28626 15444 28632 15456
rect 28684 15444 28690 15496
rect 29730 15484 29736 15496
rect 29643 15456 29736 15484
rect 29730 15444 29736 15456
rect 29788 15444 29794 15496
rect 29822 15444 29828 15496
rect 29880 15484 29886 15496
rect 29917 15487 29975 15493
rect 29917 15484 29929 15487
rect 29880 15456 29929 15484
rect 29880 15444 29886 15456
rect 29917 15453 29929 15456
rect 29963 15453 29975 15487
rect 29917 15447 29975 15453
rect 26160 15388 28580 15416
rect 31680 15416 31708 15515
rect 38102 15512 38108 15524
rect 38160 15512 38166 15564
rect 32953 15487 33011 15493
rect 32953 15453 32965 15487
rect 32999 15484 33011 15487
rect 33502 15484 33508 15496
rect 32999 15456 33508 15484
rect 32999 15453 33011 15456
rect 32953 15447 33011 15453
rect 33502 15444 33508 15456
rect 33560 15444 33566 15496
rect 34790 15444 34796 15496
rect 34848 15484 34854 15496
rect 34977 15487 35035 15493
rect 34977 15484 34989 15487
rect 34848 15456 34989 15484
rect 34848 15444 34854 15456
rect 34977 15453 34989 15456
rect 35023 15453 35035 15487
rect 37826 15484 37832 15496
rect 37787 15456 37832 15484
rect 34977 15447 35035 15453
rect 37826 15444 37832 15456
rect 37884 15444 37890 15496
rect 31680 15388 34652 15416
rect 28445 15351 28503 15357
rect 28445 15348 28457 15351
rect 25976 15320 28457 15348
rect 28445 15317 28457 15320
rect 28491 15348 28503 15351
rect 28718 15348 28724 15360
rect 28491 15320 28724 15348
rect 28491 15317 28503 15320
rect 28445 15311 28503 15317
rect 28718 15308 28724 15320
rect 28776 15308 28782 15360
rect 31110 15348 31116 15360
rect 31071 15320 31116 15348
rect 31110 15308 31116 15320
rect 31168 15308 31174 15360
rect 31481 15351 31539 15357
rect 31481 15317 31493 15351
rect 31527 15348 31539 15351
rect 31662 15348 31668 15360
rect 31527 15320 31668 15348
rect 31527 15317 31539 15320
rect 31481 15311 31539 15317
rect 31662 15308 31668 15320
rect 31720 15308 31726 15360
rect 33410 15348 33416 15360
rect 33371 15320 33416 15348
rect 33410 15308 33416 15320
rect 33468 15308 33474 15360
rect 33502 15308 33508 15360
rect 33560 15348 33566 15360
rect 34333 15351 34391 15357
rect 34333 15348 34345 15351
rect 33560 15320 34345 15348
rect 33560 15308 33566 15320
rect 34333 15317 34345 15320
rect 34379 15317 34391 15351
rect 34624 15348 34652 15388
rect 34698 15376 34704 15428
rect 34756 15416 34762 15428
rect 35222 15419 35280 15425
rect 35222 15416 35234 15419
rect 34756 15388 35234 15416
rect 34756 15376 34762 15388
rect 35222 15385 35234 15388
rect 35268 15385 35280 15419
rect 35222 15379 35280 15385
rect 38010 15348 38016 15360
rect 34624 15320 38016 15348
rect 34333 15311 34391 15317
rect 38010 15308 38016 15320
rect 38068 15308 38074 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 8846 15144 8852 15156
rect 8807 15116 8852 15144
rect 8846 15104 8852 15116
rect 8904 15104 8910 15156
rect 10042 15144 10048 15156
rect 10003 15116 10048 15144
rect 10042 15104 10048 15116
rect 10100 15104 10106 15156
rect 13725 15147 13783 15153
rect 13725 15113 13737 15147
rect 13771 15144 13783 15147
rect 14458 15144 14464 15156
rect 13771 15116 14464 15144
rect 13771 15113 13783 15116
rect 13725 15107 13783 15113
rect 14458 15104 14464 15116
rect 14516 15104 14522 15156
rect 16022 15144 16028 15156
rect 15120 15116 16028 15144
rect 15120 15076 15148 15116
rect 16022 15104 16028 15116
rect 16080 15104 16086 15156
rect 16758 15104 16764 15156
rect 16816 15144 16822 15156
rect 18969 15147 19027 15153
rect 18969 15144 18981 15147
rect 16816 15116 18981 15144
rect 16816 15104 16822 15116
rect 18969 15113 18981 15116
rect 19015 15113 19027 15147
rect 18969 15107 19027 15113
rect 20346 15104 20352 15156
rect 20404 15144 20410 15156
rect 20404 15116 25728 15144
rect 20404 15104 20410 15116
rect 11808 15048 15148 15076
rect 8757 15011 8815 15017
rect 8757 14977 8769 15011
rect 8803 15008 8815 15011
rect 9306 15008 9312 15020
rect 8803 14980 9312 15008
rect 8803 14977 8815 14980
rect 8757 14971 8815 14977
rect 9306 14968 9312 14980
rect 9364 14968 9370 15020
rect 10134 14968 10140 15020
rect 10192 15008 10198 15020
rect 10229 15011 10287 15017
rect 10229 15008 10241 15011
rect 10192 14980 10241 15008
rect 10192 14968 10198 14980
rect 10229 14977 10241 14980
rect 10275 14977 10287 15011
rect 10229 14971 10287 14977
rect 10505 15011 10563 15017
rect 10505 14977 10517 15011
rect 10551 15008 10563 15011
rect 11146 15008 11152 15020
rect 10551 14980 11152 15008
rect 10551 14977 10563 14980
rect 10505 14971 10563 14977
rect 11146 14968 11152 14980
rect 11204 14968 11210 15020
rect 11808 15017 11836 15048
rect 16574 15036 16580 15088
rect 16632 15076 16638 15088
rect 17862 15076 17868 15088
rect 16632 15048 17264 15076
rect 16632 15036 16638 15048
rect 11793 15011 11851 15017
rect 11793 14977 11805 15011
rect 11839 15008 11851 15011
rect 11882 15008 11888 15020
rect 11839 14980 11888 15008
rect 11839 14977 11851 14980
rect 11793 14971 11851 14977
rect 11882 14968 11888 14980
rect 11940 14968 11946 15020
rect 13354 15008 13360 15020
rect 13315 14980 13360 15008
rect 13354 14968 13360 14980
rect 13412 14968 13418 15020
rect 15013 15011 15071 15017
rect 15013 14977 15025 15011
rect 15059 14977 15071 15011
rect 15194 15008 15200 15020
rect 15155 14980 15200 15008
rect 15013 14971 15071 14977
rect 8294 14900 8300 14952
rect 8352 14940 8358 14952
rect 9033 14943 9091 14949
rect 9033 14940 9045 14943
rect 8352 14912 9045 14940
rect 8352 14900 8358 14912
rect 9033 14909 9045 14912
rect 9079 14940 9091 14943
rect 10413 14943 10471 14949
rect 10413 14940 10425 14943
rect 9079 14912 10425 14940
rect 9079 14909 9091 14912
rect 9033 14903 9091 14909
rect 10413 14909 10425 14912
rect 10459 14909 10471 14943
rect 10413 14903 10471 14909
rect 10594 14900 10600 14952
rect 10652 14940 10658 14952
rect 11701 14943 11759 14949
rect 11701 14940 11713 14943
rect 10652 14912 11713 14940
rect 10652 14900 10658 14912
rect 11701 14909 11713 14912
rect 11747 14909 11759 14943
rect 11701 14903 11759 14909
rect 12253 14943 12311 14949
rect 12253 14909 12265 14943
rect 12299 14940 12311 14943
rect 13446 14940 13452 14952
rect 12299 14912 12434 14940
rect 13407 14912 13452 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 12406 14872 12434 14912
rect 13446 14900 13452 14912
rect 13504 14900 13510 14952
rect 15028 14940 15056 14971
rect 15194 14968 15200 14980
rect 15252 14968 15258 15020
rect 15930 15008 15936 15020
rect 15891 14980 15936 15008
rect 15930 14968 15936 14980
rect 15988 14968 15994 15020
rect 16301 15011 16359 15017
rect 16301 14977 16313 15011
rect 16347 15008 16359 15011
rect 16850 15008 16856 15020
rect 16347 14980 16856 15008
rect 16347 14977 16359 14980
rect 16301 14971 16359 14977
rect 16850 14968 16856 14980
rect 16908 14968 16914 15020
rect 17034 14968 17040 15020
rect 17092 15017 17098 15020
rect 17236 15017 17264 15048
rect 17512 15048 17868 15076
rect 17092 15011 17141 15017
rect 17092 14977 17095 15011
rect 17129 14977 17141 15011
rect 17092 14971 17141 14977
rect 17221 15011 17279 15017
rect 17221 14977 17233 15011
rect 17267 14977 17279 15011
rect 17221 14971 17279 14977
rect 17334 15014 17392 15020
rect 17512 15017 17540 15048
rect 17862 15036 17868 15048
rect 17920 15036 17926 15088
rect 18046 15036 18052 15088
rect 18104 15076 18110 15088
rect 21082 15076 21088 15088
rect 18104 15048 19656 15076
rect 21043 15048 21088 15076
rect 18104 15036 18110 15048
rect 17334 14980 17346 15014
rect 17380 15011 17392 15014
rect 17497 15011 17555 15017
rect 17380 14983 17448 15011
rect 17380 14980 17392 14983
rect 17334 14974 17392 14980
rect 17092 14968 17098 14971
rect 17420 14940 17448 14983
rect 17497 14977 17509 15011
rect 17543 14977 17555 15011
rect 17497 14971 17555 14977
rect 17586 14968 17592 15020
rect 17644 15008 17650 15020
rect 17770 15008 17776 15020
rect 17644 14980 17776 15008
rect 17644 14968 17650 14980
rect 17770 14968 17776 14980
rect 17828 14968 17834 15020
rect 18874 14968 18880 15020
rect 18932 15008 18938 15020
rect 19199 15011 19257 15017
rect 19199 15008 19211 15011
rect 18932 14980 19211 15008
rect 18932 14968 18938 14980
rect 19199 14977 19211 14980
rect 19245 14977 19257 15011
rect 19334 15008 19340 15020
rect 19295 14980 19340 15008
rect 19199 14971 19257 14977
rect 19334 14968 19340 14980
rect 19392 14968 19398 15020
rect 19426 14968 19432 15020
rect 19484 15008 19490 15020
rect 19628 15017 19656 15048
rect 21082 15036 21088 15048
rect 21140 15036 21146 15088
rect 19613 15011 19671 15017
rect 19484 14980 19529 15008
rect 19484 14968 19490 14980
rect 19613 14977 19625 15011
rect 19659 14977 19671 15011
rect 19613 14971 19671 14977
rect 20714 14968 20720 15020
rect 20772 15008 20778 15020
rect 20809 15011 20867 15017
rect 20809 15008 20821 15011
rect 20772 14980 20821 15008
rect 20772 14968 20778 14980
rect 20809 14977 20821 14980
rect 20855 14977 20867 15011
rect 20809 14971 20867 14977
rect 20993 15011 21051 15017
rect 20993 14977 21005 15011
rect 21039 14977 21051 15011
rect 20993 14971 21051 14977
rect 21229 15011 21287 15017
rect 21229 14977 21241 15011
rect 21275 15008 21287 15011
rect 21910 15008 21916 15020
rect 21275 14980 21916 15008
rect 21275 14977 21287 14980
rect 21229 14971 21287 14977
rect 17862 14940 17868 14952
rect 15028 14912 16988 14940
rect 17420 14912 17868 14940
rect 12526 14872 12532 14884
rect 12406 14844 12532 14872
rect 12526 14832 12532 14844
rect 12584 14872 12590 14884
rect 13538 14872 13544 14884
rect 12584 14844 13544 14872
rect 12584 14832 12590 14844
rect 13538 14832 13544 14844
rect 13596 14832 13602 14884
rect 15378 14872 15384 14884
rect 15339 14844 15384 14872
rect 15378 14832 15384 14844
rect 15436 14832 15442 14884
rect 8386 14804 8392 14816
rect 8347 14776 8392 14804
rect 8386 14764 8392 14776
rect 8444 14764 8450 14816
rect 11146 14764 11152 14816
rect 11204 14804 11210 14816
rect 15286 14804 15292 14816
rect 11204 14776 15292 14804
rect 11204 14764 11210 14776
rect 15286 14764 15292 14776
rect 15344 14764 15350 14816
rect 16666 14764 16672 14816
rect 16724 14804 16730 14816
rect 16853 14807 16911 14813
rect 16853 14804 16865 14807
rect 16724 14776 16865 14804
rect 16724 14764 16730 14776
rect 16853 14773 16865 14776
rect 16899 14773 16911 14807
rect 16960 14804 16988 14912
rect 17862 14900 17868 14912
rect 17920 14900 17926 14952
rect 17954 14900 17960 14952
rect 18012 14940 18018 14952
rect 19702 14940 19708 14952
rect 18012 14912 19708 14940
rect 18012 14900 18018 14912
rect 19702 14900 19708 14912
rect 19760 14900 19766 14952
rect 17972 14872 18000 14900
rect 18322 14872 18328 14884
rect 17236 14844 18000 14872
rect 18235 14844 18328 14872
rect 17236 14804 17264 14844
rect 18322 14832 18328 14844
rect 18380 14872 18386 14884
rect 20346 14872 20352 14884
rect 18380 14844 20352 14872
rect 18380 14832 18386 14844
rect 20346 14832 20352 14844
rect 20404 14832 20410 14884
rect 20824 14872 20852 14971
rect 21008 14940 21036 14971
rect 21910 14968 21916 14980
rect 21968 14968 21974 15020
rect 22005 15011 22063 15017
rect 22005 14977 22017 15011
rect 22051 15008 22063 15011
rect 22112 15008 22140 15116
rect 25130 15036 25136 15088
rect 25188 15076 25194 15088
rect 25700 15085 25728 15116
rect 31570 15104 31576 15156
rect 31628 15144 31634 15156
rect 31628 15116 37872 15144
rect 31628 15104 31634 15116
rect 25593 15079 25651 15085
rect 25593 15076 25605 15079
rect 25188 15048 25605 15076
rect 25188 15036 25194 15048
rect 25593 15045 25605 15048
rect 25639 15045 25651 15079
rect 25593 15039 25651 15045
rect 25685 15079 25743 15085
rect 25685 15045 25697 15079
rect 25731 15076 25743 15079
rect 26234 15076 26240 15088
rect 25731 15048 26240 15076
rect 25731 15045 25743 15048
rect 25685 15039 25743 15045
rect 26234 15036 26240 15048
rect 26292 15036 26298 15088
rect 31478 15076 31484 15088
rect 31439 15048 31484 15076
rect 31478 15036 31484 15048
rect 31536 15036 31542 15088
rect 33410 15036 33416 15088
rect 33468 15076 33474 15088
rect 33468 15048 33732 15076
rect 33468 15036 33474 15048
rect 22462 15017 22468 15020
rect 22051 14980 22140 15008
rect 22189 15011 22247 15017
rect 22051 14977 22063 14980
rect 22005 14971 22063 14977
rect 22189 14977 22201 15011
rect 22235 14977 22247 15011
rect 22189 14971 22247 14977
rect 22281 15011 22339 15017
rect 22281 14977 22293 15011
rect 22327 14977 22339 15011
rect 22281 14971 22339 14977
rect 22425 15011 22468 15017
rect 22425 14977 22437 15011
rect 22425 14971 22468 14977
rect 21450 14940 21456 14952
rect 21008 14912 21456 14940
rect 21450 14900 21456 14912
rect 21508 14940 21514 14952
rect 21634 14940 21640 14952
rect 21508 14912 21640 14940
rect 21508 14900 21514 14912
rect 21634 14900 21640 14912
rect 21692 14940 21698 14952
rect 22204 14940 22232 14971
rect 21692 14912 22232 14940
rect 22296 14940 22324 14971
rect 22462 14968 22468 14971
rect 22520 14968 22526 15020
rect 22554 14968 22560 15020
rect 22612 15017 22618 15020
rect 22612 15011 22632 15017
rect 22620 14977 22632 15011
rect 22612 14971 22632 14977
rect 22612 14968 22618 14971
rect 23658 14968 23664 15020
rect 23716 15008 23722 15020
rect 24210 15008 24216 15020
rect 23716 14980 24216 15008
rect 23716 14968 23722 14980
rect 24210 14968 24216 14980
rect 24268 14968 24274 15020
rect 24489 15011 24547 15017
rect 24489 14977 24501 15011
rect 24535 15008 24547 15011
rect 24578 15008 24584 15020
rect 24535 14980 24584 15008
rect 24535 14977 24547 14980
rect 24489 14971 24547 14977
rect 24578 14968 24584 14980
rect 24636 15008 24642 15020
rect 24946 15008 24952 15020
rect 24636 14980 24952 15008
rect 24636 14968 24642 14980
rect 24946 14968 24952 14980
rect 25004 14968 25010 15020
rect 25406 15008 25412 15020
rect 25367 14980 25412 15008
rect 25406 14968 25412 14980
rect 25464 14968 25470 15020
rect 25774 14968 25780 15020
rect 25832 15017 25838 15020
rect 25832 15008 25840 15017
rect 27798 15008 27804 15020
rect 25832 14980 25877 15008
rect 27759 14980 27804 15008
rect 25832 14971 25840 14980
rect 25832 14968 25838 14971
rect 27798 14968 27804 14980
rect 27856 14968 27862 15020
rect 28074 14968 28080 15020
rect 28132 15008 28138 15020
rect 28169 15011 28227 15017
rect 28169 15008 28181 15011
rect 28132 14980 28181 15008
rect 28132 14968 28138 14980
rect 28169 14977 28181 14980
rect 28215 14977 28227 15011
rect 28169 14971 28227 14977
rect 31205 15011 31263 15017
rect 31205 14977 31217 15011
rect 31251 15008 31263 15011
rect 32306 15008 32312 15020
rect 31251 14980 32312 15008
rect 31251 14977 31263 14980
rect 31205 14971 31263 14977
rect 32306 14968 32312 14980
rect 32364 14968 32370 15020
rect 33502 15008 33508 15020
rect 33463 14980 33508 15008
rect 33502 14968 33508 14980
rect 33560 14968 33566 15020
rect 33704 15017 33732 15048
rect 37844 15017 37872 15116
rect 38102 15076 38108 15088
rect 38063 15048 38108 15076
rect 38102 15036 38108 15048
rect 38160 15036 38166 15088
rect 33689 15011 33747 15017
rect 33689 14977 33701 15011
rect 33735 14977 33747 15011
rect 33689 14971 33747 14977
rect 37829 15011 37887 15017
rect 37829 14977 37841 15011
rect 37875 14977 37887 15011
rect 37829 14971 37887 14977
rect 27430 14940 27436 14952
rect 22296 14912 27436 14940
rect 21692 14900 21698 14912
rect 27430 14900 27436 14912
rect 27488 14900 27494 14952
rect 27617 14943 27675 14949
rect 27617 14909 27629 14943
rect 27663 14940 27675 14943
rect 29086 14940 29092 14952
rect 27663 14912 29092 14940
rect 27663 14909 27675 14912
rect 27617 14903 27675 14909
rect 29086 14900 29092 14912
rect 29144 14940 29150 14952
rect 30650 14940 30656 14952
rect 29144 14912 30656 14940
rect 29144 14900 29150 14912
rect 30650 14900 30656 14912
rect 30708 14900 30714 14952
rect 23934 14872 23940 14884
rect 20824 14844 23940 14872
rect 23934 14832 23940 14844
rect 23992 14832 23998 14884
rect 25038 14832 25044 14884
rect 25096 14872 25102 14884
rect 28077 14875 28135 14881
rect 28077 14872 28089 14875
rect 25096 14844 28089 14872
rect 25096 14832 25102 14844
rect 28077 14841 28089 14844
rect 28123 14841 28135 14875
rect 28077 14835 28135 14841
rect 28994 14832 29000 14884
rect 29052 14872 29058 14884
rect 32122 14872 32128 14884
rect 29052 14844 32128 14872
rect 29052 14832 29058 14844
rect 32122 14832 32128 14844
rect 32180 14872 32186 14884
rect 35434 14872 35440 14884
rect 32180 14844 35440 14872
rect 32180 14832 32186 14844
rect 35434 14832 35440 14844
rect 35492 14832 35498 14884
rect 16960 14776 17264 14804
rect 16853 14767 16911 14773
rect 17770 14764 17776 14816
rect 17828 14804 17834 14816
rect 18417 14807 18475 14813
rect 18417 14804 18429 14807
rect 17828 14776 18429 14804
rect 17828 14764 17834 14776
rect 18417 14773 18429 14776
rect 18463 14773 18475 14807
rect 18417 14767 18475 14773
rect 20714 14764 20720 14816
rect 20772 14804 20778 14816
rect 21361 14807 21419 14813
rect 21361 14804 21373 14807
rect 20772 14776 21373 14804
rect 20772 14764 20778 14776
rect 21361 14773 21373 14776
rect 21407 14773 21419 14807
rect 21361 14767 21419 14773
rect 24029 14807 24087 14813
rect 24029 14773 24041 14807
rect 24075 14804 24087 14807
rect 24118 14804 24124 14816
rect 24075 14776 24124 14804
rect 24075 14773 24087 14776
rect 24029 14767 24087 14773
rect 24118 14764 24124 14776
rect 24176 14764 24182 14816
rect 24394 14804 24400 14816
rect 24355 14776 24400 14804
rect 24394 14764 24400 14776
rect 24452 14764 24458 14816
rect 25961 14807 26019 14813
rect 25961 14773 25973 14807
rect 26007 14804 26019 14807
rect 27890 14804 27896 14816
rect 26007 14776 27896 14804
rect 26007 14773 26019 14776
rect 25961 14767 26019 14773
rect 27890 14764 27896 14776
rect 27948 14764 27954 14816
rect 33505 14807 33563 14813
rect 33505 14773 33517 14807
rect 33551 14804 33563 14807
rect 33962 14804 33968 14816
rect 33551 14776 33968 14804
rect 33551 14773 33563 14776
rect 33505 14767 33563 14773
rect 33962 14764 33968 14776
rect 34020 14764 34026 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 13446 14600 13452 14612
rect 13407 14572 13452 14600
rect 13446 14560 13452 14572
rect 13504 14560 13510 14612
rect 16574 14560 16580 14612
rect 16632 14600 16638 14612
rect 17129 14603 17187 14609
rect 17129 14600 17141 14603
rect 16632 14572 17141 14600
rect 16632 14560 16638 14572
rect 17129 14569 17141 14572
rect 17175 14569 17187 14603
rect 17129 14563 17187 14569
rect 19334 14560 19340 14612
rect 19392 14600 19398 14612
rect 19521 14603 19579 14609
rect 19521 14600 19533 14603
rect 19392 14572 19533 14600
rect 19392 14560 19398 14572
rect 19521 14569 19533 14572
rect 19567 14569 19579 14603
rect 19521 14563 19579 14569
rect 19702 14560 19708 14612
rect 19760 14600 19766 14612
rect 25038 14600 25044 14612
rect 19760 14572 25044 14600
rect 19760 14560 19766 14572
rect 25038 14560 25044 14572
rect 25096 14560 25102 14612
rect 25406 14600 25412 14612
rect 25367 14572 25412 14600
rect 25406 14560 25412 14572
rect 25464 14560 25470 14612
rect 27798 14600 27804 14612
rect 27759 14572 27804 14600
rect 27798 14560 27804 14572
rect 27856 14560 27862 14612
rect 28810 14560 28816 14612
rect 28868 14600 28874 14612
rect 34885 14603 34943 14609
rect 28868 14572 31754 14600
rect 28868 14560 28874 14572
rect 15930 14492 15936 14544
rect 15988 14532 15994 14544
rect 15988 14504 18920 14532
rect 15988 14492 15994 14504
rect 6914 14424 6920 14476
rect 6972 14464 6978 14476
rect 7926 14464 7932 14476
rect 6972 14436 7932 14464
rect 6972 14424 6978 14436
rect 7926 14424 7932 14436
rect 7984 14464 7990 14476
rect 8389 14467 8447 14473
rect 8389 14464 8401 14467
rect 7984 14436 8401 14464
rect 7984 14424 7990 14436
rect 8389 14433 8401 14436
rect 8435 14433 8447 14467
rect 12434 14464 12440 14476
rect 8389 14427 8447 14433
rect 8680 14436 12440 14464
rect 7374 14356 7380 14408
rect 7432 14396 7438 14408
rect 7653 14399 7711 14405
rect 7653 14396 7665 14399
rect 7432 14368 7665 14396
rect 7432 14356 7438 14368
rect 7653 14365 7665 14368
rect 7699 14396 7711 14399
rect 8680 14396 8708 14436
rect 12434 14424 12440 14436
rect 12492 14424 12498 14476
rect 16390 14464 16396 14476
rect 13096 14436 16396 14464
rect 11882 14396 11888 14408
rect 7699 14368 8708 14396
rect 11843 14368 11888 14396
rect 7699 14365 7711 14368
rect 7653 14359 7711 14365
rect 11882 14356 11888 14368
rect 11940 14356 11946 14408
rect 12066 14396 12072 14408
rect 12027 14368 12072 14396
rect 12066 14356 12072 14368
rect 12124 14356 12130 14408
rect 12253 14399 12311 14405
rect 12253 14365 12265 14399
rect 12299 14396 12311 14399
rect 13096 14396 13124 14436
rect 12299 14368 13124 14396
rect 12299 14365 12311 14368
rect 12253 14359 12311 14365
rect 13170 14356 13176 14408
rect 13228 14396 13234 14408
rect 13357 14399 13415 14405
rect 13357 14396 13369 14399
rect 13228 14368 13369 14396
rect 13228 14356 13234 14368
rect 13357 14365 13369 14368
rect 13403 14365 13415 14399
rect 13357 14359 13415 14365
rect 13541 14399 13599 14405
rect 13541 14365 13553 14399
rect 13587 14396 13599 14399
rect 14642 14396 14648 14408
rect 13587 14368 14648 14396
rect 13587 14365 13599 14368
rect 13541 14359 13599 14365
rect 12986 14288 12992 14340
rect 13044 14328 13050 14340
rect 13556 14328 13584 14359
rect 14642 14356 14648 14368
rect 14700 14356 14706 14408
rect 15212 14405 15240 14436
rect 16390 14424 16396 14436
rect 16448 14464 16454 14476
rect 17770 14464 17776 14476
rect 16448 14436 17632 14464
rect 17731 14436 17776 14464
rect 16448 14424 16454 14436
rect 15197 14399 15255 14405
rect 15197 14365 15209 14399
rect 15243 14365 15255 14399
rect 15197 14359 15255 14365
rect 16850 14356 16856 14408
rect 16908 14396 16914 14408
rect 17218 14396 17224 14408
rect 16908 14368 17224 14396
rect 16908 14356 16914 14368
rect 17218 14356 17224 14368
rect 17276 14396 17282 14408
rect 17497 14399 17555 14405
rect 17497 14396 17509 14399
rect 17276 14368 17509 14396
rect 17276 14356 17282 14368
rect 17497 14365 17509 14368
rect 17543 14365 17555 14399
rect 17604 14396 17632 14436
rect 17770 14424 17776 14436
rect 17828 14424 17834 14476
rect 18046 14396 18052 14408
rect 17604 14368 18052 14396
rect 17497 14359 17555 14365
rect 18046 14356 18052 14368
rect 18104 14356 18110 14408
rect 18892 14405 18920 14504
rect 20898 14492 20904 14544
rect 20956 14532 20962 14544
rect 22005 14535 22063 14541
rect 22005 14532 22017 14535
rect 20956 14504 22017 14532
rect 20956 14492 20962 14504
rect 22005 14501 22017 14504
rect 22051 14501 22063 14535
rect 22005 14495 22063 14501
rect 24394 14492 24400 14544
rect 24452 14532 24458 14544
rect 29181 14535 29239 14541
rect 24452 14504 28764 14532
rect 24452 14492 24458 14504
rect 20162 14464 20168 14476
rect 20123 14436 20168 14464
rect 20162 14424 20168 14436
rect 20220 14424 20226 14476
rect 22738 14424 22744 14476
rect 22796 14464 22802 14476
rect 22796 14436 23704 14464
rect 22796 14424 22802 14436
rect 18693 14399 18751 14405
rect 18693 14365 18705 14399
rect 18739 14365 18751 14399
rect 18693 14359 18751 14365
rect 18877 14399 18935 14405
rect 18877 14365 18889 14399
rect 18923 14396 18935 14399
rect 18966 14396 18972 14408
rect 18923 14368 18972 14396
rect 18923 14365 18935 14368
rect 18877 14359 18935 14365
rect 13044 14300 13584 14328
rect 13044 14288 13050 14300
rect 15286 14288 15292 14340
rect 15344 14328 15350 14340
rect 15473 14331 15531 14337
rect 15473 14328 15485 14331
rect 15344 14300 15485 14328
rect 15344 14288 15350 14300
rect 15473 14297 15485 14300
rect 15519 14297 15531 14331
rect 15473 14291 15531 14297
rect 17589 14331 17647 14337
rect 17589 14297 17601 14331
rect 17635 14328 17647 14331
rect 17678 14328 17684 14340
rect 17635 14300 17684 14328
rect 17635 14297 17647 14300
rect 17589 14291 17647 14297
rect 17678 14288 17684 14300
rect 17736 14328 17742 14340
rect 18708 14328 18736 14359
rect 18966 14356 18972 14368
rect 19024 14356 19030 14408
rect 19150 14356 19156 14408
rect 19208 14396 19214 14408
rect 21450 14396 21456 14408
rect 19208 14368 21456 14396
rect 19208 14356 19214 14368
rect 21450 14356 21456 14368
rect 21508 14356 21514 14408
rect 21634 14396 21640 14408
rect 21595 14368 21640 14396
rect 21634 14356 21640 14368
rect 21692 14356 21698 14408
rect 21910 14405 21916 14408
rect 21873 14399 21916 14405
rect 21873 14396 21885 14399
rect 21823 14368 21885 14396
rect 21873 14365 21885 14368
rect 21968 14396 21974 14408
rect 22186 14396 22192 14408
rect 21968 14368 22192 14396
rect 21873 14359 21916 14365
rect 21910 14356 21916 14359
rect 21968 14356 21974 14368
rect 22186 14356 22192 14368
rect 22244 14356 22250 14408
rect 23566 14405 23572 14408
rect 23549 14399 23572 14405
rect 23549 14365 23561 14399
rect 23549 14359 23572 14365
rect 23566 14356 23572 14359
rect 23624 14356 23630 14408
rect 23676 14405 23704 14436
rect 23934 14424 23940 14476
rect 23992 14464 23998 14476
rect 24029 14467 24087 14473
rect 24029 14464 24041 14467
rect 23992 14436 24041 14464
rect 23992 14424 23998 14436
rect 24029 14433 24041 14436
rect 24075 14433 24087 14467
rect 24029 14427 24087 14433
rect 24118 14424 24124 14476
rect 24176 14464 24182 14476
rect 28736 14473 28764 14504
rect 29181 14501 29193 14535
rect 29227 14532 29239 14535
rect 31726 14532 31754 14572
rect 34885 14569 34897 14603
rect 34931 14600 34943 14603
rect 35342 14600 35348 14612
rect 34931 14572 35348 14600
rect 34931 14569 34943 14572
rect 34885 14563 34943 14569
rect 35342 14560 35348 14572
rect 35400 14560 35406 14612
rect 37918 14560 37924 14612
rect 37976 14600 37982 14612
rect 38289 14603 38347 14609
rect 38289 14600 38301 14603
rect 37976 14572 38301 14600
rect 37976 14560 37982 14572
rect 38289 14569 38301 14572
rect 38335 14569 38347 14603
rect 38289 14563 38347 14569
rect 35618 14532 35624 14544
rect 29227 14504 29868 14532
rect 31726 14504 35624 14532
rect 29227 14501 29239 14504
rect 29181 14495 29239 14501
rect 29840 14473 29868 14504
rect 35618 14492 35624 14504
rect 35676 14492 35682 14544
rect 28721 14467 28779 14473
rect 24176 14436 25452 14464
rect 24176 14424 24182 14436
rect 23661 14399 23719 14405
rect 23661 14365 23673 14399
rect 23707 14365 23719 14399
rect 24578 14396 24584 14408
rect 24539 14368 24584 14396
rect 23661 14359 23719 14365
rect 24578 14356 24584 14368
rect 24636 14356 24642 14408
rect 24765 14399 24823 14405
rect 24765 14365 24777 14399
rect 24811 14396 24823 14399
rect 25038 14396 25044 14408
rect 24811 14368 25044 14396
rect 24811 14365 24823 14368
rect 24765 14359 24823 14365
rect 25038 14356 25044 14368
rect 25096 14356 25102 14408
rect 25424 14405 25452 14436
rect 28721 14433 28733 14467
rect 28767 14433 28779 14467
rect 28721 14427 28779 14433
rect 29825 14467 29883 14473
rect 29825 14433 29837 14467
rect 29871 14433 29883 14467
rect 33318 14464 33324 14476
rect 33279 14436 33324 14464
rect 29825 14427 29883 14433
rect 33318 14424 33324 14436
rect 33376 14424 33382 14476
rect 34514 14424 34520 14476
rect 34572 14464 34578 14476
rect 35069 14467 35127 14473
rect 35069 14464 35081 14467
rect 34572 14436 35081 14464
rect 34572 14424 34578 14436
rect 35069 14433 35081 14436
rect 35115 14433 35127 14467
rect 35434 14464 35440 14476
rect 35395 14436 35440 14464
rect 35069 14427 35127 14433
rect 35434 14424 35440 14436
rect 35492 14424 35498 14476
rect 25409 14399 25467 14405
rect 25409 14365 25421 14399
rect 25455 14365 25467 14399
rect 25409 14359 25467 14365
rect 25593 14399 25651 14405
rect 25593 14365 25605 14399
rect 25639 14396 25651 14399
rect 25774 14396 25780 14408
rect 25639 14368 25780 14396
rect 25639 14365 25651 14368
rect 25593 14359 25651 14365
rect 21729 14331 21787 14337
rect 17736 14300 20024 14328
rect 17736 14288 17742 14300
rect 19996 14272 20024 14300
rect 21729 14297 21741 14331
rect 21775 14328 21787 14331
rect 23106 14328 23112 14340
rect 21775 14300 23112 14328
rect 21775 14297 21787 14300
rect 21729 14291 21787 14297
rect 23106 14288 23112 14300
rect 23164 14288 23170 14340
rect 23198 14288 23204 14340
rect 23256 14328 23262 14340
rect 23937 14331 23995 14337
rect 23937 14328 23949 14331
rect 23256 14300 23949 14328
rect 23256 14288 23262 14300
rect 23937 14297 23949 14300
rect 23983 14328 23995 14331
rect 25608 14328 25636 14359
rect 25774 14356 25780 14368
rect 25832 14356 25838 14408
rect 27709 14399 27767 14405
rect 27709 14365 27721 14399
rect 27755 14396 27767 14399
rect 27798 14396 27804 14408
rect 27755 14368 27804 14396
rect 27755 14365 27767 14368
rect 27709 14359 27767 14365
rect 27798 14356 27804 14368
rect 27856 14396 27862 14408
rect 28350 14396 28356 14408
rect 27856 14368 28356 14396
rect 27856 14356 27862 14368
rect 28350 14356 28356 14368
rect 28408 14356 28414 14408
rect 28813 14399 28871 14405
rect 28813 14365 28825 14399
rect 28859 14365 28871 14399
rect 29914 14396 29920 14408
rect 29875 14368 29920 14396
rect 28813 14359 28871 14365
rect 23983 14300 25636 14328
rect 23983 14297 23995 14300
rect 23937 14291 23995 14297
rect 27246 14288 27252 14340
rect 27304 14328 27310 14340
rect 28828 14328 28856 14359
rect 29914 14356 29920 14368
rect 29972 14356 29978 14408
rect 33229 14399 33287 14405
rect 33229 14365 33241 14399
rect 33275 14396 33287 14399
rect 33410 14396 33416 14408
rect 33275 14368 33416 14396
rect 33275 14365 33287 14368
rect 33229 14359 33287 14365
rect 33410 14356 33416 14368
rect 33468 14356 33474 14408
rect 35158 14356 35164 14408
rect 35216 14396 35222 14408
rect 35216 14368 35261 14396
rect 35216 14356 35222 14368
rect 35710 14356 35716 14408
rect 35768 14396 35774 14408
rect 37182 14405 37188 14408
rect 36909 14399 36967 14405
rect 36909 14396 36921 14399
rect 35768 14368 36921 14396
rect 35768 14356 35774 14368
rect 36909 14365 36921 14368
rect 36955 14365 36967 14399
rect 37176 14396 37188 14405
rect 37143 14368 37188 14396
rect 36909 14359 36967 14365
rect 37176 14359 37188 14368
rect 37182 14356 37188 14359
rect 37240 14356 37246 14408
rect 27304 14300 28856 14328
rect 27304 14288 27310 14300
rect 32674 14288 32680 14340
rect 32732 14328 32738 14340
rect 33502 14328 33508 14340
rect 32732 14300 33508 14328
rect 32732 14288 32738 14300
rect 33502 14288 33508 14300
rect 33560 14328 33566 14340
rect 35529 14331 35587 14337
rect 33560 14300 34836 14328
rect 33560 14288 33566 14300
rect 17034 14220 17040 14272
rect 17092 14260 17098 14272
rect 18785 14263 18843 14269
rect 18785 14260 18797 14263
rect 17092 14232 18797 14260
rect 17092 14220 17098 14232
rect 18785 14229 18797 14232
rect 18831 14260 18843 14263
rect 18874 14260 18880 14272
rect 18831 14232 18880 14260
rect 18831 14229 18843 14232
rect 18785 14223 18843 14229
rect 18874 14220 18880 14232
rect 18932 14220 18938 14272
rect 19334 14220 19340 14272
rect 19392 14260 19398 14272
rect 19889 14263 19947 14269
rect 19889 14260 19901 14263
rect 19392 14232 19901 14260
rect 19392 14220 19398 14232
rect 19889 14229 19901 14232
rect 19935 14229 19947 14263
rect 19889 14223 19947 14229
rect 19978 14220 19984 14272
rect 20036 14260 20042 14272
rect 20036 14232 20081 14260
rect 20036 14220 20042 14232
rect 20346 14220 20352 14272
rect 20404 14260 20410 14272
rect 22554 14260 22560 14272
rect 20404 14232 22560 14260
rect 20404 14220 20410 14232
rect 22554 14220 22560 14232
rect 22612 14220 22618 14272
rect 23385 14263 23443 14269
rect 23385 14229 23397 14263
rect 23431 14260 23443 14263
rect 23842 14260 23848 14272
rect 23431 14232 23848 14260
rect 23431 14229 23443 14232
rect 23385 14223 23443 14229
rect 23842 14220 23848 14232
rect 23900 14220 23906 14272
rect 24210 14220 24216 14272
rect 24268 14260 24274 14272
rect 24949 14263 25007 14269
rect 24949 14260 24961 14263
rect 24268 14232 24961 14260
rect 24268 14220 24274 14232
rect 24949 14229 24961 14232
rect 24995 14229 25007 14263
rect 24949 14223 25007 14229
rect 25038 14220 25044 14272
rect 25096 14260 25102 14272
rect 28994 14260 29000 14272
rect 25096 14232 29000 14260
rect 25096 14220 25102 14232
rect 28994 14220 29000 14232
rect 29052 14220 29058 14272
rect 30285 14263 30343 14269
rect 30285 14229 30297 14263
rect 30331 14260 30343 14263
rect 30834 14260 30840 14272
rect 30331 14232 30840 14260
rect 30331 14229 30343 14232
rect 30285 14223 30343 14229
rect 30834 14220 30840 14232
rect 30892 14220 30898 14272
rect 33597 14263 33655 14269
rect 33597 14229 33609 14263
rect 33643 14260 33655 14263
rect 34698 14260 34704 14272
rect 33643 14232 34704 14260
rect 33643 14229 33655 14232
rect 33597 14223 33655 14229
rect 34698 14220 34704 14232
rect 34756 14220 34762 14272
rect 34808 14260 34836 14300
rect 35529 14297 35541 14331
rect 35575 14328 35587 14331
rect 36446 14328 36452 14340
rect 35575 14300 36452 14328
rect 35575 14297 35587 14300
rect 35529 14291 35587 14297
rect 35544 14260 35572 14291
rect 36446 14288 36452 14300
rect 36504 14288 36510 14340
rect 34808 14232 35572 14260
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 9306 14056 9312 14068
rect 9267 14028 9312 14056
rect 9306 14016 9312 14028
rect 9364 14016 9370 14068
rect 17497 14059 17555 14065
rect 17497 14025 17509 14059
rect 17543 14056 17555 14059
rect 17862 14056 17868 14068
rect 17543 14028 17868 14056
rect 17543 14025 17555 14028
rect 17497 14019 17555 14025
rect 17862 14016 17868 14028
rect 17920 14016 17926 14068
rect 19426 14016 19432 14068
rect 19484 14056 19490 14068
rect 19889 14059 19947 14065
rect 19889 14056 19901 14059
rect 19484 14028 19901 14056
rect 19484 14016 19490 14028
rect 19889 14025 19901 14028
rect 19935 14025 19947 14059
rect 22738 14056 22744 14068
rect 22699 14028 22744 14056
rect 19889 14019 19947 14025
rect 22738 14016 22744 14028
rect 22796 14016 22802 14068
rect 24397 14059 24455 14065
rect 24397 14025 24409 14059
rect 24443 14056 24455 14059
rect 29914 14056 29920 14068
rect 24443 14028 29920 14056
rect 24443 14025 24455 14028
rect 24397 14019 24455 14025
rect 29914 14016 29920 14028
rect 29972 14016 29978 14068
rect 31662 14016 31668 14068
rect 31720 14056 31726 14068
rect 31757 14059 31815 14065
rect 31757 14056 31769 14059
rect 31720 14028 31769 14056
rect 31720 14016 31726 14028
rect 31757 14025 31769 14028
rect 31803 14025 31815 14059
rect 32766 14056 32772 14068
rect 32727 14028 32772 14056
rect 31757 14019 31815 14025
rect 32766 14016 32772 14028
rect 32824 14016 32830 14068
rect 35253 14059 35311 14065
rect 33336 14028 33732 14056
rect 8196 13991 8254 13997
rect 8196 13957 8208 13991
rect 8242 13988 8254 13991
rect 8386 13988 8392 14000
rect 8242 13960 8392 13988
rect 8242 13957 8254 13960
rect 8196 13951 8254 13957
rect 8386 13948 8392 13960
rect 8444 13948 8450 14000
rect 9324 13988 9352 14016
rect 12066 13988 12072 14000
rect 9324 13960 12072 13988
rect 7926 13920 7932 13932
rect 7887 13892 7932 13920
rect 7926 13880 7932 13892
rect 7984 13880 7990 13932
rect 10594 13920 10600 13932
rect 10555 13892 10600 13920
rect 10594 13880 10600 13892
rect 10652 13880 10658 13932
rect 11716 13929 11744 13960
rect 12066 13948 12072 13960
rect 12124 13948 12130 14000
rect 13630 13988 13636 14000
rect 12912 13960 13636 13988
rect 11701 13923 11759 13929
rect 11701 13889 11713 13923
rect 11747 13889 11759 13923
rect 11882 13920 11888 13932
rect 11843 13892 11888 13920
rect 11701 13883 11759 13889
rect 11882 13880 11888 13892
rect 11940 13880 11946 13932
rect 12912 13929 12940 13960
rect 13630 13948 13636 13960
rect 13688 13988 13694 14000
rect 16853 13991 16911 13997
rect 13688 13960 14596 13988
rect 13688 13948 13694 13960
rect 12897 13923 12955 13929
rect 12897 13889 12909 13923
rect 12943 13889 12955 13923
rect 12897 13883 12955 13889
rect 12986 13880 12992 13932
rect 13044 13920 13050 13932
rect 13044 13892 13089 13920
rect 13044 13880 13050 13892
rect 13262 13880 13268 13932
rect 13320 13920 13326 13932
rect 13357 13923 13415 13929
rect 13357 13920 13369 13923
rect 13320 13892 13369 13920
rect 13320 13880 13326 13892
rect 13357 13889 13369 13892
rect 13403 13889 13415 13923
rect 13357 13883 13415 13889
rect 13538 13880 13544 13932
rect 13596 13920 13602 13932
rect 14369 13923 14427 13929
rect 14369 13920 14381 13923
rect 13596 13892 14381 13920
rect 13596 13880 13602 13892
rect 14369 13889 14381 13892
rect 14415 13889 14427 13923
rect 14369 13883 14427 13889
rect 10686 13852 10692 13864
rect 10647 13824 10692 13852
rect 10686 13812 10692 13824
rect 10744 13812 10750 13864
rect 12069 13855 12127 13861
rect 12069 13821 12081 13855
rect 12115 13852 12127 13855
rect 12710 13852 12716 13864
rect 12115 13824 12716 13852
rect 12115 13821 12127 13824
rect 12069 13815 12127 13821
rect 12710 13812 12716 13824
rect 12768 13812 12774 13864
rect 13081 13855 13139 13861
rect 13081 13821 13093 13855
rect 13127 13852 13139 13855
rect 13170 13852 13176 13864
rect 13127 13824 13176 13852
rect 13127 13821 13139 13824
rect 13081 13815 13139 13821
rect 13170 13812 13176 13824
rect 13228 13812 13234 13864
rect 14568 13852 14596 13960
rect 16853 13957 16865 13991
rect 16899 13988 16911 13991
rect 17954 13988 17960 14000
rect 16899 13960 17960 13988
rect 16899 13957 16911 13960
rect 16853 13951 16911 13957
rect 17954 13948 17960 13960
rect 18012 13948 18018 14000
rect 18690 13948 18696 14000
rect 18748 13988 18754 14000
rect 19245 13991 19303 13997
rect 19245 13988 19257 13991
rect 18748 13960 19257 13988
rect 18748 13948 18754 13960
rect 19245 13957 19257 13960
rect 19291 13988 19303 13991
rect 20254 13988 20260 14000
rect 19291 13960 20260 13988
rect 19291 13957 19303 13960
rect 19245 13951 19303 13957
rect 20254 13948 20260 13960
rect 20312 13948 20318 14000
rect 23753 13991 23811 13997
rect 23753 13988 23765 13991
rect 22940 13960 23765 13988
rect 14829 13923 14887 13929
rect 14829 13889 14841 13923
rect 14875 13920 14887 13923
rect 15010 13920 15016 13932
rect 14875 13892 15016 13920
rect 14875 13889 14887 13892
rect 14829 13883 14887 13889
rect 15010 13880 15016 13892
rect 15068 13880 15074 13932
rect 15378 13920 15384 13932
rect 15339 13892 15384 13920
rect 15378 13880 15384 13892
rect 15436 13880 15442 13932
rect 17218 13920 17224 13932
rect 17179 13892 17224 13920
rect 17218 13880 17224 13892
rect 17276 13920 17282 13932
rect 19334 13920 19340 13932
rect 17276 13892 19340 13920
rect 17276 13880 17282 13892
rect 19334 13880 19340 13892
rect 19392 13920 19398 13932
rect 19613 13923 19671 13929
rect 19613 13920 19625 13923
rect 19392 13892 19625 13920
rect 19392 13880 19398 13892
rect 19613 13889 19625 13892
rect 19659 13889 19671 13923
rect 19613 13883 19671 13889
rect 19705 13923 19763 13929
rect 19705 13889 19717 13923
rect 19751 13920 19763 13923
rect 20070 13920 20076 13932
rect 19751 13892 20076 13920
rect 19751 13889 19763 13892
rect 19705 13883 19763 13889
rect 20070 13880 20076 13892
rect 20128 13920 20134 13932
rect 20346 13920 20352 13932
rect 20128 13892 20352 13920
rect 20128 13880 20134 13892
rect 20346 13880 20352 13892
rect 20404 13880 20410 13932
rect 22940 13929 22968 13960
rect 23753 13957 23765 13960
rect 23799 13988 23811 13991
rect 23934 13988 23940 14000
rect 23799 13960 23940 13988
rect 23799 13957 23811 13960
rect 23753 13951 23811 13957
rect 23934 13948 23940 13960
rect 23992 13988 23998 14000
rect 24949 13991 25007 13997
rect 24949 13988 24961 13991
rect 23992 13960 24961 13988
rect 23992 13948 23998 13960
rect 24949 13957 24961 13960
rect 24995 13957 25007 13991
rect 27154 13988 27160 14000
rect 27115 13960 27160 13988
rect 24949 13951 25007 13957
rect 27154 13948 27160 13960
rect 27212 13948 27218 14000
rect 27246 13948 27252 14000
rect 27304 13988 27310 14000
rect 27341 13991 27399 13997
rect 27341 13988 27353 13991
rect 27304 13960 27353 13988
rect 27304 13948 27310 13960
rect 27341 13957 27353 13960
rect 27387 13957 27399 13991
rect 33336 13988 33364 14028
rect 27341 13951 27399 13957
rect 30392 13960 33364 13988
rect 33413 13991 33471 13997
rect 22925 13923 22983 13929
rect 22925 13889 22937 13923
rect 22971 13889 22983 13923
rect 23198 13920 23204 13932
rect 23159 13892 23204 13920
rect 22925 13883 22983 13889
rect 23198 13880 23204 13892
rect 23256 13880 23262 13932
rect 24210 13920 24216 13932
rect 24171 13892 24216 13920
rect 24210 13880 24216 13892
rect 24268 13880 24274 13932
rect 24578 13880 24584 13932
rect 24636 13920 24642 13932
rect 24857 13923 24915 13929
rect 24857 13920 24869 13923
rect 24636 13892 24869 13920
rect 24636 13880 24642 13892
rect 24857 13889 24869 13892
rect 24903 13889 24915 13923
rect 25038 13920 25044 13932
rect 24999 13892 25044 13920
rect 24857 13883 24915 13889
rect 25038 13880 25044 13892
rect 25096 13880 25102 13932
rect 25866 13880 25872 13932
rect 25924 13920 25930 13932
rect 26053 13923 26111 13929
rect 26053 13920 26065 13923
rect 25924 13892 26065 13920
rect 25924 13880 25930 13892
rect 26053 13889 26065 13892
rect 26099 13889 26111 13923
rect 26326 13920 26332 13932
rect 26239 13892 26332 13920
rect 26053 13883 26111 13889
rect 26326 13880 26332 13892
rect 26384 13920 26390 13932
rect 26970 13920 26976 13932
rect 26384 13892 26976 13920
rect 26384 13880 26390 13892
rect 26970 13880 26976 13892
rect 27028 13880 27034 13932
rect 27433 13923 27491 13929
rect 27433 13889 27445 13923
rect 27479 13889 27491 13923
rect 27982 13920 27988 13932
rect 27943 13892 27988 13920
rect 27433 13883 27491 13889
rect 15194 13852 15200 13864
rect 14568 13824 15056 13852
rect 15155 13824 15200 13852
rect 10965 13787 11023 13793
rect 10965 13753 10977 13787
rect 11011 13784 11023 13787
rect 13722 13784 13728 13796
rect 11011 13756 13728 13784
rect 11011 13753 11023 13756
rect 10965 13747 11023 13753
rect 13722 13744 13728 13756
rect 13780 13744 13786 13796
rect 15028 13793 15056 13824
rect 15194 13812 15200 13824
rect 15252 13812 15258 13864
rect 17313 13855 17371 13861
rect 17313 13821 17325 13855
rect 17359 13852 17371 13855
rect 17402 13852 17408 13864
rect 17359 13824 17408 13852
rect 17359 13821 17371 13824
rect 17313 13815 17371 13821
rect 17402 13812 17408 13824
rect 17460 13852 17466 13864
rect 18322 13852 18328 13864
rect 17460 13824 18328 13852
rect 17460 13812 17466 13824
rect 18322 13812 18328 13824
rect 18380 13812 18386 13864
rect 22738 13812 22744 13864
rect 22796 13852 22802 13864
rect 23017 13855 23075 13861
rect 23017 13852 23029 13855
rect 22796 13824 23029 13852
rect 22796 13812 22802 13824
rect 23017 13821 23029 13824
rect 23063 13821 23075 13855
rect 23017 13815 23075 13821
rect 23109 13855 23167 13861
rect 23109 13821 23121 13855
rect 23155 13852 23167 13855
rect 23474 13852 23480 13864
rect 23155 13824 23480 13852
rect 23155 13821 23167 13824
rect 23109 13815 23167 13821
rect 23474 13812 23480 13824
rect 23532 13852 23538 13864
rect 24118 13852 24124 13864
rect 23532 13824 24124 13852
rect 23532 13812 23538 13824
rect 24118 13812 24124 13824
rect 24176 13812 24182 13864
rect 25501 13855 25559 13861
rect 25501 13821 25513 13855
rect 25547 13821 25559 13855
rect 25501 13815 25559 13821
rect 26513 13855 26571 13861
rect 26513 13821 26525 13855
rect 26559 13821 26571 13855
rect 27448 13852 27476 13883
rect 27982 13880 27988 13892
rect 28040 13880 28046 13932
rect 28810 13920 28816 13932
rect 28771 13892 28816 13920
rect 28810 13880 28816 13892
rect 28868 13880 28874 13932
rect 30392 13864 30420 13960
rect 33413 13957 33425 13991
rect 33459 13988 33471 13991
rect 33502 13988 33508 14000
rect 33459 13960 33508 13988
rect 33459 13957 33471 13960
rect 33413 13951 33471 13957
rect 33502 13948 33508 13960
rect 33560 13948 33566 14000
rect 30644 13923 30702 13929
rect 30644 13889 30656 13923
rect 30690 13920 30702 13923
rect 31110 13920 31116 13932
rect 30690 13892 31116 13920
rect 30690 13889 30702 13892
rect 30644 13883 30702 13889
rect 31110 13880 31116 13892
rect 31168 13880 31174 13932
rect 31202 13880 31208 13932
rect 31260 13920 31266 13932
rect 33042 13920 33048 13932
rect 31260 13892 33048 13920
rect 31260 13880 31266 13892
rect 33042 13880 33048 13892
rect 33100 13880 33106 13932
rect 27614 13852 27620 13864
rect 27448 13824 27620 13852
rect 26513 13815 26571 13821
rect 13817 13787 13875 13793
rect 13817 13753 13829 13787
rect 13863 13753 13875 13787
rect 13817 13747 13875 13753
rect 15013 13787 15071 13793
rect 15013 13753 15025 13787
rect 15059 13753 15071 13787
rect 15013 13747 15071 13753
rect 13832 13716 13860 13747
rect 15102 13744 15108 13796
rect 15160 13784 15166 13796
rect 21358 13784 21364 13796
rect 15160 13756 21364 13784
rect 15160 13744 15166 13756
rect 21358 13744 21364 13756
rect 21416 13744 21422 13796
rect 25516 13784 25544 13815
rect 22066 13756 25544 13784
rect 26528 13784 26556 13815
rect 27614 13812 27620 13824
rect 27672 13852 27678 13864
rect 28626 13852 28632 13864
rect 27672 13824 28632 13852
rect 27672 13812 27678 13824
rect 28626 13812 28632 13824
rect 28684 13812 28690 13864
rect 30374 13852 30380 13864
rect 30335 13824 30380 13852
rect 30374 13812 30380 13824
rect 30432 13812 30438 13864
rect 32858 13812 32864 13864
rect 32916 13852 32922 13864
rect 32953 13855 33011 13861
rect 32953 13852 32965 13855
rect 32916 13824 32965 13852
rect 32916 13812 32922 13824
rect 32953 13821 32965 13824
rect 32999 13821 33011 13855
rect 33318 13852 33324 13864
rect 33279 13824 33324 13852
rect 32953 13815 33011 13821
rect 33318 13812 33324 13824
rect 33376 13812 33382 13864
rect 33704 13852 33732 14028
rect 35253 14025 35265 14059
rect 35299 14056 35311 14059
rect 35526 14056 35532 14068
rect 35299 14028 35532 14056
rect 35299 14025 35311 14028
rect 35253 14019 35311 14025
rect 35526 14016 35532 14028
rect 35584 14016 35590 14068
rect 34790 13988 34796 14000
rect 33888 13960 34796 13988
rect 33888 13929 33916 13960
rect 34790 13948 34796 13960
rect 34848 13988 34854 14000
rect 35710 13988 35716 14000
rect 34848 13960 35716 13988
rect 34848 13948 34854 13960
rect 35710 13948 35716 13960
rect 35768 13948 35774 14000
rect 36446 13988 36452 14000
rect 36407 13960 36452 13988
rect 36446 13948 36452 13960
rect 36504 13948 36510 14000
rect 33873 13923 33931 13929
rect 33873 13889 33885 13923
rect 33919 13889 33931 13923
rect 33873 13883 33931 13889
rect 33888 13852 33916 13883
rect 33962 13880 33968 13932
rect 34020 13920 34026 13932
rect 34129 13923 34187 13929
rect 34129 13920 34141 13923
rect 34020 13892 34141 13920
rect 34020 13880 34026 13892
rect 34129 13889 34141 13892
rect 34175 13889 34187 13923
rect 34129 13883 34187 13889
rect 35158 13880 35164 13932
rect 35216 13920 35222 13932
rect 36081 13923 36139 13929
rect 36081 13920 36093 13923
rect 35216 13892 36093 13920
rect 35216 13880 35222 13892
rect 36081 13889 36093 13892
rect 36127 13889 36139 13923
rect 36081 13883 36139 13889
rect 36170 13880 36176 13932
rect 36228 13920 36234 13932
rect 36357 13923 36415 13929
rect 36357 13920 36369 13923
rect 36228 13892 36369 13920
rect 36228 13880 36234 13892
rect 36357 13889 36369 13892
rect 36403 13889 36415 13923
rect 36357 13883 36415 13889
rect 33704 13824 33916 13852
rect 35342 13812 35348 13864
rect 35400 13852 35406 13864
rect 35618 13852 35624 13864
rect 35400 13824 35624 13852
rect 35400 13812 35406 13824
rect 35618 13812 35624 13824
rect 35676 13852 35682 13864
rect 35989 13855 36047 13861
rect 35989 13852 36001 13855
rect 35676 13824 36001 13852
rect 35676 13812 35682 13824
rect 35989 13821 36001 13824
rect 36035 13821 36047 13855
rect 38286 13852 38292 13864
rect 38247 13824 38292 13852
rect 35989 13815 36047 13821
rect 38286 13812 38292 13824
rect 38344 13812 38350 13864
rect 27798 13784 27804 13796
rect 26528 13756 27804 13784
rect 16022 13716 16028 13728
rect 13832 13688 16028 13716
rect 16022 13676 16028 13688
rect 16080 13676 16086 13728
rect 18138 13676 18144 13728
rect 18196 13716 18202 13728
rect 22066 13716 22094 13756
rect 27798 13744 27804 13756
rect 27856 13744 27862 13796
rect 35802 13784 35808 13796
rect 35763 13756 35808 13784
rect 35802 13744 35808 13756
rect 35860 13744 35866 13796
rect 18196 13688 22094 13716
rect 18196 13676 18202 13688
rect 22830 13676 22836 13728
rect 22888 13716 22894 13728
rect 23382 13716 23388 13728
rect 22888 13688 23388 13716
rect 22888 13676 22894 13688
rect 23382 13676 23388 13688
rect 23440 13716 23446 13728
rect 25038 13716 25044 13728
rect 23440 13688 25044 13716
rect 23440 13676 23446 13688
rect 25038 13676 25044 13688
rect 25096 13676 25102 13728
rect 26970 13676 26976 13728
rect 27028 13716 27034 13728
rect 27157 13719 27215 13725
rect 27157 13716 27169 13719
rect 27028 13688 27169 13716
rect 27028 13676 27034 13688
rect 27157 13685 27169 13688
rect 27203 13685 27215 13719
rect 28166 13716 28172 13728
rect 28127 13688 28172 13716
rect 27157 13679 27215 13685
rect 28166 13676 28172 13688
rect 28224 13676 28230 13728
rect 29178 13676 29184 13728
rect 29236 13716 29242 13728
rect 29273 13719 29331 13725
rect 29273 13716 29285 13719
rect 29236 13688 29285 13716
rect 29236 13676 29242 13688
rect 29273 13685 29285 13688
rect 29319 13685 29331 13719
rect 29273 13679 29331 13685
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 10686 13512 10692 13524
rect 10647 13484 10692 13512
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 10778 13472 10784 13524
rect 10836 13512 10842 13524
rect 15102 13512 15108 13524
rect 10836 13484 15108 13512
rect 10836 13472 10842 13484
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 15194 13472 15200 13524
rect 15252 13512 15258 13524
rect 15841 13515 15899 13521
rect 15841 13512 15853 13515
rect 15252 13484 15853 13512
rect 15252 13472 15258 13484
rect 15841 13481 15853 13484
rect 15887 13481 15899 13515
rect 23566 13512 23572 13524
rect 23527 13484 23572 13512
rect 15841 13475 15899 13481
rect 23566 13472 23572 13484
rect 23624 13472 23630 13524
rect 30190 13512 30196 13524
rect 23676 13484 30196 13512
rect 15212 13444 15240 13472
rect 18138 13444 18144 13456
rect 14292 13416 15240 13444
rect 16224 13416 18144 13444
rect 10505 13379 10563 13385
rect 10505 13345 10517 13379
rect 10551 13376 10563 13379
rect 11146 13376 11152 13388
rect 10551 13348 11152 13376
rect 10551 13345 10563 13348
rect 10505 13339 10563 13345
rect 11146 13336 11152 13348
rect 11204 13336 11210 13388
rect 14292 13385 14320 13416
rect 14277 13379 14335 13385
rect 14277 13345 14289 13379
rect 14323 13345 14335 13379
rect 15378 13376 15384 13388
rect 14277 13339 14335 13345
rect 14476 13348 15384 13376
rect 10413 13311 10471 13317
rect 10413 13277 10425 13311
rect 10459 13308 10471 13311
rect 10778 13308 10784 13320
rect 10459 13280 10784 13308
rect 10459 13277 10471 13280
rect 10413 13271 10471 13277
rect 10778 13268 10784 13280
rect 10836 13268 10842 13320
rect 12161 13311 12219 13317
rect 12161 13277 12173 13311
rect 12207 13308 12219 13311
rect 12434 13308 12440 13320
rect 12207 13280 12440 13308
rect 12207 13277 12219 13280
rect 12161 13271 12219 13277
rect 12434 13268 12440 13280
rect 12492 13268 12498 13320
rect 14476 13317 14504 13348
rect 15378 13336 15384 13348
rect 15436 13336 15442 13388
rect 14461 13311 14519 13317
rect 14461 13277 14473 13311
rect 14507 13277 14519 13311
rect 14461 13271 14519 13277
rect 14829 13311 14887 13317
rect 14829 13277 14841 13311
rect 14875 13308 14887 13311
rect 15010 13308 15016 13320
rect 14875 13280 15016 13308
rect 14875 13277 14887 13280
rect 14829 13271 14887 13277
rect 15010 13268 15016 13280
rect 15068 13268 15074 13320
rect 15746 13268 15752 13320
rect 15804 13308 15810 13320
rect 16224 13317 16252 13416
rect 18138 13404 18144 13416
rect 18196 13404 18202 13456
rect 23290 13404 23296 13456
rect 23348 13444 23354 13456
rect 23676 13444 23704 13484
rect 30190 13472 30196 13484
rect 30248 13472 30254 13524
rect 36722 13472 36728 13524
rect 36780 13512 36786 13524
rect 37093 13515 37151 13521
rect 37093 13512 37105 13515
rect 36780 13484 37105 13512
rect 36780 13472 36786 13484
rect 37093 13481 37105 13484
rect 37139 13481 37151 13515
rect 37093 13475 37151 13481
rect 23348 13416 23704 13444
rect 23348 13404 23354 13416
rect 25590 13404 25596 13456
rect 25648 13444 25654 13456
rect 25869 13447 25927 13453
rect 25869 13444 25881 13447
rect 25648 13416 25881 13444
rect 25648 13404 25654 13416
rect 25869 13413 25881 13416
rect 25915 13413 25927 13447
rect 25869 13407 25927 13413
rect 27157 13447 27215 13453
rect 27157 13413 27169 13447
rect 27203 13444 27215 13447
rect 28810 13444 28816 13456
rect 27203 13416 28816 13444
rect 27203 13413 27215 13416
rect 27157 13407 27215 13413
rect 28810 13404 28816 13416
rect 28868 13404 28874 13456
rect 30926 13404 30932 13456
rect 30984 13444 30990 13456
rect 33778 13444 33784 13456
rect 30984 13416 33784 13444
rect 30984 13404 30990 13416
rect 33778 13404 33784 13416
rect 33836 13404 33842 13456
rect 17586 13376 17592 13388
rect 16500 13348 17592 13376
rect 16500 13320 16528 13348
rect 17586 13336 17592 13348
rect 17644 13376 17650 13388
rect 19978 13376 19984 13388
rect 17644 13348 17908 13376
rect 17644 13336 17650 13348
rect 16209 13311 16267 13317
rect 16209 13308 16221 13311
rect 15804 13280 16221 13308
rect 15804 13268 15810 13280
rect 16209 13277 16221 13280
rect 16255 13277 16267 13311
rect 16482 13308 16488 13320
rect 16395 13280 16488 13308
rect 16209 13271 16267 13277
rect 16482 13268 16488 13280
rect 16540 13268 16546 13320
rect 16577 13311 16635 13317
rect 16577 13277 16589 13311
rect 16623 13308 16635 13311
rect 16850 13308 16856 13320
rect 16623 13280 16712 13308
rect 16811 13280 16856 13308
rect 16623 13277 16635 13280
rect 16577 13271 16635 13277
rect 12894 13240 12900 13252
rect 12855 13212 12900 13240
rect 12894 13200 12900 13212
rect 12952 13200 12958 13252
rect 13262 13132 13268 13184
rect 13320 13172 13326 13184
rect 14461 13175 14519 13181
rect 14461 13172 14473 13175
rect 13320 13144 14473 13172
rect 13320 13132 13326 13144
rect 14461 13141 14473 13144
rect 14507 13141 14519 13175
rect 14461 13135 14519 13141
rect 14550 13132 14556 13184
rect 14608 13172 14614 13184
rect 16684 13172 16712 13280
rect 16850 13268 16856 13280
rect 16908 13268 16914 13320
rect 17880 13317 17908 13348
rect 17972 13348 19984 13376
rect 17972 13317 18000 13348
rect 19978 13336 19984 13348
rect 20036 13376 20042 13388
rect 20036 13348 21128 13376
rect 20036 13336 20042 13348
rect 17129 13311 17187 13317
rect 17129 13277 17141 13311
rect 17175 13308 17187 13311
rect 17681 13311 17739 13317
rect 17681 13308 17693 13311
rect 17175 13280 17693 13308
rect 17175 13277 17187 13280
rect 17129 13271 17187 13277
rect 17681 13277 17693 13280
rect 17727 13277 17739 13311
rect 17681 13271 17739 13277
rect 17865 13311 17923 13317
rect 17865 13277 17877 13311
rect 17911 13277 17923 13311
rect 17865 13271 17923 13277
rect 17957 13311 18015 13317
rect 17957 13277 17969 13311
rect 18003 13277 18015 13311
rect 18138 13308 18144 13320
rect 18099 13280 18144 13308
rect 17957 13271 18015 13277
rect 18138 13268 18144 13280
rect 18196 13268 18202 13320
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13277 18291 13311
rect 20898 13308 20904 13320
rect 20859 13280 20904 13308
rect 18233 13271 18291 13277
rect 17770 13200 17776 13252
rect 17828 13240 17834 13252
rect 18248 13240 18276 13271
rect 20898 13268 20904 13280
rect 20956 13268 20962 13320
rect 21100 13317 21128 13348
rect 21726 13336 21732 13388
rect 21784 13376 21790 13388
rect 21821 13379 21879 13385
rect 21821 13376 21833 13379
rect 21784 13348 21833 13376
rect 21784 13336 21790 13348
rect 21821 13345 21833 13348
rect 21867 13345 21879 13379
rect 26970 13376 26976 13388
rect 26931 13348 26976 13376
rect 21821 13339 21879 13345
rect 26970 13336 26976 13348
rect 27028 13336 27034 13388
rect 27614 13376 27620 13388
rect 27172 13348 27620 13376
rect 21085 13311 21143 13317
rect 21085 13277 21097 13311
rect 21131 13277 21143 13311
rect 21542 13308 21548 13320
rect 21503 13280 21548 13308
rect 21085 13271 21143 13277
rect 21542 13268 21548 13280
rect 21600 13268 21606 13320
rect 21634 13268 21640 13320
rect 21692 13308 21698 13320
rect 21692 13280 21737 13308
rect 21692 13268 21698 13280
rect 23474 13268 23480 13320
rect 23532 13308 23538 13320
rect 23569 13311 23627 13317
rect 23569 13308 23581 13311
rect 23532 13280 23581 13308
rect 23532 13268 23538 13280
rect 23569 13277 23581 13280
rect 23615 13277 23627 13311
rect 23569 13271 23627 13277
rect 23845 13311 23903 13317
rect 23845 13277 23857 13311
rect 23891 13308 23903 13311
rect 23934 13308 23940 13320
rect 23891 13280 23940 13308
rect 23891 13277 23903 13280
rect 23845 13271 23903 13277
rect 23934 13268 23940 13280
rect 23992 13268 23998 13320
rect 25866 13308 25872 13320
rect 25827 13280 25872 13308
rect 25866 13268 25872 13280
rect 25924 13268 25930 13320
rect 26145 13311 26203 13317
rect 26145 13277 26157 13311
rect 26191 13308 26203 13311
rect 27172 13308 27200 13348
rect 27614 13336 27620 13348
rect 27672 13336 27678 13388
rect 28445 13379 28503 13385
rect 28445 13345 28457 13379
rect 28491 13376 28503 13379
rect 28994 13376 29000 13388
rect 28491 13348 29000 13376
rect 28491 13345 28503 13348
rect 28445 13339 28503 13345
rect 28994 13336 29000 13348
rect 29052 13336 29058 13388
rect 30834 13376 30840 13388
rect 30795 13348 30840 13376
rect 30834 13336 30840 13348
rect 30892 13336 30898 13388
rect 35710 13376 35716 13388
rect 35671 13348 35716 13376
rect 35710 13336 35716 13348
rect 35768 13336 35774 13388
rect 26191 13280 27200 13308
rect 27249 13311 27307 13317
rect 26191 13277 26203 13280
rect 26145 13271 26203 13277
rect 27249 13277 27261 13311
rect 27295 13308 27307 13311
rect 27798 13308 27804 13320
rect 27295 13280 27804 13308
rect 27295 13277 27307 13280
rect 27249 13271 27307 13277
rect 27798 13268 27804 13280
rect 27856 13268 27862 13320
rect 28350 13308 28356 13320
rect 28311 13280 28356 13308
rect 28350 13268 28356 13280
rect 28408 13268 28414 13320
rect 28721 13311 28779 13317
rect 28721 13308 28733 13311
rect 28460 13280 28733 13308
rect 17828 13212 18276 13240
rect 20916 13240 20944 13268
rect 21910 13240 21916 13252
rect 20916 13212 21916 13240
rect 17828 13200 17834 13212
rect 21910 13200 21916 13212
rect 21968 13200 21974 13252
rect 22738 13200 22744 13252
rect 22796 13240 22802 13252
rect 23753 13243 23811 13249
rect 23753 13240 23765 13243
rect 22796 13212 23765 13240
rect 22796 13200 22802 13212
rect 23753 13209 23765 13212
rect 23799 13240 23811 13243
rect 24210 13240 24216 13252
rect 23799 13212 24216 13240
rect 23799 13209 23811 13212
rect 23753 13203 23811 13209
rect 24210 13200 24216 13212
rect 24268 13200 24274 13252
rect 25038 13200 25044 13252
rect 25096 13240 25102 13252
rect 26053 13243 26111 13249
rect 26053 13240 26065 13243
rect 25096 13212 26065 13240
rect 25096 13200 25102 13212
rect 26053 13209 26065 13212
rect 26099 13209 26111 13243
rect 26053 13203 26111 13209
rect 27614 13200 27620 13252
rect 27672 13240 27678 13252
rect 27709 13243 27767 13249
rect 27709 13240 27721 13243
rect 27672 13212 27721 13240
rect 27672 13200 27678 13212
rect 27709 13209 27721 13212
rect 27755 13209 27767 13243
rect 27709 13203 27767 13209
rect 28258 13200 28264 13252
rect 28316 13240 28322 13252
rect 28460 13240 28488 13280
rect 28721 13277 28733 13280
rect 28767 13277 28779 13311
rect 28721 13271 28779 13277
rect 28813 13311 28871 13317
rect 28813 13277 28825 13311
rect 28859 13277 28871 13311
rect 30926 13308 30932 13320
rect 30887 13280 30932 13308
rect 28813 13271 28871 13277
rect 28316 13212 28488 13240
rect 28316 13200 28322 13212
rect 28626 13200 28632 13252
rect 28684 13240 28690 13252
rect 28828 13240 28856 13271
rect 30926 13268 30932 13280
rect 30984 13268 30990 13320
rect 31018 13268 31024 13320
rect 31076 13308 31082 13320
rect 31113 13311 31171 13317
rect 31113 13308 31125 13311
rect 31076 13280 31125 13308
rect 31076 13268 31082 13280
rect 31113 13277 31125 13280
rect 31159 13277 31171 13311
rect 31113 13271 31171 13277
rect 34698 13268 34704 13320
rect 34756 13308 34762 13320
rect 35969 13311 36027 13317
rect 35969 13308 35981 13311
rect 34756 13280 35981 13308
rect 34756 13268 34762 13280
rect 35969 13277 35981 13280
rect 36015 13277 36027 13311
rect 35969 13271 36027 13277
rect 28684 13212 28856 13240
rect 31573 13243 31631 13249
rect 28684 13200 28690 13212
rect 31573 13209 31585 13243
rect 31619 13240 31631 13243
rect 31662 13240 31668 13252
rect 31619 13212 31668 13240
rect 31619 13209 31631 13212
rect 31573 13203 31631 13209
rect 31662 13200 31668 13212
rect 31720 13200 31726 13252
rect 19334 13172 19340 13184
rect 14608 13144 19340 13172
rect 14608 13132 14614 13144
rect 19334 13132 19340 13144
rect 19392 13132 19398 13184
rect 21082 13172 21088 13184
rect 21043 13144 21088 13172
rect 21082 13132 21088 13144
rect 21140 13132 21146 13184
rect 21821 13175 21879 13181
rect 21821 13141 21833 13175
rect 21867 13172 21879 13175
rect 22186 13172 22192 13184
rect 21867 13144 22192 13172
rect 21867 13141 21879 13144
rect 21821 13135 21879 13141
rect 22186 13132 22192 13144
rect 22244 13132 22250 13184
rect 22462 13132 22468 13184
rect 22520 13172 22526 13184
rect 26789 13175 26847 13181
rect 26789 13172 26801 13175
rect 22520 13144 26801 13172
rect 22520 13132 22526 13144
rect 26789 13141 26801 13144
rect 26835 13141 26847 13175
rect 26789 13135 26847 13141
rect 30006 13132 30012 13184
rect 30064 13172 30070 13184
rect 34514 13172 34520 13184
rect 30064 13144 34520 13172
rect 30064 13132 30070 13144
rect 34514 13132 34520 13144
rect 34572 13132 34578 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 7926 12928 7932 12980
rect 7984 12928 7990 12980
rect 9600 12940 13032 12968
rect 7944 12900 7972 12928
rect 9600 12900 9628 12940
rect 11146 12900 11152 12912
rect 7668 12872 7972 12900
rect 9416 12872 9628 12900
rect 11107 12872 11152 12900
rect 7668 12841 7696 12872
rect 7653 12835 7711 12841
rect 7653 12801 7665 12835
rect 7699 12801 7711 12835
rect 7653 12795 7711 12801
rect 7920 12835 7978 12841
rect 7920 12801 7932 12835
rect 7966 12832 7978 12835
rect 9416 12832 9444 12872
rect 11146 12860 11152 12872
rect 11204 12860 11210 12912
rect 12158 12860 12164 12912
rect 12216 12900 12222 12912
rect 12894 12900 12900 12912
rect 12216 12872 12900 12900
rect 12216 12860 12222 12872
rect 12894 12860 12900 12872
rect 12952 12860 12958 12912
rect 7966 12804 9444 12832
rect 9493 12835 9551 12841
rect 7966 12801 7978 12804
rect 7920 12795 7978 12801
rect 9493 12801 9505 12835
rect 9539 12832 9551 12835
rect 12176 12832 12204 12860
rect 9539 12804 12204 12832
rect 12529 12835 12587 12841
rect 9539 12801 9551 12804
rect 9493 12795 9551 12801
rect 12529 12801 12541 12835
rect 12575 12801 12587 12835
rect 12710 12832 12716 12844
rect 12671 12804 12716 12832
rect 12529 12795 12587 12801
rect 9766 12764 9772 12776
rect 9727 12736 9772 12764
rect 9766 12724 9772 12736
rect 9824 12724 9830 12776
rect 12544 12764 12572 12795
rect 12710 12792 12716 12804
rect 12768 12792 12774 12844
rect 12805 12835 12863 12841
rect 12805 12801 12817 12835
rect 12851 12832 12863 12835
rect 13004 12832 13032 12940
rect 13354 12928 13360 12980
rect 13412 12968 13418 12980
rect 13725 12971 13783 12977
rect 13725 12968 13737 12971
rect 13412 12940 13737 12968
rect 13412 12928 13418 12940
rect 13725 12937 13737 12940
rect 13771 12937 13783 12971
rect 13725 12931 13783 12937
rect 14369 12971 14427 12977
rect 14369 12937 14381 12971
rect 14415 12968 14427 12971
rect 14642 12968 14648 12980
rect 14415 12940 14648 12968
rect 14415 12937 14427 12940
rect 14369 12931 14427 12937
rect 14642 12928 14648 12940
rect 14700 12928 14706 12980
rect 15933 12971 15991 12977
rect 15933 12937 15945 12971
rect 15979 12968 15991 12971
rect 16850 12968 16856 12980
rect 15979 12940 16856 12968
rect 15979 12937 15991 12940
rect 15933 12931 15991 12937
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 17770 12968 17776 12980
rect 17731 12940 17776 12968
rect 17770 12928 17776 12940
rect 17828 12928 17834 12980
rect 21082 12928 21088 12980
rect 21140 12968 21146 12980
rect 29730 12968 29736 12980
rect 21140 12940 22416 12968
rect 21140 12928 21146 12940
rect 13262 12900 13268 12912
rect 13223 12872 13268 12900
rect 13262 12860 13268 12872
rect 13320 12860 13326 12912
rect 13446 12860 13452 12912
rect 13504 12900 13510 12912
rect 16482 12900 16488 12912
rect 13504 12872 14136 12900
rect 13504 12860 13510 12872
rect 13998 12832 14004 12844
rect 12851 12804 14004 12832
rect 12851 12801 12863 12804
rect 12805 12795 12863 12801
rect 13998 12792 14004 12804
rect 14056 12792 14062 12844
rect 14108 12832 14136 12872
rect 15672 12872 16488 12900
rect 14366 12835 14424 12841
rect 14366 12832 14378 12835
rect 14108 12804 14378 12832
rect 14366 12801 14378 12804
rect 14412 12832 14424 12835
rect 14550 12832 14556 12844
rect 14412 12804 14556 12832
rect 14412 12801 14424 12804
rect 14366 12795 14424 12801
rect 14550 12792 14556 12804
rect 14608 12792 14614 12844
rect 15562 12792 15568 12844
rect 15620 12832 15626 12844
rect 15672 12841 15700 12872
rect 16482 12860 16488 12872
rect 16540 12860 16546 12912
rect 22005 12903 22063 12909
rect 22005 12900 22017 12903
rect 21100 12872 22017 12900
rect 15657 12835 15715 12841
rect 15657 12832 15669 12835
rect 15620 12804 15669 12832
rect 15620 12792 15626 12804
rect 15657 12801 15669 12804
rect 15703 12801 15715 12835
rect 15657 12795 15715 12801
rect 15746 12792 15752 12844
rect 15804 12832 15810 12844
rect 15804 12804 15849 12832
rect 15804 12792 15810 12804
rect 17218 12792 17224 12844
rect 17276 12832 17282 12844
rect 17405 12835 17463 12841
rect 17405 12832 17417 12835
rect 17276 12804 17417 12832
rect 17276 12792 17282 12804
rect 17405 12801 17417 12804
rect 17451 12801 17463 12835
rect 17405 12795 17463 12801
rect 17494 12792 17500 12844
rect 17552 12832 17558 12844
rect 17589 12835 17647 12841
rect 17589 12832 17601 12835
rect 17552 12804 17601 12832
rect 17552 12792 17558 12804
rect 17589 12801 17601 12804
rect 17635 12801 17647 12835
rect 17589 12795 17647 12801
rect 19334 12792 19340 12844
rect 19392 12832 19398 12844
rect 19521 12835 19579 12841
rect 19521 12832 19533 12835
rect 19392 12804 19533 12832
rect 19392 12792 19398 12804
rect 19521 12801 19533 12804
rect 19567 12801 19579 12835
rect 19702 12832 19708 12844
rect 19663 12804 19708 12832
rect 19521 12795 19579 12801
rect 14826 12764 14832 12776
rect 12544 12736 13768 12764
rect 14787 12736 14832 12764
rect 12710 12656 12716 12708
rect 12768 12696 12774 12708
rect 13446 12696 13452 12708
rect 12768 12668 13452 12696
rect 12768 12656 12774 12668
rect 13446 12656 13452 12668
rect 13504 12656 13510 12708
rect 13630 12696 13636 12708
rect 13591 12668 13636 12696
rect 13630 12656 13636 12668
rect 13688 12656 13694 12708
rect 13740 12696 13768 12736
rect 14826 12724 14832 12736
rect 14884 12724 14890 12776
rect 15933 12767 15991 12773
rect 15933 12733 15945 12767
rect 15979 12764 15991 12767
rect 17236 12764 17264 12792
rect 19536 12764 19564 12795
rect 19702 12792 19708 12804
rect 19760 12792 19766 12844
rect 19797 12835 19855 12841
rect 19797 12801 19809 12835
rect 19843 12832 19855 12835
rect 19978 12832 19984 12844
rect 19843 12804 19984 12832
rect 19843 12801 19855 12804
rect 19797 12795 19855 12801
rect 19978 12792 19984 12804
rect 20036 12792 20042 12844
rect 21100 12841 21128 12872
rect 22005 12869 22017 12872
rect 22051 12869 22063 12903
rect 22005 12863 22063 12869
rect 21085 12835 21143 12841
rect 21085 12801 21097 12835
rect 21131 12801 21143 12835
rect 21085 12795 21143 12801
rect 21174 12792 21180 12844
rect 21232 12832 21238 12844
rect 21232 12804 21277 12832
rect 21232 12792 21238 12804
rect 21358 12792 21364 12844
rect 21416 12832 21422 12844
rect 21453 12835 21511 12841
rect 21453 12832 21465 12835
rect 21416 12804 21465 12832
rect 21416 12792 21422 12804
rect 21453 12801 21465 12804
rect 21499 12801 21511 12835
rect 22186 12832 22192 12844
rect 22147 12804 22192 12832
rect 21453 12795 21511 12801
rect 22186 12792 22192 12804
rect 22244 12792 22250 12844
rect 22388 12841 22416 12940
rect 25792 12940 29736 12968
rect 25130 12860 25136 12912
rect 25188 12900 25194 12912
rect 25792 12900 25820 12940
rect 29730 12928 29736 12940
rect 29788 12928 29794 12980
rect 32030 12928 32036 12980
rect 32088 12968 32094 12980
rect 33045 12971 33103 12977
rect 33045 12968 33057 12971
rect 32088 12940 33057 12968
rect 32088 12928 32094 12940
rect 33045 12937 33057 12940
rect 33091 12937 33103 12971
rect 33045 12931 33103 12937
rect 25188 12872 25820 12900
rect 25188 12860 25194 12872
rect 22373 12835 22431 12841
rect 22373 12801 22385 12835
rect 22419 12801 22431 12835
rect 25406 12832 25412 12844
rect 25367 12804 25412 12832
rect 22373 12795 22431 12801
rect 25406 12792 25412 12804
rect 25464 12792 25470 12844
rect 25590 12832 25596 12844
rect 25551 12804 25596 12832
rect 25590 12792 25596 12804
rect 25648 12792 25654 12844
rect 25792 12841 25820 12872
rect 28736 12872 29040 12900
rect 25777 12835 25835 12841
rect 25777 12801 25789 12835
rect 25823 12801 25835 12835
rect 25777 12795 25835 12801
rect 25869 12835 25927 12841
rect 25869 12801 25881 12835
rect 25915 12832 25927 12835
rect 27798 12832 27804 12844
rect 25915 12804 27804 12832
rect 25915 12801 25927 12804
rect 25869 12795 25927 12801
rect 27798 12792 27804 12804
rect 27856 12832 27862 12844
rect 28736 12841 28764 12872
rect 28261 12835 28319 12841
rect 28261 12832 28273 12835
rect 27856 12804 28273 12832
rect 27856 12792 27862 12804
rect 28261 12801 28273 12804
rect 28307 12801 28319 12835
rect 28261 12795 28319 12801
rect 28721 12835 28779 12841
rect 28721 12801 28733 12835
rect 28767 12801 28779 12835
rect 28721 12795 28779 12801
rect 28905 12835 28963 12841
rect 28905 12801 28917 12835
rect 28951 12801 28963 12835
rect 29012 12832 29040 12872
rect 29086 12860 29092 12912
rect 29144 12900 29150 12912
rect 29273 12903 29331 12909
rect 29273 12900 29285 12903
rect 29144 12872 29285 12900
rect 29144 12860 29150 12872
rect 29273 12869 29285 12872
rect 29319 12869 29331 12903
rect 29273 12863 29331 12869
rect 29178 12832 29184 12844
rect 29012 12804 29184 12832
rect 28905 12795 28963 12801
rect 20070 12764 20076 12776
rect 15979 12736 17816 12764
rect 19536 12736 20076 12764
rect 15979 12733 15991 12736
rect 15933 12727 15991 12733
rect 17788 12708 17816 12736
rect 20070 12724 20076 12736
rect 20128 12724 20134 12776
rect 21542 12724 21548 12776
rect 21600 12764 21606 12776
rect 22462 12764 22468 12776
rect 21600 12736 22468 12764
rect 21600 12724 21606 12736
rect 22462 12724 22468 12736
rect 22520 12724 22526 12776
rect 27982 12764 27988 12776
rect 27943 12736 27988 12764
rect 27982 12724 27988 12736
rect 28040 12724 28046 12776
rect 28276 12764 28304 12795
rect 28810 12764 28816 12776
rect 28276 12736 28816 12764
rect 28810 12724 28816 12736
rect 28868 12724 28874 12776
rect 28920 12764 28948 12795
rect 29178 12792 29184 12804
rect 29236 12792 29242 12844
rect 32953 12835 33011 12841
rect 32953 12801 32965 12835
rect 32999 12832 33011 12835
rect 33870 12832 33876 12844
rect 32999 12804 33876 12832
rect 32999 12801 33011 12804
rect 32953 12795 33011 12801
rect 33870 12792 33876 12804
rect 33928 12792 33934 12844
rect 32858 12764 32864 12776
rect 28920 12736 32864 12764
rect 16758 12696 16764 12708
rect 13740 12668 16764 12696
rect 16758 12656 16764 12668
rect 16816 12656 16822 12708
rect 17770 12656 17776 12708
rect 17828 12656 17834 12708
rect 28169 12699 28227 12705
rect 28169 12665 28181 12699
rect 28215 12696 28227 12699
rect 28920 12696 28948 12736
rect 32858 12724 32864 12736
rect 32916 12724 32922 12776
rect 33042 12724 33048 12776
rect 33100 12764 33106 12776
rect 33137 12767 33195 12773
rect 33137 12764 33149 12767
rect 33100 12736 33149 12764
rect 33100 12724 33106 12736
rect 33137 12733 33149 12736
rect 33183 12733 33195 12767
rect 33137 12727 33195 12733
rect 28215 12668 28948 12696
rect 29181 12699 29239 12705
rect 28215 12665 28227 12668
rect 28169 12659 28227 12665
rect 29181 12665 29193 12699
rect 29227 12696 29239 12699
rect 29227 12668 32996 12696
rect 29227 12665 29239 12668
rect 29181 12659 29239 12665
rect 9033 12631 9091 12637
rect 9033 12597 9045 12631
rect 9079 12628 9091 12631
rect 9214 12628 9220 12640
rect 9079 12600 9220 12628
rect 9079 12597 9091 12600
rect 9033 12591 9091 12597
rect 9214 12588 9220 12600
rect 9272 12588 9278 12640
rect 12526 12628 12532 12640
rect 12487 12600 12532 12628
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 14182 12628 14188 12640
rect 14143 12600 14188 12628
rect 14182 12588 14188 12600
rect 14240 12588 14246 12640
rect 14737 12631 14795 12637
rect 14737 12597 14749 12631
rect 14783 12628 14795 12631
rect 15654 12628 15660 12640
rect 14783 12600 15660 12628
rect 14783 12597 14795 12600
rect 14737 12591 14795 12597
rect 15654 12588 15660 12600
rect 15712 12588 15718 12640
rect 19337 12631 19395 12637
rect 19337 12597 19349 12631
rect 19383 12628 19395 12631
rect 19702 12628 19708 12640
rect 19383 12600 19708 12628
rect 19383 12597 19395 12600
rect 19337 12591 19395 12597
rect 19702 12588 19708 12600
rect 19760 12588 19766 12640
rect 20622 12588 20628 12640
rect 20680 12628 20686 12640
rect 20901 12631 20959 12637
rect 20901 12628 20913 12631
rect 20680 12600 20913 12628
rect 20680 12588 20686 12600
rect 20901 12597 20913 12600
rect 20947 12597 20959 12631
rect 20901 12591 20959 12597
rect 21361 12631 21419 12637
rect 21361 12597 21373 12631
rect 21407 12628 21419 12631
rect 21450 12628 21456 12640
rect 21407 12600 21456 12628
rect 21407 12597 21419 12600
rect 21361 12591 21419 12597
rect 21450 12588 21456 12600
rect 21508 12588 21514 12640
rect 27798 12628 27804 12640
rect 27759 12600 27804 12628
rect 27798 12588 27804 12600
rect 27856 12588 27862 12640
rect 32582 12628 32588 12640
rect 32543 12600 32588 12628
rect 32582 12588 32588 12600
rect 32640 12588 32646 12640
rect 32968 12628 32996 12668
rect 35526 12628 35532 12640
rect 32968 12600 35532 12628
rect 35526 12588 35532 12600
rect 35584 12588 35590 12640
rect 38286 12628 38292 12640
rect 38247 12600 38292 12628
rect 38286 12588 38292 12600
rect 38344 12588 38350 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 9677 12427 9735 12433
rect 9677 12393 9689 12427
rect 9723 12424 9735 12427
rect 10594 12424 10600 12436
rect 9723 12396 10600 12424
rect 9723 12393 9735 12396
rect 9677 12387 9735 12393
rect 10594 12384 10600 12396
rect 10652 12384 10658 12436
rect 13170 12424 13176 12436
rect 13131 12396 13176 12424
rect 13170 12384 13176 12396
rect 13228 12384 13234 12436
rect 15010 12424 15016 12436
rect 14971 12396 15016 12424
rect 15010 12384 15016 12396
rect 15068 12384 15074 12436
rect 15654 12384 15660 12436
rect 15712 12424 15718 12436
rect 16945 12427 17003 12433
rect 16945 12424 16957 12427
rect 15712 12396 16957 12424
rect 15712 12384 15718 12396
rect 16945 12393 16957 12396
rect 16991 12393 17003 12427
rect 16945 12387 17003 12393
rect 17034 12384 17040 12436
rect 17092 12424 17098 12436
rect 17586 12424 17592 12436
rect 17092 12396 17592 12424
rect 17092 12384 17098 12396
rect 17586 12384 17592 12396
rect 17644 12384 17650 12436
rect 18782 12384 18788 12436
rect 18840 12424 18846 12436
rect 20162 12424 20168 12436
rect 18840 12396 20168 12424
rect 18840 12384 18846 12396
rect 20162 12384 20168 12396
rect 20220 12424 20226 12436
rect 20714 12424 20720 12436
rect 20220 12396 20720 12424
rect 20220 12384 20226 12396
rect 20714 12384 20720 12396
rect 20772 12384 20778 12436
rect 20993 12427 21051 12433
rect 20993 12393 21005 12427
rect 21039 12424 21051 12427
rect 21174 12424 21180 12436
rect 21039 12396 21180 12424
rect 21039 12393 21051 12396
rect 20993 12387 21051 12393
rect 21174 12384 21180 12396
rect 21232 12384 21238 12436
rect 25409 12427 25467 12433
rect 21284 12396 24532 12424
rect 11790 12316 11796 12368
rect 11848 12356 11854 12368
rect 12345 12359 12403 12365
rect 12345 12356 12357 12359
rect 11848 12328 12357 12356
rect 11848 12316 11854 12328
rect 12345 12325 12357 12328
rect 12391 12325 12403 12359
rect 12345 12319 12403 12325
rect 15378 12316 15384 12368
rect 15436 12356 15442 12368
rect 16301 12359 16359 12365
rect 16301 12356 16313 12359
rect 15436 12328 16313 12356
rect 15436 12316 15442 12328
rect 16301 12325 16313 12328
rect 16347 12356 16359 12359
rect 21284 12356 21312 12396
rect 21542 12356 21548 12368
rect 16347 12328 16620 12356
rect 16347 12325 16359 12328
rect 16301 12319 16359 12325
rect 9214 12288 9220 12300
rect 9175 12260 9220 12288
rect 9214 12248 9220 12260
rect 9272 12248 9278 12300
rect 12437 12291 12495 12297
rect 12437 12257 12449 12291
rect 12483 12288 12495 12291
rect 12618 12288 12624 12300
rect 12483 12260 12624 12288
rect 12483 12257 12495 12260
rect 12437 12251 12495 12257
rect 12618 12248 12624 12260
rect 12676 12288 12682 12300
rect 14182 12288 14188 12300
rect 12676 12260 14188 12288
rect 12676 12248 12682 12260
rect 14182 12248 14188 12260
rect 14240 12248 14246 12300
rect 15562 12288 15568 12300
rect 15523 12260 15568 12288
rect 15562 12248 15568 12260
rect 15620 12248 15626 12300
rect 16390 12248 16396 12300
rect 16448 12288 16454 12300
rect 16485 12291 16543 12297
rect 16485 12288 16497 12291
rect 16448 12260 16497 12288
rect 16448 12248 16454 12260
rect 16485 12257 16497 12260
rect 16531 12257 16543 12291
rect 16592 12288 16620 12328
rect 17236 12328 21312 12356
rect 21376 12328 21548 12356
rect 17236 12300 17264 12328
rect 16942 12288 16948 12300
rect 16592 12260 16948 12288
rect 16485 12251 16543 12257
rect 16942 12248 16948 12260
rect 17000 12288 17006 12300
rect 17129 12291 17187 12297
rect 17129 12288 17141 12291
rect 17000 12260 17141 12288
rect 17000 12248 17006 12260
rect 17129 12257 17141 12260
rect 17175 12257 17187 12291
rect 17129 12251 17187 12257
rect 17218 12248 17224 12300
rect 17276 12288 17282 12300
rect 18673 12291 18731 12297
rect 17276 12260 17321 12288
rect 17276 12248 17282 12260
rect 18673 12257 18685 12291
rect 18719 12288 18731 12291
rect 19889 12291 19947 12297
rect 18719 12260 19656 12288
rect 18719 12257 18731 12260
rect 18673 12251 18731 12257
rect 9306 12220 9312 12232
rect 9267 12192 9312 12220
rect 9306 12180 9312 12192
rect 9364 12180 9370 12232
rect 12161 12223 12219 12229
rect 12161 12189 12173 12223
rect 12207 12189 12219 12223
rect 12161 12183 12219 12189
rect 12253 12223 12311 12229
rect 12253 12189 12265 12223
rect 12299 12220 12311 12223
rect 12342 12220 12348 12232
rect 12299 12192 12348 12220
rect 12299 12189 12311 12192
rect 12253 12183 12311 12189
rect 12176 12152 12204 12183
rect 12342 12180 12348 12192
rect 12400 12180 12406 12232
rect 13173 12223 13231 12229
rect 13173 12189 13185 12223
rect 13219 12220 13231 12223
rect 13262 12220 13268 12232
rect 13219 12192 13268 12220
rect 13219 12189 13231 12192
rect 13173 12183 13231 12189
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 13357 12223 13415 12229
rect 13357 12189 13369 12223
rect 13403 12220 13415 12223
rect 13446 12220 13452 12232
rect 13403 12192 13452 12220
rect 13403 12189 13415 12192
rect 13357 12183 13415 12189
rect 13446 12180 13452 12192
rect 13504 12180 13510 12232
rect 16209 12223 16267 12229
rect 16209 12189 16221 12223
rect 16255 12189 16267 12223
rect 16209 12183 16267 12189
rect 12434 12152 12440 12164
rect 12176 12124 12440 12152
rect 12434 12112 12440 12124
rect 12492 12112 12498 12164
rect 15289 12155 15347 12161
rect 15289 12121 15301 12155
rect 15335 12152 15347 12155
rect 15654 12152 15660 12164
rect 15335 12124 15660 12152
rect 15335 12121 15347 12124
rect 15289 12115 15347 12121
rect 15654 12112 15660 12124
rect 15712 12112 15718 12164
rect 15470 12084 15476 12096
rect 15431 12056 15476 12084
rect 15470 12044 15476 12056
rect 15528 12044 15534 12096
rect 16224 12084 16252 12183
rect 17034 12180 17040 12232
rect 17092 12220 17098 12232
rect 17313 12223 17371 12229
rect 17313 12220 17325 12223
rect 17092 12192 17325 12220
rect 17092 12180 17098 12192
rect 17313 12189 17325 12192
rect 17359 12189 17371 12223
rect 17313 12183 17371 12189
rect 17405 12223 17463 12229
rect 17405 12189 17417 12223
rect 17451 12189 17463 12223
rect 18782 12220 18788 12232
rect 18743 12192 18788 12220
rect 17405 12183 17463 12189
rect 16485 12155 16543 12161
rect 16485 12121 16497 12155
rect 16531 12152 16543 12155
rect 17420 12152 17448 12183
rect 18782 12180 18788 12192
rect 18840 12180 18846 12232
rect 18877 12223 18935 12229
rect 18877 12189 18889 12223
rect 18923 12220 18935 12223
rect 19058 12220 19064 12232
rect 18923 12192 19064 12220
rect 18923 12189 18935 12192
rect 18877 12183 18935 12189
rect 19058 12180 19064 12192
rect 19116 12180 19122 12232
rect 19628 12229 19656 12260
rect 19889 12257 19901 12291
rect 19935 12288 19947 12291
rect 21376 12288 21404 12328
rect 21542 12316 21548 12328
rect 21600 12316 21606 12368
rect 21634 12288 21640 12300
rect 19935 12260 21404 12288
rect 19935 12257 19947 12260
rect 19889 12251 19947 12257
rect 19613 12223 19671 12229
rect 19613 12189 19625 12223
rect 19659 12189 19671 12223
rect 19613 12183 19671 12189
rect 19702 12180 19708 12232
rect 19760 12220 19766 12232
rect 19981 12223 20039 12229
rect 19981 12220 19993 12223
rect 19760 12192 19805 12220
rect 19904 12192 19993 12220
rect 19760 12180 19766 12192
rect 16531 12124 17448 12152
rect 18601 12155 18659 12161
rect 16531 12121 16543 12124
rect 16485 12115 16543 12121
rect 18601 12121 18613 12155
rect 18647 12152 18659 12155
rect 19334 12152 19340 12164
rect 18647 12124 19340 12152
rect 18647 12121 18659 12124
rect 18601 12115 18659 12121
rect 19334 12112 19340 12124
rect 19392 12112 19398 12164
rect 17678 12084 17684 12096
rect 16224 12056 17684 12084
rect 17678 12044 17684 12056
rect 17736 12044 17742 12096
rect 18874 12044 18880 12096
rect 18932 12084 18938 12096
rect 19429 12087 19487 12093
rect 19429 12084 19441 12087
rect 18932 12056 19441 12084
rect 18932 12044 18938 12056
rect 19429 12053 19441 12056
rect 19475 12053 19487 12087
rect 19904 12084 19932 12192
rect 19981 12189 19993 12192
rect 20027 12189 20039 12223
rect 19981 12183 20039 12189
rect 20070 12180 20076 12232
rect 20128 12220 20134 12232
rect 21376 12229 21404 12260
rect 21468 12260 21640 12288
rect 21468 12229 21496 12260
rect 21634 12248 21640 12260
rect 21692 12288 21698 12300
rect 22005 12291 22063 12297
rect 22005 12288 22017 12291
rect 21692 12260 22017 12288
rect 21692 12248 21698 12260
rect 22005 12257 22017 12260
rect 22051 12257 22063 12291
rect 24504 12288 24532 12396
rect 25409 12393 25421 12427
rect 25455 12424 25467 12427
rect 26326 12424 26332 12436
rect 25455 12396 26332 12424
rect 25455 12393 25467 12396
rect 25409 12387 25467 12393
rect 26326 12384 26332 12396
rect 26384 12384 26390 12436
rect 27982 12384 27988 12436
rect 28040 12424 28046 12436
rect 28261 12427 28319 12433
rect 28261 12424 28273 12427
rect 28040 12396 28273 12424
rect 28040 12384 28046 12396
rect 28261 12393 28273 12396
rect 28307 12393 28319 12427
rect 28994 12424 29000 12436
rect 28955 12396 29000 12424
rect 28261 12387 28319 12393
rect 28994 12384 29000 12396
rect 29052 12384 29058 12436
rect 33226 12424 33232 12436
rect 29288 12396 33232 12424
rect 24581 12359 24639 12365
rect 24581 12325 24593 12359
rect 24627 12356 24639 12359
rect 24627 12328 25176 12356
rect 24627 12325 24639 12328
rect 24581 12319 24639 12325
rect 25148 12288 25176 12328
rect 25777 12291 25835 12297
rect 25777 12288 25789 12291
rect 24504 12260 24992 12288
rect 25148 12260 25789 12288
rect 22005 12251 22063 12257
rect 21177 12223 21235 12229
rect 21177 12220 21189 12223
rect 20128 12192 21189 12220
rect 20128 12180 20134 12192
rect 21177 12189 21189 12192
rect 21223 12189 21235 12223
rect 21177 12183 21235 12189
rect 21361 12223 21419 12229
rect 21361 12189 21373 12223
rect 21407 12189 21419 12223
rect 21361 12183 21419 12189
rect 21453 12223 21511 12229
rect 21453 12189 21465 12223
rect 21499 12189 21511 12223
rect 21910 12220 21916 12232
rect 21871 12192 21916 12220
rect 21453 12183 21511 12189
rect 21910 12180 21916 12192
rect 21968 12180 21974 12232
rect 22097 12223 22155 12229
rect 22097 12189 22109 12223
rect 22143 12189 22155 12223
rect 22097 12183 22155 12189
rect 20438 12112 20444 12164
rect 20496 12152 20502 12164
rect 22112 12152 22140 12183
rect 22278 12180 22284 12232
rect 22336 12220 22342 12232
rect 24854 12220 24860 12232
rect 22336 12192 24860 12220
rect 22336 12180 22342 12192
rect 24854 12180 24860 12192
rect 24912 12180 24918 12232
rect 24964 12220 24992 12260
rect 25777 12257 25789 12260
rect 25823 12257 25835 12291
rect 25958 12288 25964 12300
rect 25919 12260 25964 12288
rect 25777 12251 25835 12257
rect 25958 12248 25964 12260
rect 26016 12248 26022 12300
rect 28442 12248 28448 12300
rect 28500 12288 28506 12300
rect 28500 12260 28764 12288
rect 28500 12248 28506 12260
rect 27614 12220 27620 12232
rect 24964 12192 27620 12220
rect 27614 12180 27620 12192
rect 27672 12180 27678 12232
rect 28258 12220 28264 12232
rect 28219 12192 28264 12220
rect 28258 12180 28264 12192
rect 28316 12180 28322 12232
rect 28537 12223 28595 12229
rect 28537 12189 28549 12223
rect 28583 12220 28595 12223
rect 28626 12220 28632 12232
rect 28583 12192 28632 12220
rect 28583 12189 28595 12192
rect 28537 12183 28595 12189
rect 28626 12180 28632 12192
rect 28684 12180 28690 12232
rect 28736 12220 28764 12260
rect 28810 12248 28816 12300
rect 28868 12288 28874 12300
rect 28868 12260 29224 12288
rect 28868 12248 28874 12260
rect 28902 12220 28908 12232
rect 28736 12192 28908 12220
rect 28902 12180 28908 12192
rect 28960 12220 28966 12232
rect 29196 12229 29224 12260
rect 28997 12223 29055 12229
rect 28997 12220 29009 12223
rect 28960 12192 29009 12220
rect 28960 12180 28966 12192
rect 28997 12189 29009 12192
rect 29043 12189 29055 12223
rect 28997 12183 29055 12189
rect 29181 12223 29239 12229
rect 29181 12189 29193 12223
rect 29227 12189 29239 12223
rect 29181 12183 29239 12189
rect 20496 12124 22140 12152
rect 24581 12155 24639 12161
rect 20496 12112 20502 12124
rect 24581 12121 24593 12155
rect 24627 12152 24639 12155
rect 25774 12152 25780 12164
rect 24627 12124 25780 12152
rect 24627 12121 24639 12124
rect 24581 12115 24639 12121
rect 25774 12112 25780 12124
rect 25832 12112 25838 12164
rect 29288 12152 29316 12396
rect 33226 12384 33232 12396
rect 33284 12384 33290 12436
rect 33870 12424 33876 12436
rect 33831 12396 33876 12424
rect 33870 12384 33876 12396
rect 33928 12384 33934 12436
rect 30834 12248 30840 12300
rect 30892 12288 30898 12300
rect 31665 12291 31723 12297
rect 31665 12288 31677 12291
rect 30892 12260 31677 12288
rect 30892 12248 30898 12260
rect 31665 12257 31677 12260
rect 31711 12257 31723 12291
rect 31665 12251 31723 12257
rect 34422 12248 34428 12300
rect 34480 12288 34486 12300
rect 35529 12291 35587 12297
rect 35529 12288 35541 12291
rect 34480 12260 35541 12288
rect 34480 12248 34486 12260
rect 35529 12257 35541 12260
rect 35575 12257 35587 12291
rect 35529 12251 35587 12257
rect 35710 12248 35716 12300
rect 35768 12288 35774 12300
rect 36817 12291 36875 12297
rect 36817 12288 36829 12291
rect 35768 12260 36829 12288
rect 35768 12248 35774 12260
rect 36817 12257 36829 12260
rect 36863 12257 36875 12291
rect 36817 12251 36875 12257
rect 30374 12180 30380 12232
rect 30432 12220 30438 12232
rect 32490 12220 32496 12232
rect 30432 12192 32496 12220
rect 30432 12180 30438 12192
rect 32490 12180 32496 12192
rect 32548 12180 32554 12232
rect 32582 12180 32588 12232
rect 32640 12220 32646 12232
rect 32749 12223 32807 12229
rect 32749 12220 32761 12223
rect 32640 12192 32761 12220
rect 32640 12180 32646 12192
rect 32749 12189 32761 12192
rect 32795 12189 32807 12223
rect 32749 12183 32807 12189
rect 33042 12180 33048 12232
rect 33100 12220 33106 12232
rect 38194 12220 38200 12232
rect 33100 12192 38200 12220
rect 33100 12180 33106 12192
rect 38194 12180 38200 12192
rect 38252 12180 38258 12232
rect 28460 12124 29316 12152
rect 31573 12155 31631 12161
rect 20806 12084 20812 12096
rect 19904 12056 20812 12084
rect 19429 12047 19487 12053
rect 20806 12044 20812 12056
rect 20864 12084 20870 12096
rect 21358 12084 21364 12096
rect 20864 12056 21364 12084
rect 20864 12044 20870 12056
rect 21358 12044 21364 12056
rect 21416 12044 21422 12096
rect 24762 12084 24768 12096
rect 24723 12056 24768 12084
rect 24762 12044 24768 12056
rect 24820 12044 24826 12096
rect 25866 12084 25872 12096
rect 25827 12056 25872 12084
rect 25866 12044 25872 12056
rect 25924 12044 25930 12096
rect 27798 12044 27804 12096
rect 27856 12084 27862 12096
rect 28258 12084 28264 12096
rect 27856 12056 28264 12084
rect 27856 12044 27862 12056
rect 28258 12044 28264 12056
rect 28316 12084 28322 12096
rect 28460 12093 28488 12124
rect 31573 12121 31585 12155
rect 31619 12152 31631 12155
rect 32030 12152 32036 12164
rect 31619 12124 32036 12152
rect 31619 12121 31631 12124
rect 31573 12115 31631 12121
rect 32030 12112 32036 12124
rect 32088 12112 32094 12164
rect 34330 12112 34336 12164
rect 34388 12152 34394 12164
rect 35345 12155 35403 12161
rect 34388 12124 35112 12152
rect 34388 12112 34394 12124
rect 28445 12087 28503 12093
rect 28445 12084 28457 12087
rect 28316 12056 28457 12084
rect 28316 12044 28322 12056
rect 28445 12053 28457 12056
rect 28491 12053 28503 12087
rect 31110 12084 31116 12096
rect 31071 12056 31116 12084
rect 28445 12047 28503 12053
rect 31110 12044 31116 12056
rect 31168 12044 31174 12096
rect 31478 12084 31484 12096
rect 31439 12056 31484 12084
rect 31478 12044 31484 12056
rect 31536 12044 31542 12096
rect 34790 12044 34796 12096
rect 34848 12084 34854 12096
rect 34977 12087 35035 12093
rect 34977 12084 34989 12087
rect 34848 12056 34989 12084
rect 34848 12044 34854 12056
rect 34977 12053 34989 12056
rect 35023 12053 35035 12087
rect 35084 12084 35112 12124
rect 35345 12121 35357 12155
rect 35391 12152 35403 12155
rect 35802 12152 35808 12164
rect 35391 12124 35808 12152
rect 35391 12121 35403 12124
rect 35345 12115 35403 12121
rect 35802 12112 35808 12124
rect 35860 12112 35866 12164
rect 37084 12155 37142 12161
rect 37084 12121 37096 12155
rect 37130 12152 37142 12155
rect 37458 12152 37464 12164
rect 37130 12124 37464 12152
rect 37130 12121 37142 12124
rect 37084 12115 37142 12121
rect 37458 12112 37464 12124
rect 37516 12112 37522 12164
rect 35437 12087 35495 12093
rect 35437 12084 35449 12087
rect 35084 12056 35449 12084
rect 34977 12047 35035 12053
rect 35437 12053 35449 12056
rect 35483 12084 35495 12087
rect 35710 12084 35716 12096
rect 35483 12056 35716 12084
rect 35483 12053 35495 12056
rect 35437 12047 35495 12053
rect 35710 12044 35716 12056
rect 35768 12044 35774 12096
rect 37826 12044 37832 12096
rect 37884 12084 37890 12096
rect 38197 12087 38255 12093
rect 38197 12084 38209 12087
rect 37884 12056 38209 12084
rect 37884 12044 37890 12056
rect 38197 12053 38209 12056
rect 38243 12053 38255 12087
rect 38197 12047 38255 12053
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 9306 11880 9312 11892
rect 9267 11852 9312 11880
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 9766 11840 9772 11892
rect 9824 11880 9830 11892
rect 10413 11883 10471 11889
rect 10413 11880 10425 11883
rect 9824 11852 10425 11880
rect 9824 11840 9830 11852
rect 10413 11849 10425 11852
rect 10459 11849 10471 11883
rect 14737 11883 14795 11889
rect 14737 11880 14749 11883
rect 10413 11843 10471 11849
rect 12406 11852 14749 11880
rect 12406 11824 12434 11852
rect 14737 11849 14749 11852
rect 14783 11849 14795 11883
rect 14737 11843 14795 11849
rect 15105 11883 15163 11889
rect 15105 11849 15117 11883
rect 15151 11880 15163 11883
rect 15470 11880 15476 11892
rect 15151 11852 15476 11880
rect 15151 11849 15163 11852
rect 15105 11843 15163 11849
rect 15470 11840 15476 11852
rect 15528 11880 15534 11892
rect 16758 11880 16764 11892
rect 15528 11852 16764 11880
rect 15528 11840 15534 11852
rect 16758 11840 16764 11852
rect 16816 11840 16822 11892
rect 19058 11880 19064 11892
rect 19019 11852 19064 11880
rect 19058 11840 19064 11852
rect 19116 11840 19122 11892
rect 19334 11840 19340 11892
rect 19392 11880 19398 11892
rect 19613 11883 19671 11889
rect 19613 11880 19625 11883
rect 19392 11852 19625 11880
rect 19392 11840 19398 11852
rect 19613 11849 19625 11852
rect 19659 11849 19671 11883
rect 19613 11843 19671 11849
rect 19702 11840 19708 11892
rect 19760 11880 19766 11892
rect 20254 11880 20260 11892
rect 19760 11852 20260 11880
rect 19760 11840 19766 11852
rect 20254 11840 20260 11852
rect 20312 11840 20318 11892
rect 24765 11883 24823 11889
rect 24765 11849 24777 11883
rect 24811 11849 24823 11883
rect 25222 11880 25228 11892
rect 25183 11852 25228 11880
rect 24765 11843 24823 11849
rect 8196 11815 8254 11821
rect 8196 11781 8208 11815
rect 8242 11812 8254 11815
rect 11054 11812 11060 11824
rect 8242 11784 11060 11812
rect 8242 11781 8254 11784
rect 8196 11775 8254 11781
rect 11054 11772 11060 11784
rect 11112 11772 11118 11824
rect 12342 11812 12348 11824
rect 12303 11784 12348 11812
rect 12342 11772 12348 11784
rect 12400 11784 12434 11824
rect 12529 11815 12587 11821
rect 12400 11772 12406 11784
rect 12529 11781 12541 11815
rect 12575 11812 12587 11815
rect 12618 11812 12624 11824
rect 12575 11784 12624 11812
rect 12575 11781 12587 11784
rect 12529 11775 12587 11781
rect 12618 11772 12624 11784
rect 12676 11772 12682 11824
rect 17494 11812 17500 11824
rect 17407 11784 17500 11812
rect 17494 11772 17500 11784
rect 17552 11812 17558 11824
rect 21634 11812 21640 11824
rect 17552 11784 21640 11812
rect 17552 11772 17558 11784
rect 10597 11747 10655 11753
rect 10597 11744 10609 11747
rect 10428 11716 10609 11744
rect 7926 11676 7932 11688
rect 7887 11648 7932 11676
rect 7926 11636 7932 11648
rect 7984 11636 7990 11688
rect 10428 11608 10456 11716
rect 10597 11713 10609 11716
rect 10643 11713 10655 11747
rect 10778 11744 10784 11756
rect 10739 11716 10784 11744
rect 10597 11707 10655 11713
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 10873 11747 10931 11753
rect 10873 11713 10885 11747
rect 10919 11713 10931 11747
rect 10873 11707 10931 11713
rect 15197 11747 15255 11753
rect 15197 11713 15209 11747
rect 15243 11744 15255 11747
rect 15654 11744 15660 11756
rect 15243 11716 15660 11744
rect 15243 11713 15255 11716
rect 15197 11707 15255 11713
rect 10502 11636 10508 11688
rect 10560 11676 10566 11688
rect 10888 11676 10916 11707
rect 15654 11704 15660 11716
rect 15712 11704 15718 11756
rect 17681 11747 17739 11753
rect 17681 11713 17693 11747
rect 17727 11744 17739 11747
rect 17770 11744 17776 11756
rect 17727 11716 17776 11744
rect 17727 11713 17739 11716
rect 17681 11707 17739 11713
rect 17770 11704 17776 11716
rect 17828 11704 17834 11756
rect 19168 11753 19196 11784
rect 21634 11772 21640 11784
rect 21692 11772 21698 11824
rect 23474 11812 23480 11824
rect 22940 11784 23480 11812
rect 18969 11747 19027 11753
rect 18969 11713 18981 11747
rect 19015 11713 19027 11747
rect 18969 11707 19027 11713
rect 19153 11747 19211 11753
rect 19153 11713 19165 11747
rect 19199 11713 19211 11747
rect 19153 11707 19211 11713
rect 19797 11747 19855 11753
rect 19797 11713 19809 11747
rect 19843 11713 19855 11747
rect 19978 11744 19984 11756
rect 19939 11716 19984 11744
rect 19797 11707 19855 11713
rect 15378 11676 15384 11688
rect 10560 11648 10916 11676
rect 15339 11648 15384 11676
rect 10560 11636 10566 11648
rect 15378 11636 15384 11648
rect 15436 11636 15442 11688
rect 18984 11676 19012 11707
rect 19334 11676 19340 11688
rect 18984 11648 19340 11676
rect 19334 11636 19340 11648
rect 19392 11676 19398 11688
rect 19702 11676 19708 11688
rect 19392 11648 19708 11676
rect 19392 11636 19398 11648
rect 19702 11636 19708 11648
rect 19760 11636 19766 11688
rect 19812 11676 19840 11707
rect 19978 11704 19984 11716
rect 20036 11704 20042 11756
rect 20073 11747 20131 11753
rect 20073 11713 20085 11747
rect 20119 11744 20131 11747
rect 20254 11744 20260 11756
rect 20119 11716 20260 11744
rect 20119 11713 20131 11716
rect 20073 11707 20131 11713
rect 20254 11704 20260 11716
rect 20312 11704 20318 11756
rect 22002 11704 22008 11756
rect 22060 11744 22066 11756
rect 22940 11753 22968 11784
rect 23474 11772 23480 11784
rect 23532 11772 23538 11824
rect 22925 11747 22983 11753
rect 22925 11744 22937 11747
rect 22060 11716 22937 11744
rect 22060 11704 22066 11716
rect 22925 11713 22937 11716
rect 22971 11713 22983 11747
rect 22925 11707 22983 11713
rect 23192 11747 23250 11753
rect 23192 11713 23204 11747
rect 23238 11744 23250 11747
rect 24780 11744 24808 11843
rect 25222 11840 25228 11852
rect 25280 11840 25286 11892
rect 25774 11840 25780 11892
rect 25832 11880 25838 11892
rect 26329 11883 26387 11889
rect 26329 11880 26341 11883
rect 25832 11852 26341 11880
rect 25832 11840 25838 11852
rect 26329 11849 26341 11852
rect 26375 11849 26387 11883
rect 26329 11843 26387 11849
rect 34606 11840 34612 11892
rect 34664 11880 34670 11892
rect 35161 11883 35219 11889
rect 35161 11880 35173 11883
rect 34664 11852 35173 11880
rect 34664 11840 34670 11852
rect 35161 11849 35173 11852
rect 35207 11849 35219 11883
rect 37458 11880 37464 11892
rect 37419 11852 37464 11880
rect 35161 11843 35219 11849
rect 37458 11840 37464 11852
rect 37516 11840 37522 11892
rect 37826 11880 37832 11892
rect 37787 11852 37832 11880
rect 37826 11840 37832 11852
rect 37884 11840 37890 11892
rect 25958 11812 25964 11824
rect 25919 11784 25964 11812
rect 25958 11772 25964 11784
rect 26016 11772 26022 11824
rect 26050 11772 26056 11824
rect 26108 11812 26114 11824
rect 26161 11815 26219 11821
rect 26161 11812 26173 11815
rect 26108 11784 26173 11812
rect 26108 11772 26114 11784
rect 26161 11781 26173 11784
rect 26207 11781 26219 11815
rect 26161 11775 26219 11781
rect 30644 11815 30702 11821
rect 30644 11781 30656 11815
rect 30690 11812 30702 11815
rect 31110 11812 31116 11824
rect 30690 11784 31116 11812
rect 30690 11781 30702 11784
rect 30644 11775 30702 11781
rect 31110 11772 31116 11784
rect 31168 11772 31174 11824
rect 33042 11812 33048 11824
rect 31726 11784 33048 11812
rect 23238 11716 24808 11744
rect 25133 11747 25191 11753
rect 23238 11713 23250 11716
rect 23192 11707 23250 11713
rect 25133 11713 25145 11747
rect 25179 11713 25191 11747
rect 25133 11707 25191 11713
rect 29273 11747 29331 11753
rect 29273 11713 29285 11747
rect 29319 11744 29331 11747
rect 30098 11744 30104 11756
rect 29319 11716 30104 11744
rect 29319 11713 29331 11716
rect 29273 11707 29331 11713
rect 19812 11648 19932 11676
rect 11698 11608 11704 11620
rect 10428 11580 11704 11608
rect 11698 11568 11704 11580
rect 11756 11568 11762 11620
rect 17678 11568 17684 11620
rect 17736 11608 17742 11620
rect 17865 11611 17923 11617
rect 17865 11608 17877 11611
rect 17736 11580 17877 11608
rect 17736 11568 17742 11580
rect 17865 11577 17877 11580
rect 17911 11608 17923 11611
rect 19904 11608 19932 11648
rect 21726 11608 21732 11620
rect 17911 11580 21732 11608
rect 17911 11577 17923 11580
rect 17865 11571 17923 11577
rect 21726 11568 21732 11580
rect 21784 11568 21790 11620
rect 24305 11611 24363 11617
rect 24305 11577 24317 11611
rect 24351 11608 24363 11611
rect 24762 11608 24768 11620
rect 24351 11580 24768 11608
rect 24351 11577 24363 11580
rect 24305 11571 24363 11577
rect 24762 11568 24768 11580
rect 24820 11608 24826 11620
rect 25148 11608 25176 11707
rect 30098 11704 30104 11716
rect 30156 11704 30162 11756
rect 30374 11744 30380 11756
rect 30335 11716 30380 11744
rect 30374 11704 30380 11716
rect 30432 11704 30438 11756
rect 30466 11704 30472 11756
rect 30524 11744 30530 11756
rect 31726 11744 31754 11784
rect 33042 11772 33048 11784
rect 33100 11772 33106 11824
rect 32306 11744 32312 11756
rect 30524 11716 31754 11744
rect 32267 11716 32312 11744
rect 30524 11704 30530 11716
rect 32306 11704 32312 11716
rect 32364 11704 32370 11756
rect 32858 11744 32864 11756
rect 32819 11716 32864 11744
rect 32858 11704 32864 11716
rect 32916 11704 32922 11756
rect 33134 11744 33140 11756
rect 33095 11716 33140 11744
rect 33134 11704 33140 11716
rect 33192 11704 33198 11756
rect 33781 11747 33839 11753
rect 33781 11713 33793 11747
rect 33827 11744 33839 11747
rect 33870 11744 33876 11756
rect 33827 11716 33876 11744
rect 33827 11713 33839 11716
rect 33781 11707 33839 11713
rect 33870 11704 33876 11716
rect 33928 11704 33934 11756
rect 34698 11704 34704 11756
rect 34756 11744 34762 11756
rect 35069 11747 35127 11753
rect 35069 11744 35081 11747
rect 34756 11716 35081 11744
rect 34756 11704 34762 11716
rect 35069 11713 35081 11716
rect 35115 11713 35127 11747
rect 35894 11744 35900 11756
rect 35855 11716 35900 11744
rect 35069 11707 35127 11713
rect 35894 11704 35900 11716
rect 35952 11704 35958 11756
rect 36541 11747 36599 11753
rect 36541 11713 36553 11747
rect 36587 11744 36599 11747
rect 37844 11744 37872 11840
rect 36587 11716 37872 11744
rect 36587 11713 36599 11716
rect 36541 11707 36599 11713
rect 25409 11679 25467 11685
rect 25409 11645 25421 11679
rect 25455 11645 25467 11679
rect 25409 11639 25467 11645
rect 24820 11580 25176 11608
rect 25424 11608 25452 11639
rect 25774 11636 25780 11688
rect 25832 11676 25838 11688
rect 26142 11676 26148 11688
rect 25832 11648 26148 11676
rect 25832 11636 25838 11648
rect 26142 11636 26148 11648
rect 26200 11636 26206 11688
rect 26234 11636 26240 11688
rect 26292 11676 26298 11688
rect 29365 11679 29423 11685
rect 29365 11676 29377 11679
rect 26292 11648 29377 11676
rect 26292 11636 26298 11648
rect 29365 11645 29377 11648
rect 29411 11645 29423 11679
rect 29365 11639 29423 11645
rect 29457 11679 29515 11685
rect 29457 11645 29469 11679
rect 29503 11676 29515 11679
rect 30484 11676 30512 11704
rect 29503 11648 30512 11676
rect 29503 11645 29515 11648
rect 29457 11639 29515 11645
rect 29472 11608 29500 11639
rect 31478 11636 31484 11688
rect 31536 11676 31542 11688
rect 33045 11679 33103 11685
rect 33045 11676 33057 11679
rect 31536 11648 33057 11676
rect 31536 11636 31542 11648
rect 31772 11617 31800 11648
rect 33045 11645 33057 11648
rect 33091 11645 33103 11679
rect 33505 11679 33563 11685
rect 33505 11676 33517 11679
rect 33045 11639 33103 11645
rect 33428 11648 33517 11676
rect 25424 11580 29500 11608
rect 31757 11611 31815 11617
rect 24820 11568 24826 11580
rect 31757 11577 31769 11611
rect 31803 11608 31815 11611
rect 33428 11608 33456 11648
rect 33505 11645 33517 11648
rect 33551 11645 33563 11679
rect 35802 11676 35808 11688
rect 35763 11648 35808 11676
rect 33505 11639 33563 11645
rect 35802 11636 35808 11648
rect 35860 11636 35866 11688
rect 36265 11679 36323 11685
rect 36265 11645 36277 11679
rect 36311 11645 36323 11679
rect 36265 11639 36323 11645
rect 37921 11679 37979 11685
rect 37921 11645 37933 11679
rect 37967 11645 37979 11679
rect 37921 11639 37979 11645
rect 38105 11679 38163 11685
rect 38105 11645 38117 11679
rect 38151 11676 38163 11679
rect 38194 11676 38200 11688
rect 38151 11648 38200 11676
rect 38151 11645 38163 11648
rect 38105 11639 38163 11645
rect 36170 11608 36176 11620
rect 31803 11580 31837 11608
rect 33428 11580 36176 11608
rect 31803 11577 31815 11580
rect 31757 11571 31815 11577
rect 10318 11500 10324 11552
rect 10376 11540 10382 11552
rect 11238 11540 11244 11552
rect 10376 11512 11244 11540
rect 10376 11500 10382 11512
rect 11238 11500 11244 11512
rect 11296 11540 11302 11552
rect 11974 11540 11980 11552
rect 11296 11512 11980 11540
rect 11296 11500 11302 11512
rect 11974 11500 11980 11512
rect 12032 11540 12038 11552
rect 12713 11543 12771 11549
rect 12713 11540 12725 11543
rect 12032 11512 12725 11540
rect 12032 11500 12038 11512
rect 12713 11509 12725 11512
rect 12759 11509 12771 11543
rect 26142 11540 26148 11552
rect 26103 11512 26148 11540
rect 12713 11503 12771 11509
rect 26142 11500 26148 11512
rect 26200 11500 26206 11552
rect 28905 11543 28963 11549
rect 28905 11509 28917 11543
rect 28951 11540 28963 11543
rect 28994 11540 29000 11552
rect 28951 11512 29000 11540
rect 28951 11509 28963 11512
rect 28905 11503 28963 11509
rect 28994 11500 29000 11512
rect 29052 11500 29058 11552
rect 31846 11500 31852 11552
rect 31904 11540 31910 11552
rect 33428 11540 33456 11580
rect 36170 11568 36176 11580
rect 36228 11608 36234 11620
rect 36280 11608 36308 11639
rect 36228 11580 36308 11608
rect 36228 11568 36234 11580
rect 31904 11512 33456 11540
rect 31904 11500 31910 11512
rect 35710 11500 35716 11552
rect 35768 11540 35774 11552
rect 37936 11540 37964 11639
rect 38194 11636 38200 11648
rect 38252 11636 38258 11688
rect 35768 11512 37964 11540
rect 35768 11500 35774 11512
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 10778 11296 10784 11348
rect 10836 11336 10842 11348
rect 10965 11339 11023 11345
rect 10965 11336 10977 11339
rect 10836 11308 10977 11336
rect 10836 11296 10842 11308
rect 10965 11305 10977 11308
rect 11011 11305 11023 11339
rect 10965 11299 11023 11305
rect 11054 11296 11060 11348
rect 11112 11336 11118 11348
rect 12253 11339 12311 11345
rect 12253 11336 12265 11339
rect 11112 11308 12265 11336
rect 11112 11296 11118 11308
rect 12253 11305 12265 11308
rect 12299 11305 12311 11339
rect 12253 11299 12311 11305
rect 14826 11296 14832 11348
rect 14884 11336 14890 11348
rect 15013 11339 15071 11345
rect 15013 11336 15025 11339
rect 14884 11308 15025 11336
rect 14884 11296 14890 11308
rect 15013 11305 15025 11308
rect 15059 11305 15071 11339
rect 15013 11299 15071 11305
rect 19705 11339 19763 11345
rect 19705 11305 19717 11339
rect 19751 11336 19763 11339
rect 19978 11336 19984 11348
rect 19751 11308 19984 11336
rect 19751 11305 19763 11308
rect 19705 11299 19763 11305
rect 19978 11296 19984 11308
rect 20036 11296 20042 11348
rect 21450 11296 21456 11348
rect 21508 11336 21514 11348
rect 21637 11339 21695 11345
rect 21637 11336 21649 11339
rect 21508 11308 21649 11336
rect 21508 11296 21514 11308
rect 21637 11305 21649 11308
rect 21683 11305 21695 11339
rect 30834 11336 30840 11348
rect 21637 11299 21695 11305
rect 27908 11308 30840 11336
rect 15746 11268 15752 11280
rect 12406 11240 15752 11268
rect 10137 11203 10195 11209
rect 10137 11169 10149 11203
rect 10183 11200 10195 11203
rect 12406 11200 12434 11240
rect 15746 11228 15752 11240
rect 15804 11228 15810 11280
rect 17770 11268 17776 11280
rect 16408 11240 17776 11268
rect 10183 11172 12434 11200
rect 10183 11169 10195 11172
rect 10137 11163 10195 11169
rect 10045 11135 10103 11141
rect 10045 11101 10057 11135
rect 10091 11101 10103 11135
rect 10318 11132 10324 11144
rect 10279 11104 10324 11132
rect 10045 11095 10103 11101
rect 10060 11064 10088 11095
rect 10318 11092 10324 11104
rect 10376 11092 10382 11144
rect 10413 11135 10471 11141
rect 10413 11101 10425 11135
rect 10459 11132 10471 11135
rect 11054 11132 11060 11144
rect 10459 11104 11060 11132
rect 10459 11101 10471 11104
rect 10413 11095 10471 11101
rect 11054 11092 11060 11104
rect 11112 11132 11118 11144
rect 11149 11135 11207 11141
rect 11149 11132 11161 11135
rect 11112 11104 11161 11132
rect 11112 11092 11118 11104
rect 11149 11101 11161 11104
rect 11195 11101 11207 11135
rect 11149 11095 11207 11101
rect 11238 11092 11244 11144
rect 11296 11132 11302 11144
rect 11532 11141 11560 11172
rect 11425 11135 11483 11141
rect 11296 11104 11341 11132
rect 11296 11092 11302 11104
rect 11425 11101 11437 11135
rect 11471 11101 11483 11135
rect 11425 11095 11483 11101
rect 11517 11135 11575 11141
rect 11517 11101 11529 11135
rect 11563 11101 11575 11135
rect 11517 11095 11575 11101
rect 12253 11135 12311 11141
rect 12253 11101 12265 11135
rect 12299 11132 12311 11135
rect 12342 11132 12348 11144
rect 12299 11104 12348 11132
rect 12299 11101 12311 11104
rect 12253 11095 12311 11101
rect 11440 11064 11468 11095
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 12529 11135 12587 11141
rect 12529 11101 12541 11135
rect 12575 11132 12587 11135
rect 12618 11132 12624 11144
rect 12575 11104 12624 11132
rect 12575 11101 12587 11104
rect 12529 11095 12587 11101
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 13998 11092 14004 11144
rect 14056 11132 14062 11144
rect 15013 11135 15071 11141
rect 15013 11132 15025 11135
rect 14056 11104 15025 11132
rect 14056 11092 14062 11104
rect 15013 11101 15025 11104
rect 15059 11101 15071 11135
rect 15013 11095 15071 11101
rect 15289 11135 15347 11141
rect 15289 11101 15301 11135
rect 15335 11132 15347 11135
rect 15378 11132 15384 11144
rect 15335 11104 15384 11132
rect 15335 11101 15347 11104
rect 15289 11095 15347 11101
rect 15378 11092 15384 11104
rect 15436 11092 15442 11144
rect 15197 11067 15255 11073
rect 10060 11036 15153 11064
rect 10502 10996 10508 11008
rect 10463 10968 10508 10996
rect 10502 10956 10508 10968
rect 10560 10956 10566 11008
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 13354 10996 13360 11008
rect 12492 10968 13360 10996
rect 12492 10956 12498 10968
rect 13354 10956 13360 10968
rect 13412 10956 13418 11008
rect 15125 10996 15153 11036
rect 15197 11033 15209 11067
rect 15243 11064 15255 11067
rect 16408 11064 16436 11240
rect 17770 11228 17776 11240
rect 17828 11228 17834 11280
rect 18046 11268 18052 11280
rect 18007 11240 18052 11268
rect 18046 11228 18052 11240
rect 18104 11268 18110 11280
rect 18598 11268 18604 11280
rect 18104 11240 18604 11268
rect 18104 11228 18110 11240
rect 18598 11228 18604 11240
rect 18656 11228 18662 11280
rect 19334 11200 19340 11212
rect 16500 11172 19340 11200
rect 16500 11141 16528 11172
rect 19334 11160 19340 11172
rect 19392 11160 19398 11212
rect 20162 11200 20168 11212
rect 19628 11172 20168 11200
rect 16485 11135 16543 11141
rect 16485 11101 16497 11135
rect 16531 11101 16543 11135
rect 16485 11095 16543 11101
rect 16669 11135 16727 11141
rect 16669 11101 16681 11135
rect 16715 11132 16727 11135
rect 17129 11135 17187 11141
rect 16715 11104 16988 11132
rect 16715 11101 16727 11104
rect 16669 11095 16727 11101
rect 15243 11036 16436 11064
rect 16577 11067 16635 11073
rect 15243 11033 15255 11036
rect 15197 11027 15255 11033
rect 16577 11033 16589 11067
rect 16623 11064 16635 11067
rect 16850 11064 16856 11076
rect 16623 11036 16856 11064
rect 16623 11033 16635 11036
rect 16577 11027 16635 11033
rect 16850 11024 16856 11036
rect 16908 11024 16914 11076
rect 16960 11008 16988 11104
rect 17129 11101 17141 11135
rect 17175 11132 17187 11135
rect 17586 11132 17592 11144
rect 17175 11104 17592 11132
rect 17175 11101 17187 11104
rect 17129 11095 17187 11101
rect 17586 11092 17592 11104
rect 17644 11092 17650 11144
rect 19628 11141 19656 11172
rect 20162 11160 20168 11172
rect 20220 11160 20226 11212
rect 22462 11200 22468 11212
rect 21560 11172 22468 11200
rect 19613 11135 19671 11141
rect 19613 11101 19625 11135
rect 19659 11101 19671 11135
rect 19613 11095 19671 11101
rect 19797 11135 19855 11141
rect 19797 11101 19809 11135
rect 19843 11132 19855 11135
rect 20438 11132 20444 11144
rect 19843 11104 20444 11132
rect 19843 11101 19855 11104
rect 19797 11095 19855 11101
rect 17773 11067 17831 11073
rect 17773 11033 17785 11067
rect 17819 11064 17831 11067
rect 18506 11064 18512 11076
rect 17819 11036 18512 11064
rect 17819 11033 17831 11036
rect 17773 11027 17831 11033
rect 18506 11024 18512 11036
rect 18564 11024 18570 11076
rect 18966 11024 18972 11076
rect 19024 11064 19030 11076
rect 19812 11064 19840 11095
rect 20438 11092 20444 11104
rect 20496 11092 20502 11144
rect 21560 11141 21588 11172
rect 22462 11160 22468 11172
rect 22520 11200 22526 11212
rect 22922 11200 22928 11212
rect 22520 11172 22928 11200
rect 22520 11160 22526 11172
rect 22922 11160 22928 11172
rect 22980 11160 22986 11212
rect 25222 11160 25228 11212
rect 25280 11200 25286 11212
rect 25409 11203 25467 11209
rect 25409 11200 25421 11203
rect 25280 11172 25421 11200
rect 25280 11160 25286 11172
rect 25409 11169 25421 11172
rect 25455 11169 25467 11203
rect 25409 11163 25467 11169
rect 25593 11203 25651 11209
rect 25593 11169 25605 11203
rect 25639 11200 25651 11203
rect 25639 11172 26832 11200
rect 25639 11169 25651 11172
rect 25593 11163 25651 11169
rect 21545 11135 21603 11141
rect 21545 11101 21557 11135
rect 21591 11101 21603 11135
rect 21545 11095 21603 11101
rect 21634 11092 21640 11144
rect 21692 11132 21698 11144
rect 21821 11135 21879 11141
rect 21821 11132 21833 11135
rect 21692 11104 21833 11132
rect 21692 11092 21698 11104
rect 21821 11101 21833 11104
rect 21867 11101 21879 11135
rect 26694 11132 26700 11144
rect 26655 11104 26700 11132
rect 21821 11095 21879 11101
rect 26694 11092 26700 11104
rect 26752 11092 26758 11144
rect 26804 11132 26832 11172
rect 27246 11132 27252 11144
rect 26804 11104 27252 11132
rect 27246 11092 27252 11104
rect 27304 11132 27310 11144
rect 27908 11132 27936 11308
rect 30834 11296 30840 11308
rect 30892 11336 30898 11348
rect 34422 11336 34428 11348
rect 30892 11308 34428 11336
rect 30892 11296 30898 11308
rect 34422 11296 34428 11308
rect 34480 11296 34486 11348
rect 35802 11296 35808 11348
rect 35860 11336 35866 11348
rect 36265 11339 36323 11345
rect 36265 11336 36277 11339
rect 35860 11308 36277 11336
rect 35860 11296 35866 11308
rect 36265 11305 36277 11308
rect 36311 11305 36323 11339
rect 36265 11299 36323 11305
rect 28902 11228 28908 11280
rect 28960 11268 28966 11280
rect 29825 11271 29883 11277
rect 29825 11268 29837 11271
rect 28960 11240 29837 11268
rect 28960 11228 28966 11240
rect 29825 11237 29837 11240
rect 29871 11237 29883 11271
rect 33134 11268 33140 11280
rect 29825 11231 29883 11237
rect 30576 11240 33140 11268
rect 30469 11203 30527 11209
rect 30469 11200 30481 11203
rect 27304 11104 27936 11132
rect 28736 11172 30481 11200
rect 27304 11092 27310 11104
rect 19024 11036 19840 11064
rect 25317 11067 25375 11073
rect 19024 11024 19030 11036
rect 25317 11033 25329 11067
rect 25363 11064 25375 11067
rect 25958 11064 25964 11076
rect 25363 11036 25964 11064
rect 25363 11033 25375 11036
rect 25317 11027 25375 11033
rect 25958 11024 25964 11036
rect 26016 11024 26022 11076
rect 26964 11067 27022 11073
rect 26964 11033 26976 11067
rect 27010 11064 27022 11067
rect 27154 11064 27160 11076
rect 27010 11036 27160 11064
rect 27010 11033 27022 11036
rect 26964 11027 27022 11033
rect 27154 11024 27160 11036
rect 27212 11024 27218 11076
rect 15286 10996 15292 11008
rect 15125 10968 15292 10996
rect 15286 10956 15292 10968
rect 15344 10996 15350 11008
rect 16942 10996 16948 11008
rect 15344 10968 16948 10996
rect 15344 10956 15350 10968
rect 16942 10956 16948 10968
rect 17000 10956 17006 11008
rect 17218 10996 17224 11008
rect 17179 10968 17224 10996
rect 17218 10956 17224 10968
rect 17276 10956 17282 11008
rect 18230 10996 18236 11008
rect 18191 10968 18236 10996
rect 18230 10956 18236 10968
rect 18288 10956 18294 11008
rect 22002 10956 22008 11008
rect 22060 10996 22066 11008
rect 22097 10999 22155 11005
rect 22097 10996 22109 10999
rect 22060 10968 22109 10996
rect 22060 10956 22066 10968
rect 22097 10965 22109 10968
rect 22143 10965 22155 10999
rect 22097 10959 22155 10965
rect 24854 10956 24860 11008
rect 24912 10996 24918 11008
rect 24949 10999 25007 11005
rect 24949 10996 24961 10999
rect 24912 10968 24961 10996
rect 24912 10956 24918 10968
rect 24949 10965 24961 10968
rect 24995 10965 25007 10999
rect 28074 10996 28080 11008
rect 27987 10968 28080 10996
rect 24949 10959 25007 10965
rect 28074 10956 28080 10968
rect 28132 10996 28138 11008
rect 28736 10996 28764 11172
rect 30469 11169 30481 11172
rect 30515 11169 30527 11203
rect 30469 11163 30527 11169
rect 29178 11092 29184 11144
rect 29236 11132 29242 11144
rect 29733 11135 29791 11141
rect 29733 11132 29745 11135
rect 29236 11104 29745 11132
rect 29236 11092 29242 11104
rect 29733 11101 29745 11104
rect 29779 11101 29791 11135
rect 29733 11095 29791 11101
rect 30282 11092 30288 11144
rect 30340 11132 30346 11144
rect 30576 11141 30604 11240
rect 33134 11228 33140 11240
rect 33192 11268 33198 11280
rect 33594 11268 33600 11280
rect 33192 11240 33600 11268
rect 33192 11228 33198 11240
rect 33594 11228 33600 11240
rect 33652 11228 33658 11280
rect 32490 11160 32496 11212
rect 32548 11200 32554 11212
rect 32950 11200 32956 11212
rect 32548 11172 32956 11200
rect 32548 11160 32554 11172
rect 32950 11160 32956 11172
rect 33008 11200 33014 11212
rect 33873 11203 33931 11209
rect 33873 11200 33885 11203
rect 33008 11172 33885 11200
rect 33008 11160 33014 11172
rect 33873 11169 33885 11172
rect 33919 11200 33931 11203
rect 34885 11203 34943 11209
rect 34885 11200 34897 11203
rect 33919 11172 34897 11200
rect 33919 11169 33931 11172
rect 33873 11163 33931 11169
rect 34885 11169 34897 11172
rect 34931 11169 34943 11203
rect 34885 11163 34943 11169
rect 30561 11135 30619 11141
rect 30561 11132 30573 11135
rect 30340 11104 30573 11132
rect 30340 11092 30346 11104
rect 30561 11101 30573 11104
rect 30607 11101 30619 11135
rect 30561 11095 30619 11101
rect 31021 11135 31079 11141
rect 31021 11101 31033 11135
rect 31067 11101 31079 11135
rect 31386 11132 31392 11144
rect 31347 11104 31392 11132
rect 31021 11095 31079 11101
rect 30098 11024 30104 11076
rect 30156 11064 30162 11076
rect 31036 11064 31064 11095
rect 31386 11092 31392 11104
rect 31444 11092 31450 11144
rect 34900 11132 34928 11163
rect 36725 11135 36783 11141
rect 36725 11132 36737 11135
rect 34900 11104 36737 11132
rect 36725 11101 36737 11104
rect 36771 11101 36783 11135
rect 36725 11095 36783 11101
rect 30156 11036 31064 11064
rect 33137 11067 33195 11073
rect 30156 11024 30162 11036
rect 33137 11033 33149 11067
rect 33183 11064 33195 11067
rect 33226 11064 33232 11076
rect 33183 11036 33232 11064
rect 33183 11033 33195 11036
rect 33137 11027 33195 11033
rect 33226 11024 33232 11036
rect 33284 11024 33290 11076
rect 34790 11024 34796 11076
rect 34848 11064 34854 11076
rect 35130 11067 35188 11073
rect 35130 11064 35142 11067
rect 34848 11036 35142 11064
rect 34848 11024 34854 11036
rect 35130 11033 35142 11036
rect 35176 11033 35188 11067
rect 35130 11027 35188 11033
rect 36992 11067 37050 11073
rect 36992 11033 37004 11067
rect 37038 11064 37050 11067
rect 37458 11064 37464 11076
rect 37038 11036 37464 11064
rect 37038 11033 37050 11036
rect 36992 11027 37050 11033
rect 37458 11024 37464 11036
rect 37516 11024 37522 11076
rect 28132 10968 28764 10996
rect 28132 10956 28138 10968
rect 37826 10956 37832 11008
rect 37884 10996 37890 11008
rect 38105 10999 38163 11005
rect 38105 10996 38117 10999
rect 37884 10968 38117 10996
rect 37884 10956 37890 10968
rect 38105 10965 38117 10968
rect 38151 10965 38163 10999
rect 38105 10959 38163 10965
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 17218 10752 17224 10804
rect 17276 10792 17282 10804
rect 17773 10795 17831 10801
rect 17773 10792 17785 10795
rect 17276 10764 17785 10792
rect 17276 10752 17282 10764
rect 17773 10761 17785 10764
rect 17819 10761 17831 10795
rect 18506 10792 18512 10804
rect 18467 10764 18512 10792
rect 17773 10755 17831 10761
rect 18506 10752 18512 10764
rect 18564 10792 18570 10804
rect 21085 10795 21143 10801
rect 21085 10792 21097 10795
rect 18564 10764 21097 10792
rect 18564 10752 18570 10764
rect 21085 10761 21097 10764
rect 21131 10792 21143 10795
rect 24946 10792 24952 10804
rect 21131 10764 24952 10792
rect 21131 10761 21143 10764
rect 21085 10755 21143 10761
rect 24946 10752 24952 10764
rect 25004 10752 25010 10804
rect 25958 10792 25964 10804
rect 25919 10764 25964 10792
rect 25958 10752 25964 10764
rect 26016 10752 26022 10804
rect 27154 10792 27160 10804
rect 27115 10764 27160 10792
rect 27154 10752 27160 10764
rect 27212 10752 27218 10804
rect 27525 10795 27583 10801
rect 27525 10761 27537 10795
rect 27571 10792 27583 10795
rect 28074 10792 28080 10804
rect 27571 10764 28080 10792
rect 27571 10761 27583 10764
rect 27525 10755 27583 10761
rect 28074 10752 28080 10764
rect 28132 10752 28138 10804
rect 30098 10792 30104 10804
rect 30059 10764 30104 10792
rect 30098 10752 30104 10764
rect 30156 10752 30162 10804
rect 37458 10792 37464 10804
rect 37419 10764 37464 10792
rect 37458 10752 37464 10764
rect 37516 10752 37522 10804
rect 17678 10724 17684 10736
rect 17639 10696 17684 10724
rect 17678 10684 17684 10696
rect 17736 10684 17742 10736
rect 21450 10684 21456 10736
rect 21508 10724 21514 10736
rect 22281 10727 22339 10733
rect 22281 10724 22293 10727
rect 21508 10696 22293 10724
rect 21508 10684 21514 10696
rect 22281 10693 22293 10696
rect 22327 10693 22339 10727
rect 26694 10724 26700 10736
rect 22281 10687 22339 10693
rect 24596 10696 26700 10724
rect 11790 10656 11796 10668
rect 11751 10628 11796 10656
rect 11790 10616 11796 10628
rect 11848 10616 11854 10668
rect 11974 10656 11980 10668
rect 11935 10628 11980 10656
rect 11974 10616 11980 10628
rect 12032 10616 12038 10668
rect 13170 10656 13176 10668
rect 13131 10628 13176 10656
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 13354 10616 13360 10668
rect 13412 10656 13418 10668
rect 15381 10659 15439 10665
rect 15381 10656 15393 10659
rect 13412 10628 15393 10656
rect 13412 10616 13418 10628
rect 15381 10625 15393 10628
rect 15427 10656 15439 10659
rect 15470 10656 15476 10668
rect 15427 10628 15476 10656
rect 15427 10625 15439 10628
rect 15381 10619 15439 10625
rect 15470 10616 15476 10628
rect 15528 10616 15534 10668
rect 15565 10659 15623 10665
rect 15565 10625 15577 10659
rect 15611 10656 15623 10659
rect 15654 10656 15660 10668
rect 15611 10628 15660 10656
rect 15611 10625 15623 10628
rect 15565 10619 15623 10625
rect 15654 10616 15660 10628
rect 15712 10616 15718 10668
rect 18046 10616 18052 10668
rect 18104 10656 18110 10668
rect 18877 10659 18935 10665
rect 18877 10656 18889 10659
rect 18104 10628 18889 10656
rect 18104 10616 18110 10628
rect 18877 10625 18889 10628
rect 18923 10625 18935 10659
rect 18877 10619 18935 10625
rect 20806 10616 20812 10668
rect 20864 10656 20870 10668
rect 22002 10656 22008 10668
rect 20864 10628 21312 10656
rect 21963 10628 22008 10656
rect 20864 10616 20870 10628
rect 17865 10591 17923 10597
rect 17865 10557 17877 10591
rect 17911 10588 17923 10591
rect 18230 10588 18236 10600
rect 17911 10560 18236 10588
rect 17911 10557 17923 10560
rect 17865 10551 17923 10557
rect 18230 10548 18236 10560
rect 18288 10548 18294 10600
rect 21284 10597 21312 10628
rect 22002 10616 22008 10628
rect 22060 10616 22066 10668
rect 22186 10656 22192 10668
rect 22147 10628 22192 10656
rect 22186 10616 22192 10628
rect 22244 10616 22250 10668
rect 22370 10616 22376 10668
rect 22428 10656 22434 10668
rect 22428 10628 22473 10656
rect 22428 10616 22434 10628
rect 18969 10591 19027 10597
rect 18969 10557 18981 10591
rect 19015 10588 19027 10591
rect 21177 10591 21235 10597
rect 19015 10560 20852 10588
rect 19015 10557 19027 10560
rect 18969 10551 19027 10557
rect 17770 10480 17776 10532
rect 17828 10520 17834 10532
rect 18984 10520 19012 10551
rect 17828 10492 19012 10520
rect 17828 10480 17834 10492
rect 11238 10412 11244 10464
rect 11296 10452 11302 10464
rect 11885 10455 11943 10461
rect 11885 10452 11897 10455
rect 11296 10424 11897 10452
rect 11296 10412 11302 10424
rect 11885 10421 11897 10424
rect 11931 10421 11943 10455
rect 13538 10452 13544 10464
rect 13499 10424 13544 10452
rect 11885 10415 11943 10421
rect 13538 10412 13544 10424
rect 13596 10412 13602 10464
rect 15378 10452 15384 10464
rect 15339 10424 15384 10452
rect 15378 10412 15384 10424
rect 15436 10412 15442 10464
rect 17313 10455 17371 10461
rect 17313 10421 17325 10455
rect 17359 10452 17371 10455
rect 17402 10452 17408 10464
rect 17359 10424 17408 10452
rect 17359 10421 17371 10424
rect 17313 10415 17371 10421
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 17494 10412 17500 10464
rect 17552 10452 17558 10464
rect 19153 10455 19211 10461
rect 19153 10452 19165 10455
rect 17552 10424 19165 10452
rect 17552 10412 17558 10424
rect 19153 10421 19165 10424
rect 19199 10421 19211 10455
rect 20714 10452 20720 10464
rect 20675 10424 20720 10452
rect 19153 10415 19211 10421
rect 20714 10412 20720 10424
rect 20772 10412 20778 10464
rect 20824 10452 20852 10560
rect 21177 10557 21189 10591
rect 21223 10557 21235 10591
rect 21177 10551 21235 10557
rect 21269 10591 21327 10597
rect 21269 10557 21281 10591
rect 21315 10557 21327 10591
rect 21269 10551 21327 10557
rect 21192 10520 21220 10551
rect 23474 10548 23480 10600
rect 23532 10588 23538 10600
rect 24596 10597 24624 10696
rect 26694 10684 26700 10696
rect 26752 10724 26758 10736
rect 28994 10733 29000 10736
rect 28988 10724 29000 10733
rect 26752 10696 28764 10724
rect 28955 10696 29000 10724
rect 26752 10684 26758 10696
rect 24854 10665 24860 10668
rect 24848 10656 24860 10665
rect 24815 10628 24860 10656
rect 24848 10619 24860 10628
rect 24854 10616 24860 10619
rect 24912 10616 24918 10668
rect 26234 10616 26240 10668
rect 26292 10656 26298 10668
rect 27522 10656 27528 10668
rect 26292 10628 27528 10656
rect 26292 10616 26298 10628
rect 27522 10616 27528 10628
rect 27580 10656 27586 10668
rect 28736 10665 28764 10696
rect 28988 10687 29000 10696
rect 28994 10684 29000 10687
rect 29052 10684 29058 10736
rect 37921 10727 37979 10733
rect 37921 10724 37933 10727
rect 34348 10696 37933 10724
rect 27617 10659 27675 10665
rect 27617 10656 27629 10659
rect 27580 10628 27629 10656
rect 27580 10616 27586 10628
rect 27617 10625 27629 10628
rect 27663 10625 27675 10659
rect 27617 10619 27675 10625
rect 28721 10659 28779 10665
rect 28721 10625 28733 10659
rect 28767 10625 28779 10659
rect 34238 10656 34244 10668
rect 34199 10628 34244 10656
rect 28721 10619 28779 10625
rect 34238 10616 34244 10628
rect 34296 10616 34302 10668
rect 24581 10591 24639 10597
rect 24581 10588 24593 10591
rect 23532 10560 24593 10588
rect 23532 10548 23538 10560
rect 24581 10557 24593 10560
rect 24627 10557 24639 10591
rect 24581 10551 24639 10557
rect 27246 10548 27252 10600
rect 27304 10588 27310 10600
rect 27709 10591 27767 10597
rect 27709 10588 27721 10591
rect 27304 10560 27721 10588
rect 27304 10548 27310 10560
rect 27709 10557 27721 10560
rect 27755 10557 27767 10591
rect 33318 10588 33324 10600
rect 27709 10551 27767 10557
rect 31726 10560 33324 10588
rect 22557 10523 22615 10529
rect 22557 10520 22569 10523
rect 21192 10492 22569 10520
rect 22557 10489 22569 10492
rect 22603 10489 22615 10523
rect 22557 10483 22615 10489
rect 22646 10452 22652 10464
rect 20824 10424 22652 10452
rect 22646 10412 22652 10424
rect 22704 10412 22710 10464
rect 25682 10412 25688 10464
rect 25740 10452 25746 10464
rect 31726 10452 31754 10560
rect 33318 10548 33324 10560
rect 33376 10588 33382 10600
rect 34348 10597 34376 10696
rect 37921 10693 37933 10696
rect 37967 10724 37979 10727
rect 38010 10724 38016 10736
rect 37967 10696 38016 10724
rect 37967 10693 37979 10696
rect 37921 10687 37979 10693
rect 38010 10684 38016 10696
rect 38068 10684 38074 10736
rect 37366 10616 37372 10668
rect 37424 10656 37430 10668
rect 37826 10656 37832 10668
rect 37424 10628 37832 10656
rect 37424 10616 37430 10628
rect 37826 10616 37832 10628
rect 37884 10616 37890 10668
rect 34333 10591 34391 10597
rect 34333 10588 34345 10591
rect 33376 10560 34345 10588
rect 33376 10548 33382 10560
rect 34333 10557 34345 10560
rect 34379 10557 34391 10591
rect 34333 10551 34391 10557
rect 34422 10548 34428 10600
rect 34480 10588 34486 10600
rect 38105 10591 38163 10597
rect 34480 10560 34525 10588
rect 34480 10548 34486 10560
rect 38105 10557 38117 10591
rect 38151 10588 38163 10591
rect 38194 10588 38200 10600
rect 38151 10560 38200 10588
rect 38151 10557 38163 10560
rect 38105 10551 38163 10557
rect 38194 10548 38200 10560
rect 38252 10548 38258 10600
rect 25740 10424 31754 10452
rect 25740 10412 25746 10424
rect 33502 10412 33508 10464
rect 33560 10452 33566 10464
rect 33873 10455 33931 10461
rect 33873 10452 33885 10455
rect 33560 10424 33885 10452
rect 33560 10412 33566 10424
rect 33873 10421 33885 10424
rect 33919 10421 33931 10455
rect 33873 10415 33931 10421
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 10686 10248 10692 10260
rect 10647 10220 10692 10248
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 12526 10208 12532 10260
rect 12584 10248 12590 10260
rect 12894 10248 12900 10260
rect 12584 10220 12900 10248
rect 12584 10208 12590 10220
rect 12894 10208 12900 10220
rect 12952 10248 12958 10260
rect 13173 10251 13231 10257
rect 13173 10248 13185 10251
rect 12952 10220 13185 10248
rect 12952 10208 12958 10220
rect 13173 10217 13185 10220
rect 13219 10217 13231 10251
rect 13173 10211 13231 10217
rect 13354 10208 13360 10260
rect 13412 10248 13418 10260
rect 20530 10248 20536 10260
rect 13412 10220 20536 10248
rect 13412 10208 13418 10220
rect 20530 10208 20536 10220
rect 20588 10208 20594 10260
rect 21913 10251 21971 10257
rect 21913 10217 21925 10251
rect 21959 10248 21971 10251
rect 22186 10248 22192 10260
rect 21959 10220 22192 10248
rect 21959 10217 21971 10220
rect 21913 10211 21971 10217
rect 22186 10208 22192 10220
rect 22244 10208 22250 10260
rect 24854 10248 24860 10260
rect 24815 10220 24860 10248
rect 24854 10208 24860 10220
rect 24912 10208 24918 10260
rect 24949 10251 25007 10257
rect 24949 10217 24961 10251
rect 24995 10248 25007 10251
rect 25866 10248 25872 10260
rect 24995 10220 25872 10248
rect 24995 10217 25007 10220
rect 24949 10211 25007 10217
rect 25866 10208 25872 10220
rect 25924 10208 25930 10260
rect 31849 10251 31907 10257
rect 31849 10217 31861 10251
rect 31895 10248 31907 10251
rect 32306 10248 32312 10260
rect 31895 10220 32312 10248
rect 31895 10217 31907 10220
rect 31849 10211 31907 10217
rect 32306 10208 32312 10220
rect 32364 10208 32370 10260
rect 14826 10140 14832 10192
rect 14884 10180 14890 10192
rect 17221 10183 17279 10189
rect 17221 10180 17233 10183
rect 14884 10152 17233 10180
rect 14884 10140 14890 10152
rect 17221 10149 17233 10152
rect 17267 10149 17279 10183
rect 17221 10143 17279 10149
rect 21726 10140 21732 10192
rect 21784 10140 21790 10192
rect 21821 10183 21879 10189
rect 21821 10149 21833 10183
rect 21867 10180 21879 10183
rect 22370 10180 22376 10192
rect 21867 10152 22376 10180
rect 21867 10149 21879 10152
rect 21821 10143 21879 10149
rect 22370 10140 22376 10152
rect 22428 10180 22434 10192
rect 22557 10183 22615 10189
rect 22557 10180 22569 10183
rect 22428 10152 22569 10180
rect 22428 10140 22434 10152
rect 22557 10149 22569 10152
rect 22603 10149 22615 10183
rect 22557 10143 22615 10149
rect 34238 10140 34244 10192
rect 34296 10180 34302 10192
rect 34333 10183 34391 10189
rect 34333 10180 34345 10183
rect 34296 10152 34345 10180
rect 34296 10140 34302 10152
rect 34333 10149 34345 10152
rect 34379 10149 34391 10183
rect 34333 10143 34391 10149
rect 7926 10072 7932 10124
rect 7984 10112 7990 10124
rect 9125 10115 9183 10121
rect 9125 10112 9137 10115
rect 7984 10084 9137 10112
rect 7984 10072 7990 10084
rect 9125 10081 9137 10084
rect 9171 10081 9183 10115
rect 13262 10112 13268 10124
rect 13223 10084 13268 10112
rect 9125 10075 9183 10081
rect 13262 10072 13268 10084
rect 13320 10112 13326 10124
rect 14458 10112 14464 10124
rect 13320 10084 14464 10112
rect 13320 10072 13326 10084
rect 14458 10072 14464 10084
rect 14516 10112 14522 10124
rect 15657 10115 15715 10121
rect 14516 10084 15240 10112
rect 14516 10072 14522 10084
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10044 9459 10047
rect 10870 10044 10876 10056
rect 9447 10016 10876 10044
rect 9447 10013 9459 10016
rect 9401 10007 9459 10013
rect 10870 10004 10876 10016
rect 10928 10004 10934 10056
rect 11238 10044 11244 10056
rect 11199 10016 11244 10044
rect 11238 10004 11244 10016
rect 11296 10004 11302 10056
rect 11517 10047 11575 10053
rect 11517 10013 11529 10047
rect 11563 10044 11575 10047
rect 13170 10044 13176 10056
rect 11563 10016 12434 10044
rect 13083 10016 13176 10044
rect 11563 10013 11575 10016
rect 11517 10007 11575 10013
rect 11422 9976 11428 9988
rect 11383 9948 11428 9976
rect 11422 9936 11428 9948
rect 11480 9936 11486 9988
rect 12406 9920 12434 10016
rect 13170 10004 13176 10016
rect 13228 10004 13234 10056
rect 13188 9976 13216 10004
rect 15212 9976 15240 10084
rect 15657 10081 15669 10115
rect 15703 10112 15715 10115
rect 20346 10112 20352 10124
rect 15703 10084 20352 10112
rect 15703 10081 15715 10084
rect 15657 10075 15715 10081
rect 20346 10072 20352 10084
rect 20404 10072 20410 10124
rect 21744 10112 21772 10140
rect 22005 10115 22063 10121
rect 22005 10112 22017 10115
rect 21744 10084 22017 10112
rect 22005 10081 22017 10084
rect 22051 10081 22063 10115
rect 22005 10075 22063 10081
rect 25041 10115 25099 10121
rect 25041 10081 25053 10115
rect 25087 10112 25099 10115
rect 26326 10112 26332 10124
rect 25087 10084 26332 10112
rect 25087 10081 25099 10084
rect 25041 10075 25099 10081
rect 26326 10072 26332 10084
rect 26384 10072 26390 10124
rect 26694 10072 26700 10124
rect 26752 10112 26758 10124
rect 26881 10115 26939 10121
rect 26881 10112 26893 10115
rect 26752 10084 26893 10112
rect 26752 10072 26758 10084
rect 26881 10081 26893 10084
rect 26927 10081 26939 10115
rect 32950 10112 32956 10124
rect 32911 10084 32956 10112
rect 26881 10075 26939 10081
rect 32950 10072 32956 10084
rect 33008 10072 33014 10124
rect 34348 10112 34376 10143
rect 34514 10140 34520 10192
rect 34572 10180 34578 10192
rect 35069 10183 35127 10189
rect 35069 10180 35081 10183
rect 34572 10152 35081 10180
rect 34572 10140 34578 10152
rect 35069 10149 35081 10152
rect 35115 10149 35127 10183
rect 35069 10143 35127 10149
rect 35713 10115 35771 10121
rect 35713 10112 35725 10115
rect 34348 10084 35725 10112
rect 35713 10081 35725 10084
rect 35759 10081 35771 10115
rect 36170 10112 36176 10124
rect 36131 10084 36176 10112
rect 35713 10075 35771 10081
rect 36170 10072 36176 10084
rect 36228 10072 36234 10124
rect 37366 10112 37372 10124
rect 36464 10084 37372 10112
rect 15378 10044 15384 10056
rect 15339 10016 15384 10044
rect 15378 10004 15384 10016
rect 15436 10044 15442 10056
rect 16393 10047 16451 10053
rect 16393 10044 16405 10047
rect 15436 10016 16405 10044
rect 15436 10004 15442 10016
rect 16393 10013 16405 10016
rect 16439 10013 16451 10047
rect 16758 10044 16764 10056
rect 16719 10016 16764 10044
rect 16393 10007 16451 10013
rect 16758 10004 16764 10016
rect 16816 10004 16822 10056
rect 17402 10044 17408 10056
rect 17363 10016 17408 10044
rect 17402 10004 17408 10016
rect 17460 10004 17466 10056
rect 18690 10044 18696 10056
rect 18651 10016 18696 10044
rect 18690 10004 18696 10016
rect 18748 10004 18754 10056
rect 18877 10047 18935 10053
rect 18877 10013 18889 10047
rect 18923 10044 18935 10047
rect 20806 10044 20812 10056
rect 18923 10016 20812 10044
rect 18923 10013 18935 10016
rect 18877 10007 18935 10013
rect 16209 9979 16267 9985
rect 16209 9976 16221 9979
rect 13188 9948 15056 9976
rect 15212 9948 16221 9976
rect 11330 9908 11336 9920
rect 11291 9880 11336 9908
rect 11330 9868 11336 9880
rect 11388 9868 11394 9920
rect 12406 9880 12440 9920
rect 12434 9868 12440 9880
rect 12492 9908 12498 9920
rect 15028 9917 15056 9948
rect 16209 9945 16221 9948
rect 16255 9945 16267 9979
rect 16209 9939 16267 9945
rect 16942 9936 16948 9988
rect 17000 9976 17006 9988
rect 17773 9979 17831 9985
rect 17000 9948 17632 9976
rect 17000 9936 17006 9948
rect 13541 9911 13599 9917
rect 13541 9908 13553 9911
rect 12492 9880 13553 9908
rect 12492 9868 12498 9880
rect 13541 9877 13553 9880
rect 13587 9877 13599 9911
rect 13541 9871 13599 9877
rect 15013 9911 15071 9917
rect 15013 9877 15025 9911
rect 15059 9877 15071 9911
rect 15013 9871 15071 9877
rect 15473 9911 15531 9917
rect 15473 9877 15485 9911
rect 15519 9908 15531 9911
rect 15654 9908 15660 9920
rect 15519 9880 15660 9908
rect 15519 9877 15531 9880
rect 15473 9871 15531 9877
rect 15654 9868 15660 9880
rect 15712 9868 15718 9920
rect 17494 9908 17500 9920
rect 17455 9880 17500 9908
rect 17494 9868 17500 9880
rect 17552 9868 17558 9920
rect 17604 9917 17632 9948
rect 17773 9945 17785 9979
rect 17819 9976 17831 9979
rect 18785 9979 18843 9985
rect 18785 9976 18797 9979
rect 17819 9948 18797 9976
rect 17819 9945 17831 9948
rect 17773 9939 17831 9945
rect 18785 9945 18797 9948
rect 18831 9945 18843 9979
rect 18785 9939 18843 9945
rect 17589 9911 17647 9917
rect 17589 9877 17601 9911
rect 17635 9908 17647 9911
rect 18892 9908 18920 10007
rect 20806 10004 20812 10016
rect 20864 10004 20870 10056
rect 21450 10004 21456 10056
rect 21508 10044 21514 10056
rect 21729 10047 21787 10053
rect 21729 10044 21741 10047
rect 21508 10016 21741 10044
rect 21508 10004 21514 10016
rect 21729 10013 21741 10016
rect 21775 10013 21787 10047
rect 22462 10044 22468 10056
rect 22423 10016 22468 10044
rect 21729 10007 21787 10013
rect 22462 10004 22468 10016
rect 22520 10004 22526 10056
rect 22646 10044 22652 10056
rect 22607 10016 22652 10044
rect 22646 10004 22652 10016
rect 22704 10004 22710 10056
rect 24762 10044 24768 10056
rect 24723 10016 24768 10044
rect 24762 10004 24768 10016
rect 24820 10004 24826 10056
rect 32122 10044 32128 10056
rect 32083 10016 32128 10044
rect 32122 10004 32128 10016
rect 32180 10004 32186 10056
rect 32217 10047 32275 10053
rect 32217 10013 32229 10047
rect 32263 10013 32275 10047
rect 32217 10007 32275 10013
rect 32309 10047 32367 10053
rect 32309 10013 32321 10047
rect 32355 10044 32367 10047
rect 32493 10047 32551 10053
rect 32355 10016 32444 10044
rect 32355 10013 32367 10016
rect 32309 10007 32367 10013
rect 22094 9936 22100 9988
rect 22152 9976 22158 9988
rect 26145 9979 26203 9985
rect 26145 9976 26157 9979
rect 22152 9948 26157 9976
rect 22152 9936 22158 9948
rect 26145 9945 26157 9948
rect 26191 9976 26203 9979
rect 26234 9976 26240 9988
rect 26191 9948 26240 9976
rect 26191 9945 26203 9948
rect 26145 9939 26203 9945
rect 26234 9936 26240 9948
rect 26292 9936 26298 9988
rect 31938 9936 31944 9988
rect 31996 9976 32002 9988
rect 32232 9976 32260 10007
rect 31996 9948 32260 9976
rect 31996 9936 32002 9948
rect 17635 9880 18920 9908
rect 32416 9908 32444 10016
rect 32493 10013 32505 10047
rect 32539 10013 32551 10047
rect 32493 10007 32551 10013
rect 33220 10047 33278 10053
rect 33220 10013 33232 10047
rect 33266 10044 33278 10047
rect 33502 10044 33508 10056
rect 33266 10016 33508 10044
rect 33266 10013 33278 10016
rect 33220 10007 33278 10013
rect 32508 9976 32536 10007
rect 33502 10004 33508 10016
rect 33560 10004 33566 10056
rect 34514 10004 34520 10056
rect 34572 10044 34578 10056
rect 34977 10047 35035 10053
rect 34977 10044 34989 10047
rect 34572 10016 34989 10044
rect 34572 10004 34578 10016
rect 34977 10013 34989 10016
rect 35023 10013 35035 10047
rect 35894 10044 35900 10056
rect 35807 10016 35900 10044
rect 34977 10007 35035 10013
rect 35894 10004 35900 10016
rect 35952 10004 35958 10056
rect 36464 10053 36492 10084
rect 37366 10072 37372 10084
rect 37424 10072 37430 10124
rect 38102 10112 38108 10124
rect 38063 10084 38108 10112
rect 38102 10072 38108 10084
rect 38160 10072 38166 10124
rect 36449 10047 36507 10053
rect 36449 10013 36461 10047
rect 36495 10013 36507 10047
rect 37826 10044 37832 10056
rect 37787 10016 37832 10044
rect 36449 10007 36507 10013
rect 37826 10004 37832 10016
rect 37884 10004 37890 10056
rect 33410 9976 33416 9988
rect 32508 9948 33416 9976
rect 33410 9936 33416 9948
rect 33468 9936 33474 9988
rect 33594 9936 33600 9988
rect 33652 9976 33658 9988
rect 35912 9976 35940 10004
rect 33652 9948 35940 9976
rect 33652 9936 33658 9948
rect 32766 9908 32772 9920
rect 32416 9880 32772 9908
rect 17635 9877 17647 9880
rect 17589 9871 17647 9877
rect 32766 9868 32772 9880
rect 32824 9868 32830 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 12434 9704 12440 9716
rect 12406 9664 12440 9704
rect 12492 9664 12498 9716
rect 15378 9664 15384 9716
rect 15436 9704 15442 9716
rect 15473 9707 15531 9713
rect 15473 9704 15485 9707
rect 15436 9676 15485 9704
rect 15436 9664 15442 9676
rect 15473 9673 15485 9676
rect 15519 9673 15531 9707
rect 15473 9667 15531 9673
rect 24121 9707 24179 9713
rect 24121 9673 24133 9707
rect 24167 9673 24179 9707
rect 24121 9667 24179 9673
rect 11057 9639 11115 9645
rect 11057 9605 11069 9639
rect 11103 9636 11115 9639
rect 12406 9636 12434 9664
rect 11103 9608 12434 9636
rect 14645 9639 14703 9645
rect 11103 9605 11115 9608
rect 11057 9599 11115 9605
rect 14645 9605 14657 9639
rect 14691 9636 14703 9639
rect 14734 9636 14740 9648
rect 14691 9608 14740 9636
rect 14691 9605 14703 9608
rect 14645 9599 14703 9605
rect 14734 9596 14740 9608
rect 14792 9596 14798 9648
rect 14918 9596 14924 9648
rect 14976 9636 14982 9648
rect 23474 9636 23480 9648
rect 14976 9608 18368 9636
rect 14976 9596 14982 9608
rect 10873 9571 10931 9577
rect 10873 9537 10885 9571
rect 10919 9537 10931 9571
rect 10873 9531 10931 9537
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9568 11207 9571
rect 11422 9568 11428 9580
rect 11195 9540 11428 9568
rect 11195 9537 11207 9540
rect 11149 9531 11207 9537
rect 10888 9500 10916 9531
rect 11422 9528 11428 9540
rect 11480 9568 11486 9580
rect 11790 9568 11796 9580
rect 11480 9540 11796 9568
rect 11480 9528 11486 9540
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 11977 9571 12035 9577
rect 11977 9537 11989 9571
rect 12023 9537 12035 9571
rect 11977 9531 12035 9537
rect 12069 9571 12127 9577
rect 12069 9537 12081 9571
rect 12115 9537 12127 9571
rect 12069 9531 12127 9537
rect 11238 9500 11244 9512
rect 10888 9472 11244 9500
rect 11238 9460 11244 9472
rect 11296 9460 11302 9512
rect 11330 9460 11336 9512
rect 11388 9500 11394 9512
rect 11992 9500 12020 9531
rect 11388 9472 12020 9500
rect 11388 9460 11394 9472
rect 10689 9435 10747 9441
rect 10689 9401 10701 9435
rect 10735 9432 10747 9435
rect 11054 9432 11060 9444
rect 10735 9404 11060 9432
rect 10735 9401 10747 9404
rect 10689 9395 10747 9401
rect 11054 9392 11060 9404
rect 11112 9392 11118 9444
rect 11698 9432 11704 9444
rect 11659 9404 11704 9432
rect 11698 9392 11704 9404
rect 11756 9392 11762 9444
rect 12084 9432 12112 9531
rect 12158 9528 12164 9580
rect 12216 9568 12222 9580
rect 13265 9571 13323 9577
rect 13265 9568 13277 9571
rect 12216 9540 12261 9568
rect 12452 9540 13277 9568
rect 12216 9528 12222 9540
rect 12452 9512 12480 9540
rect 13265 9537 13277 9540
rect 13311 9537 13323 9571
rect 13265 9531 13323 9537
rect 15565 9571 15623 9577
rect 15565 9537 15577 9571
rect 15611 9568 15623 9571
rect 15654 9568 15660 9580
rect 15611 9540 15660 9568
rect 15611 9537 15623 9540
rect 15565 9531 15623 9537
rect 15654 9528 15660 9540
rect 15712 9568 15718 9580
rect 18340 9577 18368 9608
rect 18524 9608 19334 9636
rect 18325 9571 18383 9577
rect 15712 9540 18184 9568
rect 15712 9528 15718 9540
rect 12434 9460 12440 9512
rect 12492 9500 12498 9512
rect 12986 9500 12992 9512
rect 12492 9472 12537 9500
rect 12947 9472 12992 9500
rect 12492 9460 12498 9472
rect 12986 9460 12992 9472
rect 13044 9460 13050 9512
rect 15749 9503 15807 9509
rect 15749 9469 15761 9503
rect 15795 9500 15807 9503
rect 18046 9500 18052 9512
rect 15795 9472 18052 9500
rect 15795 9469 15807 9472
rect 15749 9463 15807 9469
rect 18046 9460 18052 9472
rect 18104 9460 18110 9512
rect 18156 9500 18184 9540
rect 18325 9537 18337 9571
rect 18371 9568 18383 9571
rect 18414 9568 18420 9580
rect 18371 9540 18420 9568
rect 18371 9537 18383 9540
rect 18325 9531 18383 9537
rect 18414 9528 18420 9540
rect 18472 9528 18478 9580
rect 18524 9500 18552 9608
rect 19150 9568 19156 9580
rect 19111 9540 19156 9568
rect 19150 9528 19156 9540
rect 19208 9528 19214 9580
rect 18156 9472 18552 9500
rect 19306 9500 19334 9608
rect 19536 9608 22692 9636
rect 19536 9577 19564 9608
rect 19521 9571 19579 9577
rect 19521 9537 19533 9571
rect 19567 9537 19579 9571
rect 21082 9568 21088 9580
rect 21043 9540 21088 9568
rect 19521 9531 19579 9537
rect 21082 9528 21088 9540
rect 21140 9528 21146 9580
rect 21177 9571 21235 9577
rect 21177 9537 21189 9571
rect 21223 9568 21235 9571
rect 21266 9568 21272 9580
rect 21223 9540 21272 9568
rect 21223 9537 21235 9540
rect 21177 9531 21235 9537
rect 21266 9528 21272 9540
rect 21324 9568 21330 9580
rect 22278 9568 22284 9580
rect 21324 9540 22284 9568
rect 21324 9528 21330 9540
rect 22278 9528 22284 9540
rect 22336 9528 22342 9580
rect 19886 9500 19892 9512
rect 19306 9472 19892 9500
rect 19886 9460 19892 9472
rect 19944 9460 19950 9512
rect 21361 9503 21419 9509
rect 21361 9469 21373 9503
rect 21407 9500 21419 9503
rect 22462 9500 22468 9512
rect 21407 9472 22468 9500
rect 21407 9469 21419 9472
rect 21361 9463 21419 9469
rect 22462 9460 22468 9472
rect 22520 9460 22526 9512
rect 22554 9432 22560 9444
rect 12084 9404 13032 9432
rect 11974 9324 11980 9376
rect 12032 9364 12038 9376
rect 12345 9367 12403 9373
rect 12345 9364 12357 9367
rect 12032 9336 12357 9364
rect 12032 9324 12038 9336
rect 12345 9333 12357 9336
rect 12391 9333 12403 9367
rect 13004 9364 13032 9404
rect 13924 9404 15332 9432
rect 13924 9364 13952 9404
rect 13004 9336 13952 9364
rect 12345 9327 12403 9333
rect 14642 9324 14648 9376
rect 14700 9364 14706 9376
rect 15105 9367 15163 9373
rect 15105 9364 15117 9367
rect 14700 9336 15117 9364
rect 14700 9324 14706 9336
rect 15105 9333 15117 9336
rect 15151 9333 15163 9367
rect 15304 9364 15332 9404
rect 19306 9404 22560 9432
rect 15562 9364 15568 9376
rect 15304 9336 15568 9364
rect 15105 9327 15163 9333
rect 15562 9324 15568 9336
rect 15620 9364 15626 9376
rect 18322 9364 18328 9376
rect 15620 9336 18328 9364
rect 15620 9324 15626 9336
rect 18322 9324 18328 9336
rect 18380 9324 18386 9376
rect 18414 9324 18420 9376
rect 18472 9364 18478 9376
rect 19306 9364 19334 9404
rect 22554 9392 22560 9404
rect 22612 9392 22618 9444
rect 18472 9336 19334 9364
rect 18472 9324 18478 9336
rect 20530 9324 20536 9376
rect 20588 9364 20594 9376
rect 20717 9367 20775 9373
rect 20717 9364 20729 9367
rect 20588 9336 20729 9364
rect 20588 9324 20594 9336
rect 20717 9333 20729 9336
rect 20763 9333 20775 9367
rect 22664 9364 22692 9608
rect 22756 9608 23480 9636
rect 22756 9577 22784 9608
rect 23474 9596 23480 9608
rect 23532 9596 23538 9648
rect 24136 9636 24164 9667
rect 24854 9664 24860 9716
rect 24912 9704 24918 9716
rect 24912 9676 26188 9704
rect 24912 9664 24918 9676
rect 24762 9636 24768 9648
rect 24136 9608 24768 9636
rect 24762 9596 24768 9608
rect 24820 9636 24826 9648
rect 24949 9639 25007 9645
rect 24949 9636 24961 9639
rect 24820 9608 24961 9636
rect 24820 9596 24826 9608
rect 24949 9605 24961 9608
rect 24995 9605 25007 9639
rect 24949 9599 25007 9605
rect 25041 9639 25099 9645
rect 25041 9605 25053 9639
rect 25087 9636 25099 9639
rect 25222 9636 25228 9648
rect 25087 9608 25228 9636
rect 25087 9605 25099 9608
rect 25041 9599 25099 9605
rect 25222 9596 25228 9608
rect 25280 9596 25286 9648
rect 26160 9636 26188 9676
rect 26234 9664 26240 9716
rect 26292 9704 26298 9716
rect 33226 9704 33232 9716
rect 26292 9676 33232 9704
rect 26292 9664 26298 9676
rect 33226 9664 33232 9676
rect 33284 9664 33290 9716
rect 33594 9704 33600 9716
rect 33555 9676 33600 9704
rect 33594 9664 33600 9676
rect 33652 9664 33658 9716
rect 26329 9639 26387 9645
rect 26329 9636 26341 9639
rect 26160 9608 26341 9636
rect 26329 9605 26341 9608
rect 26375 9636 26387 9639
rect 26418 9636 26424 9648
rect 26375 9608 26424 9636
rect 26375 9605 26387 9608
rect 26329 9599 26387 9605
rect 26418 9596 26424 9608
rect 26476 9596 26482 9648
rect 29178 9636 29184 9648
rect 29139 9608 29184 9636
rect 29178 9596 29184 9608
rect 29236 9596 29242 9648
rect 30190 9596 30196 9648
rect 30248 9636 30254 9648
rect 30834 9636 30840 9648
rect 30248 9608 30420 9636
rect 30795 9608 30840 9636
rect 30248 9596 30254 9608
rect 22741 9571 22799 9577
rect 22741 9537 22753 9571
rect 22787 9537 22799 9571
rect 22741 9531 22799 9537
rect 23008 9571 23066 9577
rect 23008 9537 23020 9571
rect 23054 9568 23066 9571
rect 25869 9571 25927 9577
rect 25869 9568 25881 9571
rect 23054 9540 24624 9568
rect 23054 9537 23066 9540
rect 23008 9531 23066 9537
rect 24596 9441 24624 9540
rect 25792 9540 25881 9568
rect 25225 9503 25283 9509
rect 25225 9469 25237 9503
rect 25271 9500 25283 9503
rect 25314 9500 25320 9512
rect 25271 9472 25320 9500
rect 25271 9469 25283 9472
rect 25225 9463 25283 9469
rect 25314 9460 25320 9472
rect 25372 9460 25378 9512
rect 24581 9435 24639 9441
rect 24581 9401 24593 9435
rect 24627 9401 24639 9435
rect 24581 9395 24639 9401
rect 25792 9364 25820 9540
rect 25869 9537 25881 9540
rect 25915 9537 25927 9571
rect 25869 9531 25927 9537
rect 26694 9528 26700 9580
rect 26752 9568 26758 9580
rect 27341 9571 27399 9577
rect 27341 9568 27353 9571
rect 26752 9540 27353 9568
rect 26752 9528 26758 9540
rect 27341 9537 27353 9540
rect 27387 9537 27399 9571
rect 27341 9531 27399 9537
rect 27608 9571 27666 9577
rect 27608 9537 27620 9571
rect 27654 9568 27666 9571
rect 27982 9568 27988 9580
rect 27654 9540 27988 9568
rect 27654 9537 27666 9540
rect 27608 9531 27666 9537
rect 27982 9528 27988 9540
rect 28040 9528 28046 9580
rect 29457 9571 29515 9577
rect 29457 9537 29469 9571
rect 29503 9537 29515 9571
rect 29457 9531 29515 9537
rect 29549 9571 29607 9577
rect 29549 9537 29561 9571
rect 29595 9537 29607 9571
rect 29549 9531 29607 9537
rect 28350 9392 28356 9444
rect 28408 9432 28414 9444
rect 28721 9435 28779 9441
rect 28721 9432 28733 9435
rect 28408 9404 28733 9432
rect 28408 9392 28414 9404
rect 28721 9401 28733 9404
rect 28767 9432 28779 9435
rect 29472 9432 29500 9531
rect 28767 9404 29500 9432
rect 29564 9432 29592 9531
rect 29638 9528 29644 9580
rect 29696 9568 29702 9580
rect 29822 9568 29828 9580
rect 29696 9540 29741 9568
rect 29783 9540 29828 9568
rect 29696 9528 29702 9540
rect 29822 9528 29828 9540
rect 29880 9528 29886 9580
rect 30282 9568 30288 9580
rect 30243 9540 30288 9568
rect 30282 9528 30288 9540
rect 30340 9528 30346 9580
rect 30392 9577 30420 9608
rect 30834 9596 30840 9608
rect 30892 9596 30898 9648
rect 32122 9596 32128 9648
rect 32180 9636 32186 9648
rect 32582 9636 32588 9648
rect 32180 9608 32588 9636
rect 32180 9596 32186 9608
rect 32582 9596 32588 9608
rect 32640 9636 32646 9648
rect 32677 9639 32735 9645
rect 32677 9636 32689 9639
rect 32640 9608 32689 9636
rect 32640 9596 32646 9608
rect 32677 9605 32689 9608
rect 32723 9605 32735 9639
rect 32677 9599 32735 9605
rect 32766 9596 32772 9648
rect 32824 9636 32830 9648
rect 38102 9636 38108 9648
rect 32824 9608 34744 9636
rect 38063 9608 38108 9636
rect 32824 9596 32830 9608
rect 30377 9571 30435 9577
rect 30377 9537 30389 9571
rect 30423 9537 30435 9571
rect 30377 9531 30435 9537
rect 32030 9528 32036 9580
rect 32088 9568 32094 9580
rect 34146 9568 34152 9580
rect 32088 9540 32812 9568
rect 34107 9540 34152 9568
rect 32088 9528 32094 9540
rect 32784 9512 32812 9540
rect 34146 9528 34152 9540
rect 34204 9528 34210 9580
rect 34716 9577 34744 9608
rect 38102 9596 38108 9608
rect 38160 9596 38166 9648
rect 34701 9571 34759 9577
rect 34701 9537 34713 9571
rect 34747 9568 34759 9571
rect 35526 9568 35532 9580
rect 34747 9540 35532 9568
rect 34747 9537 34759 9540
rect 34701 9531 34759 9537
rect 35526 9528 35532 9540
rect 35584 9528 35590 9580
rect 37826 9568 37832 9580
rect 37787 9540 37832 9568
rect 37826 9528 37832 9540
rect 37884 9528 37890 9580
rect 30742 9460 30748 9512
rect 30800 9500 30806 9512
rect 32766 9500 32772 9512
rect 30800 9472 32536 9500
rect 32727 9472 32772 9500
rect 30800 9460 30806 9472
rect 29914 9432 29920 9444
rect 29564 9404 29920 9432
rect 28767 9401 28779 9404
rect 28721 9395 28779 9401
rect 29564 9364 29592 9404
rect 29914 9392 29920 9404
rect 29972 9432 29978 9444
rect 32508 9432 32536 9472
rect 32766 9460 32772 9472
rect 32824 9460 32830 9512
rect 32861 9503 32919 9509
rect 32861 9469 32873 9503
rect 32907 9469 32919 9503
rect 32861 9463 32919 9469
rect 32876 9432 32904 9463
rect 29972 9404 32444 9432
rect 32508 9404 32904 9432
rect 29972 9392 29978 9404
rect 22664 9336 29592 9364
rect 20717 9327 20775 9333
rect 31754 9324 31760 9376
rect 31812 9364 31818 9376
rect 32309 9367 32367 9373
rect 32309 9364 32321 9367
rect 31812 9336 32321 9364
rect 31812 9324 31818 9336
rect 32309 9333 32321 9336
rect 32355 9333 32367 9367
rect 32416 9364 32444 9404
rect 34146 9364 34152 9376
rect 32416 9336 34152 9364
rect 32309 9327 32367 9333
rect 34146 9324 34152 9336
rect 34204 9324 34210 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 10870 9160 10876 9172
rect 10831 9132 10876 9160
rect 10870 9120 10876 9132
rect 10928 9120 10934 9172
rect 17126 9120 17132 9172
rect 17184 9160 17190 9172
rect 26237 9163 26295 9169
rect 17184 9132 20944 9160
rect 17184 9120 17190 9132
rect 16758 9052 16764 9104
rect 16816 9092 16822 9104
rect 16816 9064 17540 9092
rect 16816 9052 16822 9064
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 9024 10563 9027
rect 11054 9024 11060 9036
rect 10551 8996 11060 9024
rect 10551 8993 10563 8996
rect 10505 8987 10563 8993
rect 11054 8984 11060 8996
rect 11112 9024 11118 9036
rect 12158 9024 12164 9036
rect 11112 8996 12164 9024
rect 11112 8984 11118 8996
rect 12158 8984 12164 8996
rect 12216 8984 12222 9036
rect 12526 8984 12532 9036
rect 12584 9024 12590 9036
rect 12621 9027 12679 9033
rect 12621 9024 12633 9027
rect 12584 8996 12633 9024
rect 12584 8984 12590 8996
rect 12621 8993 12633 8996
rect 12667 8993 12679 9027
rect 12621 8987 12679 8993
rect 12894 8984 12900 9036
rect 12952 9024 12958 9036
rect 12989 9027 13047 9033
rect 12989 9024 13001 9027
rect 12952 8996 13001 9024
rect 12952 8984 12958 8996
rect 12989 8993 13001 8996
rect 13035 8993 13047 9027
rect 12989 8987 13047 8993
rect 13081 9027 13139 9033
rect 13081 8993 13093 9027
rect 13127 9024 13139 9027
rect 13538 9024 13544 9036
rect 13127 8996 13544 9024
rect 13127 8993 13139 8996
rect 13081 8987 13139 8993
rect 13538 8984 13544 8996
rect 13596 8984 13602 9036
rect 16945 9027 17003 9033
rect 16945 8993 16957 9027
rect 16991 9024 17003 9027
rect 17310 9024 17316 9036
rect 16991 8996 17316 9024
rect 16991 8993 17003 8996
rect 16945 8987 17003 8993
rect 17310 8984 17316 8996
rect 17368 8984 17374 9036
rect 10689 8959 10747 8965
rect 10689 8925 10701 8959
rect 10735 8956 10747 8959
rect 11330 8956 11336 8968
rect 10735 8928 11336 8956
rect 10735 8925 10747 8928
rect 10689 8919 10747 8925
rect 11330 8916 11336 8928
rect 11388 8916 11394 8968
rect 14458 8956 14464 8968
rect 14419 8928 14464 8956
rect 14458 8916 14464 8928
rect 14516 8916 14522 8968
rect 14642 8956 14648 8968
rect 14603 8928 14648 8956
rect 14642 8916 14648 8928
rect 14700 8916 14706 8968
rect 15654 8956 15660 8968
rect 15615 8928 15660 8956
rect 15654 8916 15660 8928
rect 15712 8916 15718 8968
rect 15749 8959 15807 8965
rect 15749 8925 15761 8959
rect 15795 8956 15807 8959
rect 16758 8956 16764 8968
rect 15795 8928 16764 8956
rect 15795 8925 15807 8928
rect 15749 8919 15807 8925
rect 16758 8916 16764 8928
rect 16816 8916 16822 8968
rect 17512 8965 17540 9064
rect 18414 9052 18420 9104
rect 18472 9092 18478 9104
rect 18509 9095 18567 9101
rect 18509 9092 18521 9095
rect 18472 9064 18521 9092
rect 18472 9052 18478 9064
rect 18509 9061 18521 9064
rect 18555 9061 18567 9095
rect 18509 9055 18567 9061
rect 19429 9095 19487 9101
rect 19429 9061 19441 9095
rect 19475 9061 19487 9095
rect 20806 9092 20812 9104
rect 20767 9064 20812 9092
rect 19429 9055 19487 9061
rect 18693 9027 18751 9033
rect 18693 8993 18705 9027
rect 18739 9024 18751 9027
rect 18782 9024 18788 9036
rect 18739 8996 18788 9024
rect 18739 8993 18751 8996
rect 18693 8987 18751 8993
rect 18782 8984 18788 8996
rect 18840 8984 18846 9036
rect 17497 8959 17555 8965
rect 17497 8925 17509 8959
rect 17543 8956 17555 8959
rect 17862 8956 17868 8968
rect 17543 8928 17868 8956
rect 17543 8925 17555 8928
rect 17497 8919 17555 8925
rect 17862 8916 17868 8928
rect 17920 8916 17926 8968
rect 18506 8956 18512 8968
rect 18419 8928 18512 8956
rect 18506 8916 18512 8928
rect 18564 8956 18570 8968
rect 19444 8956 19472 9055
rect 20806 9052 20812 9064
rect 20864 9052 20870 9104
rect 20916 9092 20944 9132
rect 26237 9129 26249 9163
rect 26283 9160 26295 9163
rect 26326 9160 26332 9172
rect 26283 9132 26332 9160
rect 26283 9129 26295 9132
rect 26237 9123 26295 9129
rect 26326 9120 26332 9132
rect 26384 9120 26390 9172
rect 27982 9160 27988 9172
rect 27943 9132 27988 9160
rect 27982 9120 27988 9132
rect 28040 9120 28046 9172
rect 29546 9120 29552 9172
rect 29604 9160 29610 9172
rect 31478 9160 31484 9172
rect 29604 9132 31484 9160
rect 29604 9120 29610 9132
rect 31478 9120 31484 9132
rect 31536 9120 31542 9172
rect 32582 9160 32588 9172
rect 32543 9132 32588 9160
rect 32582 9120 32588 9132
rect 32640 9120 32646 9172
rect 33410 9160 33416 9172
rect 33371 9132 33416 9160
rect 33410 9120 33416 9132
rect 33468 9120 33474 9172
rect 29638 9092 29644 9104
rect 20916 9064 29644 9092
rect 29638 9052 29644 9064
rect 29696 9052 29702 9104
rect 35342 9052 35348 9104
rect 35400 9092 35406 9104
rect 35437 9095 35495 9101
rect 35437 9092 35449 9095
rect 35400 9064 35449 9092
rect 35400 9052 35406 9064
rect 35437 9061 35449 9064
rect 35483 9061 35495 9095
rect 35437 9055 35495 9061
rect 36170 9052 36176 9104
rect 36228 9092 36234 9104
rect 36228 9064 36584 9092
rect 36228 9052 36234 9064
rect 20073 9027 20131 9033
rect 20073 8993 20085 9027
rect 20119 9024 20131 9027
rect 20162 9024 20168 9036
rect 20119 8996 20168 9024
rect 20119 8993 20131 8996
rect 20073 8987 20131 8993
rect 20162 8984 20168 8996
rect 20220 8984 20226 9036
rect 21361 9027 21419 9033
rect 21361 8993 21373 9027
rect 21407 9024 21419 9027
rect 21910 9024 21916 9036
rect 21407 8996 21916 9024
rect 21407 8993 21419 8996
rect 21361 8987 21419 8993
rect 21910 8984 21916 8996
rect 21968 8984 21974 9036
rect 25222 8984 25228 9036
rect 25280 9024 25286 9036
rect 25501 9027 25559 9033
rect 25501 9024 25513 9027
rect 25280 8996 25513 9024
rect 25280 8984 25286 8996
rect 25501 8993 25513 8996
rect 25547 8993 25559 9027
rect 25682 9024 25688 9036
rect 25643 8996 25688 9024
rect 25501 8987 25559 8993
rect 25682 8984 25688 8996
rect 25740 8984 25746 9036
rect 26050 8984 26056 9036
rect 26108 9024 26114 9036
rect 26108 8996 26740 9024
rect 26108 8984 26114 8996
rect 24210 8956 24216 8968
rect 18564 8928 19472 8956
rect 19720 8928 24216 8956
rect 18564 8916 18570 8928
rect 14829 8891 14887 8897
rect 14829 8857 14841 8891
rect 14875 8888 14887 8891
rect 14918 8888 14924 8900
rect 14875 8860 14924 8888
rect 14875 8857 14887 8860
rect 14829 8851 14887 8857
rect 14918 8848 14924 8860
rect 14976 8848 14982 8900
rect 16669 8891 16727 8897
rect 16669 8857 16681 8891
rect 16715 8888 16727 8891
rect 17589 8891 17647 8897
rect 17589 8888 17601 8891
rect 16715 8860 17601 8888
rect 16715 8857 16727 8860
rect 16669 8851 16727 8857
rect 17589 8857 17601 8860
rect 17635 8857 17647 8891
rect 18874 8888 18880 8900
rect 18835 8860 18880 8888
rect 17589 8851 17647 8857
rect 18874 8848 18880 8860
rect 18932 8848 18938 8900
rect 19242 8848 19248 8900
rect 19300 8888 19306 8900
rect 19720 8888 19748 8928
rect 24210 8916 24216 8928
rect 24268 8916 24274 8968
rect 25409 8959 25467 8965
rect 25409 8925 25421 8959
rect 25455 8956 25467 8959
rect 25866 8956 25872 8968
rect 25455 8928 25872 8956
rect 25455 8925 25467 8928
rect 25409 8919 25467 8925
rect 25866 8916 25872 8928
rect 25924 8956 25930 8968
rect 26712 8965 26740 8996
rect 27522 8984 27528 9036
rect 27580 9024 27586 9036
rect 28445 9027 28503 9033
rect 28445 9024 28457 9027
rect 27580 8996 28457 9024
rect 27580 8984 27586 8996
rect 28445 8993 28457 8996
rect 28491 8993 28503 9027
rect 28445 8987 28503 8993
rect 28537 9027 28595 9033
rect 28537 8993 28549 9027
rect 28583 8993 28595 9027
rect 36078 9024 36084 9036
rect 36039 8996 36084 9024
rect 28537 8987 28595 8993
rect 26421 8959 26479 8965
rect 26421 8956 26433 8959
rect 25924 8928 26433 8956
rect 25924 8916 25930 8928
rect 26421 8925 26433 8928
rect 26467 8925 26479 8959
rect 26421 8919 26479 8925
rect 26697 8959 26755 8965
rect 26697 8925 26709 8959
rect 26743 8925 26755 8959
rect 28350 8956 28356 8968
rect 28311 8928 28356 8956
rect 26697 8919 26755 8925
rect 28350 8916 28356 8928
rect 28408 8916 28414 8968
rect 28552 8956 28580 8987
rect 36078 8984 36084 8996
rect 36136 8984 36142 9036
rect 36556 9033 36584 9064
rect 36541 9027 36599 9033
rect 36541 8993 36553 9027
rect 36587 8993 36599 9027
rect 36541 8987 36599 8993
rect 28460 8928 28580 8956
rect 30009 8959 30067 8965
rect 21082 8888 21088 8900
rect 19300 8860 19748 8888
rect 19812 8860 21088 8888
rect 19300 8848 19306 8860
rect 12710 8780 12716 8832
rect 12768 8820 12774 8832
rect 13265 8823 13323 8829
rect 13265 8820 13277 8823
rect 12768 8792 13277 8820
rect 12768 8780 12774 8792
rect 13265 8789 13277 8792
rect 13311 8789 13323 8823
rect 16298 8820 16304 8832
rect 16259 8792 16304 8820
rect 13265 8783 13323 8789
rect 16298 8780 16304 8792
rect 16356 8780 16362 8832
rect 17862 8780 17868 8832
rect 17920 8820 17926 8832
rect 19812 8829 19840 8860
rect 21082 8848 21088 8860
rect 21140 8848 21146 8900
rect 21266 8888 21272 8900
rect 21227 8860 21272 8888
rect 21266 8848 21272 8860
rect 21324 8848 21330 8900
rect 24228 8888 24256 8916
rect 26142 8888 26148 8900
rect 24228 8860 26148 8888
rect 26142 8848 26148 8860
rect 26200 8888 26206 8900
rect 26605 8891 26663 8897
rect 26605 8888 26617 8891
rect 26200 8860 26617 8888
rect 26200 8848 26206 8860
rect 26605 8857 26617 8860
rect 26651 8857 26663 8891
rect 26605 8851 26663 8857
rect 19797 8823 19855 8829
rect 19797 8820 19809 8823
rect 17920 8792 19809 8820
rect 17920 8780 17926 8792
rect 19797 8789 19809 8792
rect 19843 8789 19855 8823
rect 19797 8783 19855 8789
rect 19886 8780 19892 8832
rect 19944 8820 19950 8832
rect 21284 8820 21312 8848
rect 28460 8832 28488 8928
rect 30009 8925 30021 8959
rect 30055 8925 30067 8959
rect 30009 8919 30067 8925
rect 30101 8959 30159 8965
rect 30101 8925 30113 8959
rect 30147 8956 30159 8959
rect 30190 8956 30196 8968
rect 30147 8928 30196 8956
rect 30147 8925 30159 8928
rect 30101 8919 30159 8925
rect 25038 8820 25044 8832
rect 19944 8792 21312 8820
rect 24999 8792 25044 8820
rect 19944 8780 19950 8792
rect 25038 8780 25044 8792
rect 25096 8780 25102 8832
rect 25314 8780 25320 8832
rect 25372 8820 25378 8832
rect 28442 8820 28448 8832
rect 25372 8792 28448 8820
rect 25372 8780 25378 8792
rect 28442 8780 28448 8792
rect 28500 8780 28506 8832
rect 30024 8820 30052 8919
rect 30190 8916 30196 8928
rect 30248 8916 30254 8968
rect 31202 8956 31208 8968
rect 31163 8928 31208 8956
rect 31202 8916 31208 8928
rect 31260 8916 31266 8968
rect 31472 8959 31530 8965
rect 31472 8925 31484 8959
rect 31518 8956 31530 8959
rect 31754 8956 31760 8968
rect 31518 8928 31760 8956
rect 31518 8925 31530 8928
rect 31472 8919 31530 8925
rect 31754 8916 31760 8928
rect 31812 8916 31818 8968
rect 32858 8916 32864 8968
rect 32916 8956 32922 8968
rect 33229 8959 33287 8965
rect 33229 8956 33241 8959
rect 32916 8928 33241 8956
rect 32916 8916 32922 8928
rect 33229 8925 33241 8928
rect 33275 8925 33287 8959
rect 35434 8956 35440 8968
rect 35395 8928 35440 8956
rect 33229 8919 33287 8925
rect 35434 8916 35440 8928
rect 35492 8916 35498 8968
rect 35894 8916 35900 8968
rect 35952 8956 35958 8968
rect 36173 8959 36231 8965
rect 36173 8956 36185 8959
rect 35952 8928 36185 8956
rect 35952 8916 35958 8928
rect 36173 8925 36185 8928
rect 36219 8925 36231 8959
rect 36173 8919 36231 8925
rect 36817 8959 36875 8965
rect 36817 8925 36829 8959
rect 36863 8925 36875 8959
rect 36817 8919 36875 8925
rect 37829 8959 37887 8965
rect 37829 8925 37841 8959
rect 37875 8925 37887 8959
rect 37829 8919 37887 8925
rect 30466 8848 30472 8900
rect 30524 8888 30530 8900
rect 30561 8891 30619 8897
rect 30561 8888 30573 8891
rect 30524 8860 30573 8888
rect 30524 8848 30530 8860
rect 30561 8857 30573 8860
rect 30607 8857 30619 8891
rect 30561 8851 30619 8857
rect 30926 8848 30932 8900
rect 30984 8888 30990 8900
rect 33045 8891 33103 8897
rect 33045 8888 33057 8891
rect 30984 8860 33057 8888
rect 30984 8848 30990 8860
rect 33045 8857 33057 8860
rect 33091 8888 33103 8891
rect 33870 8888 33876 8900
rect 33091 8860 33876 8888
rect 33091 8857 33103 8860
rect 33045 8851 33103 8857
rect 33870 8848 33876 8860
rect 33928 8848 33934 8900
rect 36832 8888 36860 8919
rect 37734 8888 37740 8900
rect 36832 8860 37740 8888
rect 37734 8848 37740 8860
rect 37792 8848 37798 8900
rect 31386 8820 31392 8832
rect 30024 8792 31392 8820
rect 31386 8780 31392 8792
rect 31444 8780 31450 8832
rect 31478 8780 31484 8832
rect 31536 8820 31542 8832
rect 37844 8820 37872 8919
rect 38102 8888 38108 8900
rect 38063 8860 38108 8888
rect 38102 8848 38108 8860
rect 38160 8848 38166 8900
rect 31536 8792 37872 8820
rect 31536 8780 31542 8792
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 12069 8619 12127 8625
rect 12069 8585 12081 8619
rect 12115 8616 12127 8619
rect 12434 8616 12440 8628
rect 12115 8588 12440 8616
rect 12115 8585 12127 8588
rect 12069 8579 12127 8585
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 14458 8576 14464 8628
rect 14516 8616 14522 8628
rect 16945 8619 17003 8625
rect 16945 8616 16957 8619
rect 14516 8588 16957 8616
rect 14516 8576 14522 8588
rect 16945 8585 16957 8588
rect 16991 8585 17003 8619
rect 21361 8619 21419 8625
rect 21361 8616 21373 8619
rect 16945 8579 17003 8585
rect 17052 8588 21373 8616
rect 14918 8548 14924 8560
rect 13924 8520 14924 8548
rect 11790 8480 11796 8492
rect 11751 8452 11796 8480
rect 11790 8440 11796 8452
rect 11848 8440 11854 8492
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8480 11943 8483
rect 12802 8480 12808 8492
rect 11931 8452 12808 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 12802 8440 12808 8452
rect 12860 8440 12866 8492
rect 13924 8489 13952 8520
rect 14918 8508 14924 8520
rect 14976 8508 14982 8560
rect 17052 8548 17080 8588
rect 21361 8585 21373 8588
rect 21407 8616 21419 8619
rect 25866 8616 25872 8628
rect 21407 8588 22232 8616
rect 25827 8588 25872 8616
rect 21407 8585 21419 8588
rect 21361 8579 21419 8585
rect 18506 8548 18512 8560
rect 15028 8520 17080 8548
rect 18467 8520 18512 8548
rect 13909 8483 13967 8489
rect 13909 8449 13921 8483
rect 13955 8449 13967 8483
rect 14826 8480 14832 8492
rect 14787 8452 14832 8480
rect 13909 8443 13967 8449
rect 14826 8440 14832 8452
rect 14884 8440 14890 8492
rect 14458 8372 14464 8424
rect 14516 8412 14522 8424
rect 15028 8412 15056 8520
rect 18506 8508 18512 8520
rect 18564 8508 18570 8560
rect 22204 8557 22232 8588
rect 25866 8576 25872 8588
rect 25924 8576 25930 8628
rect 27522 8576 27528 8628
rect 27580 8616 27586 8628
rect 27617 8619 27675 8625
rect 27617 8616 27629 8619
rect 27580 8588 27629 8616
rect 27580 8576 27586 8588
rect 27617 8585 27629 8588
rect 27663 8585 27675 8619
rect 27617 8579 27675 8585
rect 29178 8576 29184 8628
rect 29236 8616 29242 8628
rect 31386 8616 31392 8628
rect 29236 8588 30972 8616
rect 31347 8588 31392 8616
rect 29236 8576 29242 8588
rect 20165 8551 20223 8557
rect 20165 8517 20177 8551
rect 20211 8548 20223 8551
rect 22005 8551 22063 8557
rect 22005 8548 22017 8551
rect 20211 8520 22017 8548
rect 20211 8517 20223 8520
rect 20165 8511 20223 8517
rect 22005 8517 22017 8520
rect 22051 8517 22063 8551
rect 22005 8511 22063 8517
rect 22189 8551 22247 8557
rect 22189 8517 22201 8551
rect 22235 8517 22247 8551
rect 22189 8511 22247 8517
rect 24756 8551 24814 8557
rect 24756 8517 24768 8551
rect 24802 8548 24814 8551
rect 25038 8548 25044 8560
rect 24802 8520 25044 8548
rect 24802 8517 24814 8520
rect 24756 8511 24814 8517
rect 25038 8508 25044 8520
rect 25096 8508 25102 8560
rect 28442 8508 28448 8560
rect 28500 8548 28506 8560
rect 29825 8551 29883 8557
rect 29825 8548 29837 8551
rect 28500 8520 29837 8548
rect 28500 8508 28506 8520
rect 29825 8517 29837 8520
rect 29871 8548 29883 8551
rect 30742 8548 30748 8560
rect 29871 8520 30748 8548
rect 29871 8517 29883 8520
rect 29825 8511 29883 8517
rect 30742 8508 30748 8520
rect 30800 8508 30806 8560
rect 30944 8548 30972 8588
rect 31386 8576 31392 8588
rect 31444 8576 31450 8628
rect 32766 8576 32772 8628
rect 32824 8616 32830 8628
rect 32953 8619 33011 8625
rect 32953 8616 32965 8619
rect 32824 8588 32965 8616
rect 32824 8576 32830 8588
rect 32953 8585 32965 8588
rect 32999 8585 33011 8619
rect 32953 8579 33011 8585
rect 36078 8576 36084 8628
rect 36136 8616 36142 8628
rect 36173 8619 36231 8625
rect 36173 8616 36185 8619
rect 36136 8588 36185 8616
rect 36136 8576 36142 8588
rect 36173 8585 36185 8588
rect 36219 8585 36231 8619
rect 36173 8579 36231 8585
rect 37734 8576 37740 8628
rect 37792 8616 37798 8628
rect 37829 8619 37887 8625
rect 37829 8616 37841 8619
rect 37792 8588 37841 8616
rect 37792 8576 37798 8588
rect 37829 8585 37841 8588
rect 37875 8585 37887 8619
rect 37829 8579 37887 8585
rect 33781 8551 33839 8557
rect 30944 8520 31064 8548
rect 16117 8483 16175 8489
rect 16117 8449 16129 8483
rect 16163 8449 16175 8483
rect 16117 8443 16175 8449
rect 14516 8384 15056 8412
rect 14516 8372 14522 8384
rect 15562 8304 15568 8356
rect 15620 8344 15626 8356
rect 16132 8344 16160 8443
rect 16758 8440 16764 8492
rect 16816 8480 16822 8492
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 16816 8452 16865 8480
rect 16816 8440 16822 8452
rect 16853 8449 16865 8452
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 17037 8483 17095 8489
rect 17037 8449 17049 8483
rect 17083 8449 17095 8483
rect 17037 8443 17095 8449
rect 18693 8483 18751 8489
rect 18693 8449 18705 8483
rect 18739 8480 18751 8483
rect 18874 8480 18880 8492
rect 18739 8452 18880 8480
rect 18739 8449 18751 8452
rect 18693 8443 18751 8449
rect 16209 8415 16267 8421
rect 16209 8381 16221 8415
rect 16255 8412 16267 8415
rect 16482 8412 16488 8424
rect 16255 8384 16488 8412
rect 16255 8381 16267 8384
rect 16209 8375 16267 8381
rect 16482 8372 16488 8384
rect 16540 8412 16546 8424
rect 17052 8412 17080 8443
rect 18874 8440 18880 8452
rect 18932 8440 18938 8492
rect 20349 8483 20407 8489
rect 20349 8449 20361 8483
rect 20395 8480 20407 8483
rect 20714 8480 20720 8492
rect 20395 8452 20720 8480
rect 20395 8449 20407 8452
rect 20349 8443 20407 8449
rect 20714 8440 20720 8452
rect 20772 8480 20778 8492
rect 21085 8483 21143 8489
rect 21085 8480 21097 8483
rect 20772 8452 21097 8480
rect 20772 8440 20778 8452
rect 21085 8449 21097 8452
rect 21131 8449 21143 8483
rect 21269 8483 21327 8489
rect 21269 8480 21281 8483
rect 21085 8443 21143 8449
rect 21192 8452 21281 8480
rect 16540 8384 17080 8412
rect 16540 8372 16546 8384
rect 18782 8372 18788 8424
rect 18840 8372 18846 8424
rect 20530 8412 20536 8424
rect 20491 8384 20536 8412
rect 20530 8372 20536 8384
rect 20588 8372 20594 8424
rect 20625 8415 20683 8421
rect 20625 8381 20637 8415
rect 20671 8412 20683 8415
rect 20898 8412 20904 8424
rect 20671 8384 20904 8412
rect 20671 8381 20683 8384
rect 20625 8375 20683 8381
rect 20898 8372 20904 8384
rect 20956 8372 20962 8424
rect 18800 8344 18828 8372
rect 15620 8316 18828 8344
rect 15620 8304 15626 8316
rect 19978 8304 19984 8356
rect 20036 8344 20042 8356
rect 20548 8344 20576 8372
rect 21192 8344 21220 8452
rect 21269 8449 21281 8452
rect 21315 8449 21327 8483
rect 21269 8443 21327 8449
rect 23474 8440 23480 8492
rect 23532 8480 23538 8492
rect 24489 8483 24547 8489
rect 24489 8480 24501 8483
rect 23532 8452 24501 8480
rect 23532 8440 23538 8452
rect 24489 8449 24501 8452
rect 24535 8449 24547 8483
rect 24489 8443 24547 8449
rect 27525 8483 27583 8489
rect 27525 8449 27537 8483
rect 27571 8480 27583 8483
rect 27890 8480 27896 8492
rect 27571 8452 27896 8480
rect 27571 8449 27583 8452
rect 27525 8443 27583 8449
rect 27890 8440 27896 8452
rect 27948 8440 27954 8492
rect 29178 8440 29184 8492
rect 29236 8480 29242 8492
rect 29273 8483 29331 8489
rect 29273 8480 29285 8483
rect 29236 8452 29285 8480
rect 29236 8440 29242 8452
rect 29273 8449 29285 8452
rect 29319 8449 29331 8483
rect 29273 8443 29331 8449
rect 29365 8483 29423 8489
rect 29365 8449 29377 8483
rect 29411 8480 29423 8483
rect 29638 8480 29644 8492
rect 29411 8452 29644 8480
rect 29411 8449 29423 8452
rect 29365 8443 29423 8449
rect 29638 8440 29644 8452
rect 29696 8480 29702 8492
rect 30190 8480 30196 8492
rect 29696 8452 30196 8480
rect 29696 8440 29702 8452
rect 30190 8440 30196 8452
rect 30248 8440 30254 8492
rect 30926 8480 30932 8492
rect 30887 8452 30932 8480
rect 30926 8440 30932 8452
rect 30984 8440 30990 8492
rect 31036 8489 31064 8520
rect 33781 8517 33793 8551
rect 33827 8548 33839 8551
rect 33870 8548 33876 8560
rect 33827 8520 33876 8548
rect 33827 8517 33839 8520
rect 33781 8511 33839 8517
rect 33870 8508 33876 8520
rect 33928 8508 33934 8560
rect 31021 8483 31079 8489
rect 31021 8449 31033 8483
rect 31067 8480 31079 8483
rect 32674 8480 32680 8492
rect 31067 8452 32680 8480
rect 31067 8449 31079 8452
rect 31021 8443 31079 8449
rect 32674 8440 32680 8452
rect 32732 8440 32738 8492
rect 32858 8480 32864 8492
rect 32819 8452 32864 8480
rect 32858 8440 32864 8452
rect 32916 8440 32922 8492
rect 33962 8480 33968 8492
rect 33923 8452 33968 8480
rect 33962 8440 33968 8452
rect 34020 8440 34026 8492
rect 35060 8483 35118 8489
rect 35060 8449 35072 8483
rect 35106 8480 35118 8483
rect 35342 8480 35348 8492
rect 35106 8452 35348 8480
rect 35106 8449 35118 8452
rect 35060 8443 35118 8449
rect 35342 8440 35348 8452
rect 35400 8440 35406 8492
rect 25682 8372 25688 8424
rect 25740 8412 25746 8424
rect 26510 8412 26516 8424
rect 25740 8384 26516 8412
rect 25740 8372 25746 8384
rect 26510 8372 26516 8384
rect 26568 8412 26574 8424
rect 27709 8415 27767 8421
rect 27709 8412 27721 8415
rect 26568 8384 27721 8412
rect 26568 8372 26574 8384
rect 27709 8381 27721 8384
rect 27755 8381 27767 8415
rect 27709 8375 27767 8381
rect 22373 8347 22431 8353
rect 22373 8344 22385 8347
rect 20036 8316 20484 8344
rect 20548 8316 21220 8344
rect 21468 8316 22385 8344
rect 20036 8304 20042 8316
rect 14182 8276 14188 8288
rect 14143 8248 14188 8276
rect 14182 8236 14188 8248
rect 14240 8236 14246 8288
rect 18690 8236 18696 8288
rect 18748 8276 18754 8288
rect 18785 8279 18843 8285
rect 18785 8276 18797 8279
rect 18748 8248 18797 8276
rect 18748 8236 18754 8248
rect 18785 8245 18797 8248
rect 18831 8245 18843 8279
rect 20456 8276 20484 8316
rect 21468 8276 21496 8316
rect 22373 8313 22385 8316
rect 22419 8313 22431 8347
rect 27724 8344 27752 8375
rect 28350 8372 28356 8424
rect 28408 8412 28414 8424
rect 29089 8415 29147 8421
rect 29089 8412 29101 8415
rect 28408 8384 29101 8412
rect 28408 8372 28414 8384
rect 29089 8381 29101 8384
rect 29135 8412 29147 8415
rect 30944 8412 30972 8440
rect 29135 8384 30972 8412
rect 29135 8381 29147 8384
rect 29089 8375 29147 8381
rect 31386 8372 31392 8424
rect 31444 8412 31450 8424
rect 31846 8412 31852 8424
rect 31444 8384 31852 8412
rect 31444 8372 31450 8384
rect 31846 8372 31852 8384
rect 31904 8372 31910 8424
rect 33045 8415 33103 8421
rect 33045 8381 33057 8415
rect 33091 8381 33103 8415
rect 34790 8412 34796 8424
rect 34751 8384 34796 8412
rect 33045 8375 33103 8381
rect 29546 8344 29552 8356
rect 27724 8316 29552 8344
rect 22373 8307 22431 8313
rect 29546 8304 29552 8316
rect 29604 8344 29610 8356
rect 33060 8344 33088 8375
rect 34790 8372 34796 8384
rect 34848 8372 34854 8424
rect 37918 8412 37924 8424
rect 37879 8384 37924 8412
rect 37918 8372 37924 8384
rect 37976 8372 37982 8424
rect 38105 8415 38163 8421
rect 38105 8381 38117 8415
rect 38151 8412 38163 8415
rect 38194 8412 38200 8424
rect 38151 8384 38200 8412
rect 38151 8381 38163 8384
rect 38105 8375 38163 8381
rect 38194 8372 38200 8384
rect 38252 8372 38258 8424
rect 29604 8316 33088 8344
rect 34149 8347 34207 8353
rect 29604 8304 29610 8316
rect 34149 8313 34161 8347
rect 34195 8344 34207 8347
rect 34606 8344 34612 8356
rect 34195 8316 34612 8344
rect 34195 8313 34207 8316
rect 34149 8307 34207 8313
rect 34606 8304 34612 8316
rect 34664 8304 34670 8356
rect 37182 8304 37188 8356
rect 37240 8344 37246 8356
rect 37461 8347 37519 8353
rect 37461 8344 37473 8347
rect 37240 8316 37473 8344
rect 37240 8304 37246 8316
rect 37461 8313 37473 8316
rect 37507 8313 37519 8347
rect 37461 8307 37519 8313
rect 27154 8276 27160 8288
rect 20456 8248 21496 8276
rect 27115 8248 27160 8276
rect 18785 8239 18843 8245
rect 27154 8236 27160 8248
rect 27212 8236 27218 8288
rect 32490 8276 32496 8288
rect 32451 8248 32496 8276
rect 32490 8236 32496 8248
rect 32548 8236 32554 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 11790 8072 11796 8084
rect 11751 8044 11796 8072
rect 11790 8032 11796 8044
rect 11848 8032 11854 8084
rect 12802 8072 12808 8084
rect 12763 8044 12808 8072
rect 12802 8032 12808 8044
rect 12860 8032 12866 8084
rect 15562 8072 15568 8084
rect 15523 8044 15568 8072
rect 15562 8032 15568 8044
rect 15620 8032 15626 8084
rect 16666 8032 16672 8084
rect 16724 8072 16730 8084
rect 17589 8075 17647 8081
rect 17589 8072 17601 8075
rect 16724 8044 17601 8072
rect 16724 8032 16730 8044
rect 17589 8041 17601 8044
rect 17635 8041 17647 8075
rect 17589 8035 17647 8041
rect 18782 8032 18788 8084
rect 18840 8072 18846 8084
rect 20898 8072 20904 8084
rect 18840 8044 20904 8072
rect 18840 8032 18846 8044
rect 20898 8032 20904 8044
rect 20956 8032 20962 8084
rect 23014 8072 23020 8084
rect 22975 8044 23020 8072
rect 23014 8032 23020 8044
rect 23072 8032 23078 8084
rect 27890 8072 27896 8084
rect 27851 8044 27896 8072
rect 27890 8032 27896 8044
rect 27948 8032 27954 8084
rect 28721 8075 28779 8081
rect 28721 8041 28733 8075
rect 28767 8072 28779 8075
rect 29822 8072 29828 8084
rect 28767 8044 29828 8072
rect 28767 8041 28779 8044
rect 28721 8035 28779 8041
rect 29822 8032 29828 8044
rect 29880 8032 29886 8084
rect 32033 8075 32091 8081
rect 32033 8041 32045 8075
rect 32079 8072 32091 8075
rect 32858 8072 32864 8084
rect 32079 8044 32864 8072
rect 32079 8041 32091 8044
rect 32033 8035 32091 8041
rect 32858 8032 32864 8044
rect 32916 8032 32922 8084
rect 35069 8075 35127 8081
rect 35069 8041 35081 8075
rect 35115 8072 35127 8075
rect 35342 8072 35348 8084
rect 35115 8044 35348 8072
rect 35115 8041 35127 8044
rect 35069 8035 35127 8041
rect 35342 8032 35348 8044
rect 35400 8032 35406 8084
rect 37826 8032 37832 8084
rect 37884 8072 37890 8084
rect 38289 8075 38347 8081
rect 38289 8072 38301 8075
rect 37884 8044 38301 8072
rect 37884 8032 37890 8044
rect 38289 8041 38301 8044
rect 38335 8041 38347 8075
rect 38289 8035 38347 8041
rect 31662 7964 31668 8016
rect 31720 7964 31726 8016
rect 34422 7964 34428 8016
rect 34480 8004 34486 8016
rect 34480 7976 35664 8004
rect 34480 7964 34486 7976
rect 14826 7936 14832 7948
rect 12268 7908 12940 7936
rect 12268 7880 12296 7908
rect 11977 7871 12035 7877
rect 11977 7837 11989 7871
rect 12023 7837 12035 7871
rect 12250 7868 12256 7880
rect 12211 7840 12256 7868
rect 11977 7831 12035 7837
rect 11992 7800 12020 7831
rect 12250 7828 12256 7840
rect 12308 7828 12314 7880
rect 12710 7868 12716 7880
rect 12406 7840 12716 7868
rect 12406 7800 12434 7840
rect 12710 7828 12716 7840
rect 12768 7828 12774 7880
rect 12912 7812 12940 7908
rect 14292 7908 14832 7936
rect 12989 7871 13047 7877
rect 12989 7837 13001 7871
rect 13035 7868 13047 7871
rect 14182 7868 14188 7880
rect 13035 7840 14188 7868
rect 13035 7837 13047 7840
rect 12989 7831 13047 7837
rect 12894 7800 12900 7812
rect 11992 7772 12434 7800
rect 12855 7772 12900 7800
rect 12894 7760 12900 7772
rect 12952 7760 12958 7812
rect 12161 7735 12219 7741
rect 12161 7701 12173 7735
rect 12207 7732 12219 7735
rect 13004 7732 13032 7831
rect 14182 7828 14188 7840
rect 14240 7828 14246 7880
rect 14292 7877 14320 7908
rect 14826 7896 14832 7908
rect 14884 7896 14890 7948
rect 18509 7939 18567 7945
rect 16408 7908 17448 7936
rect 14277 7871 14335 7877
rect 14277 7837 14289 7871
rect 14323 7837 14335 7871
rect 14918 7868 14924 7880
rect 14879 7840 14924 7868
rect 14277 7831 14335 7837
rect 14918 7828 14924 7840
rect 14976 7828 14982 7880
rect 16298 7828 16304 7880
rect 16356 7868 16362 7880
rect 16408 7877 16436 7908
rect 16393 7871 16451 7877
rect 16393 7868 16405 7871
rect 16356 7840 16405 7868
rect 16356 7828 16362 7840
rect 16393 7837 16405 7840
rect 16439 7837 16451 7871
rect 16393 7831 16451 7837
rect 16482 7828 16488 7880
rect 16540 7868 16546 7880
rect 16666 7868 16672 7880
rect 16540 7840 16585 7868
rect 16627 7840 16672 7868
rect 16540 7828 16546 7840
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 16761 7871 16819 7877
rect 16761 7837 16773 7871
rect 16807 7868 16819 7871
rect 16850 7868 16856 7880
rect 16807 7840 16856 7868
rect 16807 7837 16819 7840
rect 16761 7831 16819 7837
rect 16850 7828 16856 7840
rect 16908 7828 16914 7880
rect 17420 7877 17448 7908
rect 18509 7905 18521 7939
rect 18555 7936 18567 7939
rect 18598 7936 18604 7948
rect 18555 7908 18604 7936
rect 18555 7905 18567 7908
rect 18509 7899 18567 7905
rect 18598 7896 18604 7908
rect 18656 7896 18662 7948
rect 20622 7896 20628 7948
rect 20680 7936 20686 7948
rect 31680 7936 31708 7964
rect 35250 7936 35256 7948
rect 20680 7908 20760 7936
rect 31680 7908 35256 7936
rect 20680 7896 20686 7908
rect 17405 7871 17463 7877
rect 17405 7837 17417 7871
rect 17451 7837 17463 7871
rect 17405 7831 17463 7837
rect 17681 7871 17739 7877
rect 17681 7837 17693 7871
rect 17727 7837 17739 7871
rect 18414 7868 18420 7880
rect 18375 7840 18420 7868
rect 17681 7831 17739 7837
rect 14734 7800 14740 7812
rect 14695 7772 14740 7800
rect 14734 7760 14740 7772
rect 14792 7760 14798 7812
rect 16868 7800 16896 7828
rect 17696 7800 17724 7831
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 18690 7868 18696 7880
rect 18651 7840 18696 7868
rect 18690 7828 18696 7840
rect 18748 7828 18754 7880
rect 19521 7871 19579 7877
rect 19521 7837 19533 7871
rect 19567 7837 19579 7871
rect 19521 7831 19579 7837
rect 19613 7871 19671 7877
rect 19613 7837 19625 7871
rect 19659 7868 19671 7871
rect 20441 7871 20499 7877
rect 20441 7868 20453 7871
rect 19659 7840 20453 7868
rect 19659 7837 19671 7840
rect 19613 7831 19671 7837
rect 20441 7837 20453 7840
rect 20487 7837 20499 7871
rect 20441 7831 20499 7837
rect 16868 7772 17724 7800
rect 19536 7800 19564 7831
rect 20530 7828 20536 7880
rect 20588 7868 20594 7880
rect 20732 7877 20760 7908
rect 35250 7896 35256 7908
rect 35308 7896 35314 7948
rect 35342 7896 35348 7948
rect 35400 7936 35406 7948
rect 35526 7936 35532 7948
rect 35400 7908 35532 7936
rect 35400 7896 35406 7908
rect 35526 7896 35532 7908
rect 35584 7896 35590 7948
rect 35636 7945 35664 7976
rect 35621 7939 35679 7945
rect 35621 7905 35633 7939
rect 35667 7905 35679 7939
rect 35621 7899 35679 7905
rect 20717 7871 20775 7877
rect 20588 7840 20633 7868
rect 20588 7828 20594 7840
rect 20717 7837 20729 7871
rect 20763 7837 20775 7871
rect 20717 7831 20775 7837
rect 21637 7871 21695 7877
rect 21637 7837 21649 7871
rect 21683 7868 21695 7871
rect 22462 7868 22468 7880
rect 21683 7840 22468 7868
rect 21683 7837 21695 7840
rect 21637 7831 21695 7837
rect 22462 7828 22468 7840
rect 22520 7828 22526 7880
rect 26513 7871 26571 7877
rect 26513 7837 26525 7871
rect 26559 7868 26571 7871
rect 26602 7868 26608 7880
rect 26559 7840 26608 7868
rect 26559 7837 26571 7840
rect 26513 7831 26571 7837
rect 26602 7828 26608 7840
rect 26660 7828 26666 7880
rect 26780 7871 26838 7877
rect 26780 7837 26792 7871
rect 26826 7868 26838 7871
rect 27154 7868 27160 7880
rect 26826 7840 27160 7868
rect 26826 7837 26838 7840
rect 26780 7831 26838 7837
rect 27154 7828 27160 7840
rect 27212 7828 27218 7880
rect 27890 7828 27896 7880
rect 27948 7868 27954 7880
rect 28537 7871 28595 7877
rect 28537 7868 28549 7871
rect 27948 7840 28549 7868
rect 27948 7828 27954 7840
rect 28537 7837 28549 7840
rect 28583 7837 28595 7871
rect 28537 7831 28595 7837
rect 30653 7871 30711 7877
rect 30653 7837 30665 7871
rect 30699 7868 30711 7871
rect 31202 7868 31208 7880
rect 30699 7840 31208 7868
rect 30699 7837 30711 7840
rect 30653 7831 30711 7837
rect 31202 7828 31208 7840
rect 31260 7868 31266 7880
rect 31662 7868 31668 7880
rect 31260 7840 31668 7868
rect 31260 7828 31266 7840
rect 31662 7828 31668 7840
rect 31720 7868 31726 7880
rect 33226 7868 33232 7880
rect 31720 7840 33088 7868
rect 33187 7840 33232 7868
rect 31720 7828 31726 7840
rect 20806 7800 20812 7812
rect 19536 7772 20812 7800
rect 20806 7760 20812 7772
rect 20864 7760 20870 7812
rect 21177 7803 21235 7809
rect 21177 7769 21189 7803
rect 21223 7769 21235 7803
rect 21177 7763 21235 7769
rect 16206 7732 16212 7744
rect 12207 7704 13032 7732
rect 16167 7704 16212 7732
rect 12207 7701 12219 7704
rect 12161 7695 12219 7701
rect 16206 7692 16212 7704
rect 16264 7692 16270 7744
rect 16574 7692 16580 7744
rect 16632 7732 16638 7744
rect 17221 7735 17279 7741
rect 17221 7732 17233 7735
rect 16632 7704 17233 7732
rect 16632 7692 16638 7704
rect 17221 7701 17233 7704
rect 17267 7701 17279 7735
rect 17221 7695 17279 7701
rect 20254 7692 20260 7744
rect 20312 7732 20318 7744
rect 21192 7732 21220 7763
rect 21726 7760 21732 7812
rect 21784 7800 21790 7812
rect 21882 7803 21940 7809
rect 21882 7800 21894 7803
rect 21784 7772 21894 7800
rect 21784 7760 21790 7772
rect 21882 7769 21894 7772
rect 21928 7769 21940 7803
rect 28350 7800 28356 7812
rect 28311 7772 28356 7800
rect 21882 7763 21940 7769
rect 28350 7760 28356 7772
rect 28408 7760 28414 7812
rect 30920 7803 30978 7809
rect 30920 7769 30932 7803
rect 30966 7800 30978 7803
rect 32490 7800 32496 7812
rect 30966 7772 32496 7800
rect 30966 7769 30978 7772
rect 30920 7763 30978 7769
rect 32490 7760 32496 7772
rect 32548 7760 32554 7812
rect 33060 7800 33088 7840
rect 33226 7828 33232 7840
rect 33284 7828 33290 7880
rect 36722 7868 36728 7880
rect 34808 7840 35204 7868
rect 34808 7812 34836 7840
rect 33965 7803 34023 7809
rect 33965 7800 33977 7803
rect 33060 7772 33977 7800
rect 33965 7769 33977 7772
rect 34011 7800 34023 7803
rect 34790 7800 34796 7812
rect 34011 7772 34796 7800
rect 34011 7769 34023 7772
rect 33965 7763 34023 7769
rect 34790 7760 34796 7772
rect 34848 7760 34854 7812
rect 35176 7800 35204 7840
rect 35360 7840 36728 7868
rect 35360 7800 35388 7840
rect 36722 7828 36728 7840
rect 36780 7868 36786 7880
rect 37182 7877 37188 7880
rect 36909 7871 36967 7877
rect 36909 7868 36921 7871
rect 36780 7840 36921 7868
rect 36780 7828 36786 7840
rect 36909 7837 36921 7840
rect 36955 7837 36967 7871
rect 37176 7868 37188 7877
rect 37143 7840 37188 7868
rect 36909 7831 36967 7837
rect 37176 7831 37188 7840
rect 37182 7828 37188 7831
rect 37240 7828 37246 7880
rect 35176 7772 35388 7800
rect 35437 7803 35495 7809
rect 35437 7769 35449 7803
rect 35483 7800 35495 7803
rect 36078 7800 36084 7812
rect 35483 7772 36084 7800
rect 35483 7769 35495 7772
rect 35437 7763 35495 7769
rect 36078 7760 36084 7772
rect 36136 7760 36142 7812
rect 20312 7704 21220 7732
rect 20312 7692 20318 7704
rect 34606 7692 34612 7744
rect 34664 7732 34670 7744
rect 35158 7732 35164 7744
rect 34664 7704 35164 7732
rect 34664 7692 34670 7704
rect 35158 7692 35164 7704
rect 35216 7692 35222 7744
rect 35250 7692 35256 7744
rect 35308 7732 35314 7744
rect 35529 7735 35587 7741
rect 35529 7732 35541 7735
rect 35308 7704 35541 7732
rect 35308 7692 35314 7704
rect 35529 7701 35541 7704
rect 35575 7732 35587 7735
rect 35894 7732 35900 7744
rect 35575 7704 35900 7732
rect 35575 7701 35587 7704
rect 35529 7695 35587 7701
rect 35894 7692 35900 7704
rect 35952 7732 35958 7744
rect 37918 7732 37924 7744
rect 35952 7704 37924 7732
rect 35952 7692 35958 7704
rect 37918 7692 37924 7704
rect 37976 7692 37982 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 20530 7488 20536 7540
rect 20588 7528 20594 7540
rect 21453 7531 21511 7537
rect 21453 7528 21465 7531
rect 20588 7500 21465 7528
rect 20588 7488 20594 7500
rect 21453 7497 21465 7500
rect 21499 7497 21511 7531
rect 21453 7491 21511 7497
rect 22554 7488 22560 7540
rect 22612 7528 22618 7540
rect 24229 7531 24287 7537
rect 24229 7528 24241 7531
rect 22612 7500 24241 7528
rect 22612 7488 22618 7500
rect 24229 7497 24241 7500
rect 24275 7528 24287 7531
rect 26050 7528 26056 7540
rect 24275 7500 26056 7528
rect 24275 7497 24287 7500
rect 24229 7491 24287 7497
rect 26050 7488 26056 7500
rect 26108 7488 26114 7540
rect 33781 7531 33839 7537
rect 33781 7497 33793 7531
rect 33827 7528 33839 7531
rect 33962 7528 33968 7540
rect 33827 7500 33968 7528
rect 33827 7497 33839 7500
rect 33781 7491 33839 7497
rect 33962 7488 33968 7500
rect 34020 7488 34026 7540
rect 34514 7528 34520 7540
rect 34475 7500 34520 7528
rect 34514 7488 34520 7500
rect 34572 7488 34578 7540
rect 37826 7528 37832 7540
rect 34808 7500 37832 7528
rect 13354 7460 13360 7472
rect 13315 7432 13360 7460
rect 13354 7420 13360 7432
rect 13412 7420 13418 7472
rect 15930 7460 15936 7472
rect 14108 7432 15936 7460
rect 11701 7395 11759 7401
rect 11701 7361 11713 7395
rect 11747 7392 11759 7395
rect 12986 7392 12992 7404
rect 11747 7364 12992 7392
rect 11747 7361 11759 7364
rect 11701 7355 11759 7361
rect 12986 7352 12992 7364
rect 13044 7392 13050 7404
rect 14108 7392 14136 7432
rect 15930 7420 15936 7432
rect 15988 7420 15994 7472
rect 18690 7460 18696 7472
rect 17236 7432 18696 7460
rect 14366 7392 14372 7404
rect 13044 7364 14136 7392
rect 14327 7364 14372 7392
rect 13044 7352 13050 7364
rect 14366 7352 14372 7364
rect 14424 7352 14430 7404
rect 14458 7352 14464 7404
rect 14516 7392 14522 7404
rect 14734 7392 14740 7404
rect 14516 7364 14561 7392
rect 14695 7364 14740 7392
rect 14516 7352 14522 7364
rect 14734 7352 14740 7364
rect 14792 7352 14798 7404
rect 17236 7401 17264 7432
rect 18690 7420 18696 7432
rect 18748 7460 18754 7472
rect 18748 7432 19104 7460
rect 18748 7420 18754 7432
rect 14921 7395 14979 7401
rect 14921 7361 14933 7395
rect 14967 7361 14979 7395
rect 14921 7355 14979 7361
rect 17221 7395 17279 7401
rect 17221 7361 17233 7395
rect 17267 7361 17279 7395
rect 17221 7355 17279 7361
rect 17405 7395 17463 7401
rect 17405 7361 17417 7395
rect 17451 7392 17463 7395
rect 18509 7395 18567 7401
rect 18509 7392 18521 7395
rect 17451 7364 18521 7392
rect 17451 7361 17463 7364
rect 17405 7355 17463 7361
rect 18509 7361 18521 7364
rect 18555 7392 18567 7395
rect 18598 7392 18604 7404
rect 18555 7364 18604 7392
rect 18555 7361 18567 7364
rect 18509 7355 18567 7361
rect 11974 7324 11980 7336
rect 11935 7296 11980 7324
rect 11974 7284 11980 7296
rect 12032 7284 12038 7336
rect 14182 7284 14188 7336
rect 14240 7324 14246 7336
rect 14936 7324 14964 7355
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 19076 7401 19104 7432
rect 20806 7420 20812 7472
rect 20864 7460 20870 7472
rect 21085 7463 21143 7469
rect 21085 7460 21097 7463
rect 20864 7432 21097 7460
rect 20864 7420 20870 7432
rect 21085 7429 21097 7432
rect 21131 7429 21143 7463
rect 24026 7460 24032 7472
rect 23987 7432 24032 7460
rect 21085 7423 21143 7429
rect 24026 7420 24032 7432
rect 24084 7420 24090 7472
rect 29178 7420 29184 7472
rect 29236 7460 29242 7472
rect 29549 7463 29607 7469
rect 29549 7460 29561 7463
rect 29236 7432 29561 7460
rect 29236 7420 29242 7432
rect 29549 7429 29561 7432
rect 29595 7429 29607 7463
rect 29549 7423 29607 7429
rect 19061 7395 19119 7401
rect 19061 7361 19073 7395
rect 19107 7361 19119 7395
rect 20254 7392 20260 7404
rect 20167 7364 20260 7392
rect 19061 7355 19119 7361
rect 20254 7352 20260 7364
rect 20312 7352 20318 7404
rect 20349 7395 20407 7401
rect 20349 7361 20361 7395
rect 20395 7361 20407 7395
rect 20622 7392 20628 7404
rect 20583 7364 20628 7392
rect 20349 7355 20407 7361
rect 14240 7296 14964 7324
rect 17497 7327 17555 7333
rect 14240 7284 14246 7296
rect 17497 7293 17509 7327
rect 17543 7324 17555 7327
rect 18138 7324 18144 7336
rect 17543 7296 18144 7324
rect 17543 7293 17555 7296
rect 17497 7287 17555 7293
rect 18138 7284 18144 7296
rect 18196 7284 18202 7336
rect 18782 7324 18788 7336
rect 18743 7296 18788 7324
rect 18782 7284 18788 7296
rect 18840 7324 18846 7336
rect 20272 7324 20300 7352
rect 18840 7296 20300 7324
rect 18840 7284 18846 7296
rect 12894 7216 12900 7268
rect 12952 7256 12958 7268
rect 14553 7259 14611 7265
rect 14553 7256 14565 7259
rect 12952 7228 14565 7256
rect 12952 7216 12958 7228
rect 14553 7225 14565 7228
rect 14599 7225 14611 7259
rect 14553 7219 14611 7225
rect 17954 7216 17960 7268
rect 18012 7256 18018 7268
rect 18693 7259 18751 7265
rect 18693 7256 18705 7259
rect 18012 7228 18705 7256
rect 18012 7216 18018 7228
rect 18693 7225 18705 7228
rect 18739 7225 18751 7259
rect 20364 7256 20392 7355
rect 20622 7352 20628 7364
rect 20680 7352 20686 7404
rect 20533 7327 20591 7333
rect 20533 7293 20545 7327
rect 20579 7324 20591 7327
rect 20824 7324 20852 7420
rect 20898 7352 20904 7404
rect 20956 7392 20962 7404
rect 21269 7395 21327 7401
rect 21269 7392 21281 7395
rect 20956 7364 21281 7392
rect 20956 7352 20962 7364
rect 21269 7361 21281 7364
rect 21315 7361 21327 7395
rect 21269 7355 21327 7361
rect 29638 7352 29644 7404
rect 29696 7392 29702 7404
rect 29696 7364 29741 7392
rect 29696 7352 29702 7364
rect 31662 7352 31668 7404
rect 31720 7392 31726 7404
rect 32401 7395 32459 7401
rect 32401 7392 32413 7395
rect 31720 7364 32413 7392
rect 31720 7352 31726 7364
rect 32401 7361 32413 7364
rect 32447 7361 32459 7395
rect 32401 7355 32459 7361
rect 32668 7395 32726 7401
rect 32668 7361 32680 7395
rect 32714 7392 32726 7395
rect 32950 7392 32956 7404
rect 32714 7364 32956 7392
rect 32714 7361 32726 7364
rect 32668 7355 32726 7361
rect 32950 7352 32956 7364
rect 33008 7352 33014 7404
rect 34808 7401 34836 7500
rect 37826 7488 37832 7500
rect 37884 7488 37890 7540
rect 37921 7531 37979 7537
rect 37921 7497 37933 7531
rect 37967 7528 37979 7531
rect 38010 7528 38016 7540
rect 37967 7500 38016 7528
rect 37967 7497 37979 7500
rect 37921 7491 37979 7497
rect 38010 7488 38016 7500
rect 38068 7488 38074 7540
rect 34793 7395 34851 7401
rect 34793 7361 34805 7395
rect 34839 7361 34851 7395
rect 34793 7355 34851 7361
rect 34885 7395 34943 7401
rect 34885 7361 34897 7395
rect 34931 7361 34943 7395
rect 34885 7355 34943 7361
rect 34977 7395 35035 7401
rect 34977 7361 34989 7395
rect 35023 7392 35035 7395
rect 35066 7392 35072 7404
rect 35023 7364 35072 7392
rect 35023 7361 35035 7364
rect 34977 7355 35035 7361
rect 20579 7296 20852 7324
rect 20579 7293 20591 7296
rect 20533 7287 20591 7293
rect 18693 7219 18751 7225
rect 18800 7228 20392 7256
rect 17037 7191 17095 7197
rect 17037 7157 17049 7191
rect 17083 7188 17095 7191
rect 18230 7188 18236 7200
rect 17083 7160 18236 7188
rect 17083 7157 17095 7160
rect 17037 7151 17095 7157
rect 18230 7148 18236 7160
rect 18288 7188 18294 7200
rect 18800 7188 18828 7228
rect 20070 7188 20076 7200
rect 18288 7160 18828 7188
rect 20031 7160 20076 7188
rect 18288 7148 18294 7160
rect 20070 7148 20076 7160
rect 20128 7148 20134 7200
rect 24210 7188 24216 7200
rect 24171 7160 24216 7188
rect 24210 7148 24216 7160
rect 24268 7148 24274 7200
rect 24394 7188 24400 7200
rect 24355 7160 24400 7188
rect 24394 7148 24400 7160
rect 24452 7148 24458 7200
rect 29086 7148 29092 7200
rect 29144 7188 29150 7200
rect 29365 7191 29423 7197
rect 29365 7188 29377 7191
rect 29144 7160 29377 7188
rect 29144 7148 29150 7160
rect 29365 7157 29377 7160
rect 29411 7157 29423 7191
rect 29365 7151 29423 7157
rect 29546 7148 29552 7200
rect 29604 7188 29610 7200
rect 29825 7191 29883 7197
rect 29825 7188 29837 7191
rect 29604 7160 29837 7188
rect 29604 7148 29610 7160
rect 29825 7157 29837 7160
rect 29871 7157 29883 7191
rect 29825 7151 29883 7157
rect 31018 7148 31024 7200
rect 31076 7188 31082 7200
rect 31938 7188 31944 7200
rect 31076 7160 31944 7188
rect 31076 7148 31082 7160
rect 31938 7148 31944 7160
rect 31996 7188 32002 7200
rect 34790 7188 34796 7200
rect 31996 7160 34796 7188
rect 31996 7148 32002 7160
rect 34790 7148 34796 7160
rect 34848 7188 34854 7200
rect 34900 7188 34928 7355
rect 35066 7352 35072 7364
rect 35124 7352 35130 7404
rect 35158 7352 35164 7404
rect 35216 7392 35222 7404
rect 35216 7364 35261 7392
rect 35216 7352 35222 7364
rect 38010 7324 38016 7336
rect 37971 7296 38016 7324
rect 38010 7284 38016 7296
rect 38068 7284 38074 7336
rect 34848 7160 34928 7188
rect 34848 7148 34854 7160
rect 36998 7148 37004 7200
rect 37056 7188 37062 7200
rect 37461 7191 37519 7197
rect 37461 7188 37473 7191
rect 37056 7160 37473 7188
rect 37056 7148 37062 7160
rect 37461 7157 37473 7160
rect 37507 7157 37519 7191
rect 37461 7151 37519 7157
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 14458 6944 14464 6996
rect 14516 6984 14522 6996
rect 21637 6987 21695 6993
rect 14516 6956 14872 6984
rect 14516 6944 14522 6956
rect 14277 6919 14335 6925
rect 14277 6916 14289 6919
rect 13372 6888 14289 6916
rect 11974 6808 11980 6860
rect 12032 6848 12038 6860
rect 12529 6851 12587 6857
rect 12529 6848 12541 6851
rect 12032 6820 12541 6848
rect 12032 6808 12038 6820
rect 12529 6817 12541 6820
rect 12575 6817 12587 6851
rect 12529 6811 12587 6817
rect 12250 6780 12256 6792
rect 12211 6752 12256 6780
rect 12250 6740 12256 6752
rect 12308 6740 12314 6792
rect 12345 6783 12403 6789
rect 12345 6749 12357 6783
rect 12391 6780 12403 6783
rect 13372 6780 13400 6888
rect 14277 6885 14289 6888
rect 14323 6885 14335 6919
rect 14277 6879 14335 6885
rect 14734 6876 14740 6928
rect 14792 6876 14798 6928
rect 14752 6848 14780 6876
rect 14476 6820 14780 6848
rect 14476 6789 14504 6820
rect 12391 6752 13400 6780
rect 14461 6783 14519 6789
rect 12391 6749 12403 6752
rect 12345 6743 12403 6749
rect 14461 6749 14473 6783
rect 14507 6749 14519 6783
rect 14461 6743 14519 6749
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6749 14611 6783
rect 14734 6780 14740 6792
rect 14695 6752 14740 6780
rect 14553 6743 14611 6749
rect 14182 6672 14188 6724
rect 14240 6712 14246 6724
rect 14568 6712 14596 6743
rect 14734 6740 14740 6752
rect 14792 6740 14798 6792
rect 14844 6789 14872 6956
rect 21637 6953 21649 6987
rect 21683 6984 21695 6987
rect 21726 6984 21732 6996
rect 21683 6956 21732 6984
rect 21683 6953 21695 6956
rect 21637 6947 21695 6953
rect 21726 6944 21732 6956
rect 21784 6944 21790 6996
rect 23845 6987 23903 6993
rect 23845 6953 23857 6987
rect 23891 6984 23903 6987
rect 24026 6984 24032 6996
rect 23891 6956 24032 6984
rect 23891 6953 23903 6956
rect 23845 6947 23903 6953
rect 24026 6944 24032 6956
rect 24084 6944 24090 6996
rect 25130 6984 25136 6996
rect 25091 6956 25136 6984
rect 25130 6944 25136 6956
rect 25188 6944 25194 6996
rect 32950 6984 32956 6996
rect 32911 6956 32956 6984
rect 32950 6944 32956 6956
rect 33008 6944 33014 6996
rect 34885 6987 34943 6993
rect 34885 6953 34897 6987
rect 34931 6984 34943 6987
rect 35434 6984 35440 6996
rect 34931 6956 35440 6984
rect 34931 6953 34943 6956
rect 34885 6947 34943 6953
rect 35434 6944 35440 6956
rect 35492 6944 35498 6996
rect 37826 6944 37832 6996
rect 37884 6984 37890 6996
rect 38105 6987 38163 6993
rect 38105 6984 38117 6987
rect 37884 6956 38117 6984
rect 37884 6944 37890 6956
rect 38105 6953 38117 6956
rect 38151 6953 38163 6987
rect 38105 6947 38163 6953
rect 26050 6876 26056 6928
rect 26108 6916 26114 6928
rect 26108 6888 27743 6916
rect 26108 6876 26114 6888
rect 16206 6808 16212 6860
rect 16264 6848 16270 6860
rect 16301 6851 16359 6857
rect 16301 6848 16313 6851
rect 16264 6820 16313 6848
rect 16264 6808 16270 6820
rect 16301 6817 16313 6820
rect 16347 6817 16359 6851
rect 17954 6848 17960 6860
rect 17915 6820 17960 6848
rect 16301 6811 16359 6817
rect 17954 6808 17960 6820
rect 18012 6808 18018 6860
rect 18414 6848 18420 6860
rect 18064 6820 18420 6848
rect 14829 6783 14887 6789
rect 14829 6749 14841 6783
rect 14875 6749 14887 6783
rect 14829 6743 14887 6749
rect 15657 6783 15715 6789
rect 15657 6749 15669 6783
rect 15703 6749 15715 6783
rect 16022 6780 16028 6792
rect 15983 6752 16028 6780
rect 15657 6743 15715 6749
rect 14240 6684 14596 6712
rect 15672 6712 15700 6743
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 17402 6780 17408 6792
rect 17363 6752 17408 6780
rect 17402 6740 17408 6752
rect 17460 6740 17466 6792
rect 17681 6783 17739 6789
rect 17681 6749 17693 6783
rect 17727 6780 17739 6783
rect 18064 6780 18092 6820
rect 18414 6808 18420 6820
rect 18472 6808 18478 6860
rect 18509 6851 18567 6857
rect 18509 6817 18521 6851
rect 18555 6848 18567 6851
rect 20438 6848 20444 6860
rect 18555 6820 20444 6848
rect 18555 6817 18567 6820
rect 18509 6811 18567 6817
rect 20438 6808 20444 6820
rect 20496 6848 20502 6860
rect 20809 6851 20867 6857
rect 20809 6848 20821 6851
rect 20496 6820 20821 6848
rect 20496 6808 20502 6820
rect 20809 6817 20821 6820
rect 20855 6817 20867 6851
rect 20809 6811 20867 6817
rect 25685 6851 25743 6857
rect 25685 6817 25697 6851
rect 25731 6848 25743 6851
rect 25774 6848 25780 6860
rect 25731 6820 25780 6848
rect 25731 6817 25743 6820
rect 25685 6811 25743 6817
rect 17727 6752 18092 6780
rect 18233 6783 18291 6789
rect 17727 6749 17739 6752
rect 17681 6743 17739 6749
rect 18233 6749 18245 6783
rect 18279 6780 18291 6783
rect 18322 6780 18328 6792
rect 18279 6752 18328 6780
rect 18279 6749 18291 6752
rect 18233 6743 18291 6749
rect 18322 6740 18328 6752
rect 18380 6740 18386 6792
rect 19978 6780 19984 6792
rect 19939 6752 19984 6780
rect 19978 6740 19984 6752
rect 20036 6740 20042 6792
rect 20070 6740 20076 6792
rect 20128 6780 20134 6792
rect 20530 6780 20536 6792
rect 20128 6752 20536 6780
rect 20128 6740 20134 6752
rect 20530 6740 20536 6752
rect 20588 6740 20594 6792
rect 20824 6780 20852 6811
rect 25774 6808 25780 6820
rect 25832 6808 25838 6860
rect 26142 6808 26148 6860
rect 26200 6848 26206 6860
rect 27617 6851 27675 6857
rect 27617 6848 27629 6851
rect 26200 6820 27629 6848
rect 26200 6808 26206 6820
rect 27617 6817 27629 6820
rect 27663 6817 27675 6851
rect 27617 6811 27675 6817
rect 21545 6783 21603 6789
rect 21545 6780 21557 6783
rect 20824 6752 21557 6780
rect 21545 6749 21557 6752
rect 21591 6749 21603 6783
rect 21545 6743 21603 6749
rect 21729 6783 21787 6789
rect 21729 6749 21741 6783
rect 21775 6749 21787 6783
rect 22462 6780 22468 6792
rect 22375 6752 22468 6780
rect 21729 6743 21787 6749
rect 16574 6712 16580 6724
rect 15672 6684 16580 6712
rect 14240 6672 14246 6684
rect 16574 6672 16580 6684
rect 16632 6672 16638 6724
rect 18046 6712 18052 6724
rect 17144 6684 18052 6712
rect 15565 6647 15623 6653
rect 15565 6613 15577 6647
rect 15611 6644 15623 6647
rect 17144 6644 17172 6684
rect 18046 6672 18052 6684
rect 18104 6672 18110 6724
rect 20548 6712 20576 6740
rect 21744 6712 21772 6743
rect 22462 6740 22468 6752
rect 22520 6780 22526 6792
rect 23198 6780 23204 6792
rect 22520 6752 23204 6780
rect 22520 6740 22526 6752
rect 23198 6740 23204 6752
rect 23256 6740 23262 6792
rect 20548 6684 21772 6712
rect 22732 6715 22790 6721
rect 22732 6681 22744 6715
rect 22778 6712 22790 6715
rect 23290 6712 23296 6724
rect 22778 6684 23296 6712
rect 22778 6681 22790 6684
rect 22732 6675 22790 6681
rect 23290 6672 23296 6684
rect 23348 6672 23354 6724
rect 25406 6712 25412 6724
rect 25367 6684 25412 6712
rect 25406 6672 25412 6684
rect 25464 6672 25470 6724
rect 25792 6712 25820 6808
rect 26234 6780 26240 6792
rect 26195 6752 26240 6780
rect 26234 6740 26240 6752
rect 26292 6740 26298 6792
rect 27715 6789 27743 6888
rect 34146 6876 34152 6928
rect 34204 6916 34210 6928
rect 34204 6888 35296 6916
rect 34204 6876 34210 6888
rect 28169 6851 28227 6857
rect 28169 6817 28181 6851
rect 28215 6848 28227 6851
rect 28350 6848 28356 6860
rect 28215 6820 28356 6848
rect 28215 6817 28227 6820
rect 28169 6811 28227 6817
rect 28350 6808 28356 6820
rect 28408 6808 28414 6860
rect 29730 6808 29736 6860
rect 29788 6848 29794 6860
rect 29788 6820 30328 6848
rect 29788 6808 29794 6820
rect 27709 6783 27767 6789
rect 27709 6749 27721 6783
rect 27755 6749 27767 6783
rect 27709 6743 27767 6749
rect 29270 6740 29276 6792
rect 29328 6780 29334 6792
rect 30009 6783 30067 6789
rect 30009 6780 30021 6783
rect 29328 6752 30021 6780
rect 29328 6740 29334 6752
rect 30009 6749 30021 6752
rect 30055 6749 30067 6783
rect 30009 6743 30067 6749
rect 30098 6740 30104 6792
rect 30156 6780 30162 6792
rect 30300 6789 30328 6820
rect 30650 6808 30656 6860
rect 30708 6848 30714 6860
rect 30745 6851 30803 6857
rect 30745 6848 30757 6851
rect 30708 6820 30757 6848
rect 30708 6808 30714 6820
rect 30745 6817 30757 6820
rect 30791 6817 30803 6851
rect 30745 6811 30803 6817
rect 33042 6808 33048 6860
rect 33100 6848 33106 6860
rect 33505 6851 33563 6857
rect 33505 6848 33517 6851
rect 33100 6820 33517 6848
rect 33100 6808 33106 6820
rect 33505 6817 33517 6820
rect 33551 6817 33563 6851
rect 33505 6811 33563 6817
rect 30285 6783 30343 6789
rect 30156 6752 30201 6780
rect 30156 6740 30162 6752
rect 30285 6749 30297 6783
rect 30331 6780 30343 6783
rect 33321 6783 33379 6789
rect 30331 6752 31754 6780
rect 30331 6749 30343 6752
rect 30285 6743 30343 6749
rect 27065 6715 27123 6721
rect 25792 6684 27016 6712
rect 15611 6616 17172 6644
rect 15611 6613 15623 6616
rect 15565 6607 15623 6613
rect 18690 6604 18696 6656
rect 18748 6644 18754 6656
rect 20073 6647 20131 6653
rect 20073 6644 20085 6647
rect 18748 6616 20085 6644
rect 18748 6604 18754 6616
rect 20073 6613 20085 6616
rect 20119 6644 20131 6647
rect 21358 6644 21364 6656
rect 20119 6616 21364 6644
rect 20119 6613 20131 6616
rect 20073 6607 20131 6613
rect 21358 6604 21364 6616
rect 21416 6604 21422 6656
rect 25593 6647 25651 6653
rect 25593 6613 25605 6647
rect 25639 6644 25651 6647
rect 25958 6644 25964 6656
rect 25639 6616 25964 6644
rect 25639 6613 25651 6616
rect 25593 6607 25651 6613
rect 25958 6604 25964 6616
rect 26016 6604 26022 6656
rect 26988 6644 27016 6684
rect 27065 6681 27077 6715
rect 27111 6712 27123 6715
rect 27430 6712 27436 6724
rect 27111 6684 27436 6712
rect 27111 6681 27123 6684
rect 27065 6675 27123 6681
rect 27430 6672 27436 6684
rect 27488 6672 27494 6724
rect 31726 6712 31754 6752
rect 33321 6749 33333 6783
rect 33367 6780 33379 6783
rect 33962 6780 33968 6792
rect 33367 6752 33968 6780
rect 33367 6749 33379 6752
rect 33321 6743 33379 6749
rect 33962 6740 33968 6752
rect 34020 6740 34026 6792
rect 35066 6740 35072 6792
rect 35124 6789 35130 6792
rect 35268 6789 35296 6888
rect 36722 6848 36728 6860
rect 36683 6820 36728 6848
rect 36722 6808 36728 6820
rect 36780 6808 36786 6860
rect 35124 6783 35173 6789
rect 35124 6749 35127 6783
rect 35161 6749 35173 6783
rect 35124 6743 35173 6749
rect 35253 6783 35311 6789
rect 35253 6749 35265 6783
rect 35299 6749 35311 6783
rect 35253 6743 35311 6749
rect 35345 6783 35403 6789
rect 35345 6749 35357 6783
rect 35391 6749 35403 6783
rect 35526 6780 35532 6792
rect 35487 6752 35532 6780
rect 35345 6743 35403 6749
rect 35124 6740 35130 6743
rect 35360 6712 35388 6743
rect 35526 6740 35532 6752
rect 35584 6740 35590 6792
rect 36998 6789 37004 6792
rect 36992 6780 37004 6789
rect 36959 6752 37004 6780
rect 36992 6743 37004 6752
rect 36998 6740 37004 6743
rect 37056 6740 37062 6792
rect 31726 6684 35388 6712
rect 29178 6644 29184 6656
rect 26988 6616 29184 6644
rect 29178 6604 29184 6616
rect 29236 6604 29242 6656
rect 33318 6604 33324 6656
rect 33376 6644 33382 6656
rect 33413 6647 33471 6653
rect 33413 6644 33425 6647
rect 33376 6616 33425 6644
rect 33376 6604 33382 6616
rect 33413 6613 33425 6616
rect 33459 6613 33471 6647
rect 33413 6607 33471 6613
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 20438 6400 20444 6452
rect 20496 6440 20502 6452
rect 20549 6443 20607 6449
rect 20549 6440 20561 6443
rect 20496 6412 20561 6440
rect 20496 6400 20502 6412
rect 20549 6409 20561 6412
rect 20595 6409 20607 6443
rect 20549 6403 20607 6409
rect 20717 6443 20775 6449
rect 20717 6409 20729 6443
rect 20763 6409 20775 6443
rect 23290 6440 23296 6452
rect 23251 6412 23296 6440
rect 20717 6403 20775 6409
rect 18972 6384 19024 6390
rect 16574 6372 16580 6384
rect 15580 6344 16580 6372
rect 15580 6313 15608 6344
rect 16574 6332 16580 6344
rect 16632 6332 16638 6384
rect 18414 6332 18420 6384
rect 18472 6372 18478 6384
rect 18472 6344 18972 6372
rect 18472 6332 18478 6344
rect 19978 6332 19984 6384
rect 20036 6372 20042 6384
rect 20349 6375 20407 6381
rect 20349 6372 20361 6375
rect 20036 6344 20361 6372
rect 20036 6332 20042 6344
rect 20349 6341 20361 6344
rect 20395 6341 20407 6375
rect 20349 6335 20407 6341
rect 18972 6326 19024 6332
rect 15565 6307 15623 6313
rect 15565 6273 15577 6307
rect 15611 6273 15623 6307
rect 15565 6267 15623 6273
rect 16025 6307 16083 6313
rect 16025 6273 16037 6307
rect 16071 6304 16083 6307
rect 16206 6304 16212 6316
rect 16071 6276 16212 6304
rect 16071 6273 16083 6276
rect 16025 6267 16083 6273
rect 16206 6264 16212 6276
rect 16264 6264 16270 6316
rect 18138 6304 18144 6316
rect 18099 6276 18144 6304
rect 18138 6264 18144 6276
rect 18196 6264 18202 6316
rect 18598 6304 18604 6316
rect 18559 6276 18604 6304
rect 18598 6264 18604 6276
rect 18656 6264 18662 6316
rect 20732 6304 20760 6403
rect 23290 6400 23296 6412
rect 23348 6400 23354 6452
rect 23661 6443 23719 6449
rect 23661 6409 23673 6443
rect 23707 6440 23719 6443
rect 24026 6440 24032 6452
rect 23707 6412 24032 6440
rect 23707 6409 23719 6412
rect 23661 6403 23719 6409
rect 24026 6400 24032 6412
rect 24084 6400 24090 6452
rect 24587 6443 24645 6449
rect 24587 6409 24599 6443
rect 24633 6440 24645 6443
rect 25406 6440 25412 6452
rect 24633 6412 25412 6440
rect 24633 6409 24645 6412
rect 24587 6403 24645 6409
rect 25406 6400 25412 6412
rect 25464 6400 25470 6452
rect 26142 6400 26148 6452
rect 26200 6440 26206 6452
rect 26237 6443 26295 6449
rect 26237 6440 26249 6443
rect 26200 6412 26249 6440
rect 26200 6400 26206 6412
rect 26237 6409 26249 6412
rect 26283 6409 26295 6443
rect 26237 6403 26295 6409
rect 28813 6443 28871 6449
rect 28813 6409 28825 6443
rect 28859 6409 28871 6443
rect 29270 6440 29276 6452
rect 29231 6412 29276 6440
rect 28813 6403 28871 6409
rect 23753 6375 23811 6381
rect 23753 6341 23765 6375
rect 23799 6372 23811 6375
rect 23842 6372 23848 6384
rect 23799 6344 23848 6372
rect 23799 6341 23811 6344
rect 23753 6335 23811 6341
rect 23842 6332 23848 6344
rect 23900 6332 23906 6384
rect 24394 6332 24400 6384
rect 24452 6372 24458 6384
rect 24489 6375 24547 6381
rect 24489 6372 24501 6375
rect 24452 6344 24501 6372
rect 24452 6332 24458 6344
rect 24489 6341 24501 6344
rect 24535 6341 24547 6375
rect 26418 6372 26424 6384
rect 24489 6335 24547 6341
rect 24780 6344 26424 6372
rect 21177 6307 21235 6313
rect 21177 6304 21189 6307
rect 20732 6276 21189 6304
rect 21177 6273 21189 6276
rect 21223 6273 21235 6307
rect 21358 6304 21364 6316
rect 21319 6276 21364 6304
rect 21177 6267 21235 6273
rect 21358 6264 21364 6276
rect 21416 6264 21422 6316
rect 24670 6304 24676 6316
rect 24631 6276 24676 6304
rect 24670 6264 24676 6276
rect 24728 6264 24734 6316
rect 24780 6313 24808 6344
rect 26418 6332 26424 6344
rect 26476 6372 26482 6384
rect 26476 6344 28396 6372
rect 26476 6332 26482 6344
rect 24765 6307 24823 6313
rect 24765 6273 24777 6307
rect 24811 6273 24823 6307
rect 24765 6267 24823 6273
rect 26053 6307 26111 6313
rect 26053 6273 26065 6307
rect 26099 6273 26111 6307
rect 26053 6267 26111 6273
rect 23937 6239 23995 6245
rect 23937 6205 23949 6239
rect 23983 6205 23995 6239
rect 26068 6236 26096 6267
rect 26142 6264 26148 6316
rect 26200 6304 26206 6316
rect 26329 6307 26387 6313
rect 26329 6304 26341 6307
rect 26200 6276 26341 6304
rect 26200 6264 26206 6276
rect 26329 6273 26341 6276
rect 26375 6273 26387 6307
rect 26329 6267 26387 6273
rect 27700 6307 27758 6313
rect 27700 6273 27712 6307
rect 27746 6304 27758 6307
rect 28074 6304 28080 6316
rect 27746 6276 28080 6304
rect 27746 6273 27758 6276
rect 27700 6267 27758 6273
rect 28074 6264 28080 6276
rect 28132 6264 28138 6316
rect 28368 6304 28396 6344
rect 28442 6332 28448 6384
rect 28500 6372 28506 6384
rect 28828 6372 28856 6403
rect 29270 6400 29276 6412
rect 29328 6400 29334 6452
rect 30098 6400 30104 6452
rect 30156 6440 30162 6452
rect 30469 6443 30527 6449
rect 30469 6440 30481 6443
rect 30156 6412 30481 6440
rect 30156 6400 30162 6412
rect 30469 6409 30481 6412
rect 30515 6409 30527 6443
rect 30469 6403 30527 6409
rect 33965 6443 34023 6449
rect 33965 6409 33977 6443
rect 34011 6440 34023 6443
rect 35526 6440 35532 6452
rect 34011 6412 35532 6440
rect 34011 6409 34023 6412
rect 33965 6403 34023 6409
rect 35526 6400 35532 6412
rect 35584 6400 35590 6452
rect 29641 6375 29699 6381
rect 29641 6372 29653 6375
rect 28500 6344 29653 6372
rect 28500 6332 28506 6344
rect 29641 6341 29653 6344
rect 29687 6341 29699 6375
rect 29641 6335 29699 6341
rect 33597 6375 33655 6381
rect 33597 6341 33609 6375
rect 33643 6372 33655 6375
rect 33870 6372 33876 6384
rect 33643 6344 33876 6372
rect 33643 6341 33655 6344
rect 33597 6335 33655 6341
rect 33870 6332 33876 6344
rect 33928 6332 33934 6384
rect 34698 6332 34704 6384
rect 34756 6372 34762 6384
rect 34793 6375 34851 6381
rect 34793 6372 34805 6375
rect 34756 6344 34805 6372
rect 34756 6332 34762 6344
rect 34793 6341 34805 6344
rect 34839 6341 34851 6375
rect 34793 6335 34851 6341
rect 34882 6332 34888 6384
rect 34940 6372 34946 6384
rect 35342 6372 35348 6384
rect 34940 6344 35204 6372
rect 34940 6332 34946 6344
rect 29086 6304 29092 6316
rect 28368 6276 29092 6304
rect 29086 6264 29092 6276
rect 29144 6264 29150 6316
rect 30834 6304 30840 6316
rect 30795 6276 30840 6304
rect 30834 6264 30840 6276
rect 30892 6264 30898 6316
rect 33778 6304 33784 6316
rect 33739 6276 33784 6304
rect 33778 6264 33784 6276
rect 33836 6264 33842 6316
rect 35176 6313 35204 6344
rect 35268 6344 35348 6372
rect 35268 6313 35296 6344
rect 35342 6332 35348 6344
rect 35400 6332 35406 6384
rect 38102 6372 38108 6384
rect 38063 6344 38108 6372
rect 38102 6332 38108 6344
rect 38160 6332 38166 6384
rect 35069 6307 35127 6313
rect 35069 6273 35081 6307
rect 35115 6273 35127 6307
rect 35069 6267 35127 6273
rect 35161 6307 35219 6313
rect 35161 6273 35173 6307
rect 35207 6273 35219 6307
rect 35161 6267 35219 6273
rect 35253 6307 35311 6313
rect 35253 6273 35265 6307
rect 35299 6273 35311 6307
rect 35434 6304 35440 6316
rect 35395 6276 35440 6304
rect 35253 6267 35311 6273
rect 27430 6236 27436 6248
rect 26068 6208 26280 6236
rect 27391 6208 27436 6236
rect 23937 6199 23995 6205
rect 23952 6168 23980 6199
rect 26252 6180 26280 6208
rect 27430 6196 27436 6208
rect 27488 6196 27494 6248
rect 23952 6140 26188 6168
rect 15470 6060 15476 6112
rect 15528 6100 15534 6112
rect 15657 6103 15715 6109
rect 15657 6100 15669 6103
rect 15528 6072 15669 6100
rect 15528 6060 15534 6072
rect 15657 6069 15669 6072
rect 15703 6069 15715 6103
rect 20530 6100 20536 6112
rect 20491 6072 20536 6100
rect 15657 6063 15715 6069
rect 20530 6060 20536 6072
rect 20588 6060 20594 6112
rect 21174 6100 21180 6112
rect 21135 6072 21180 6100
rect 21174 6060 21180 6072
rect 21232 6060 21238 6112
rect 25869 6103 25927 6109
rect 25869 6069 25881 6103
rect 25915 6100 25927 6103
rect 26050 6100 26056 6112
rect 25915 6072 26056 6100
rect 25915 6069 25927 6072
rect 25869 6063 25927 6069
rect 26050 6060 26056 6072
rect 26108 6060 26114 6112
rect 26160 6100 26188 6140
rect 26234 6128 26240 6180
rect 26292 6128 26298 6180
rect 29104 6168 29132 6264
rect 29730 6236 29736 6248
rect 29691 6208 29736 6236
rect 29730 6196 29736 6208
rect 29788 6196 29794 6248
rect 29914 6236 29920 6248
rect 29875 6208 29920 6236
rect 29914 6196 29920 6208
rect 29972 6196 29978 6248
rect 30926 6236 30932 6248
rect 30887 6208 30932 6236
rect 30926 6196 30932 6208
rect 30984 6196 30990 6248
rect 31018 6196 31024 6248
rect 31076 6236 31082 6248
rect 35084 6236 35112 6267
rect 35434 6264 35440 6276
rect 35492 6264 35498 6316
rect 35618 6264 35624 6316
rect 35676 6304 35682 6316
rect 37829 6307 37887 6313
rect 37829 6304 37841 6307
rect 35676 6276 37841 6304
rect 35676 6264 35682 6276
rect 37829 6273 37841 6276
rect 37875 6273 37887 6307
rect 37829 6267 37887 6273
rect 38286 6236 38292 6248
rect 31076 6208 31169 6236
rect 35084 6208 38292 6236
rect 31076 6196 31082 6208
rect 38286 6196 38292 6208
rect 38344 6196 38350 6248
rect 31036 6168 31064 6196
rect 29104 6140 31064 6168
rect 27246 6100 27252 6112
rect 26160 6072 27252 6100
rect 27246 6060 27252 6072
rect 27304 6060 27310 6112
rect 35066 6060 35072 6112
rect 35124 6100 35130 6112
rect 36630 6100 36636 6112
rect 35124 6072 36636 6100
rect 35124 6060 35130 6072
rect 36630 6060 36636 6072
rect 36688 6060 36694 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 17129 5899 17187 5905
rect 17129 5865 17141 5899
rect 17175 5896 17187 5899
rect 17402 5896 17408 5908
rect 17175 5868 17408 5896
rect 17175 5865 17187 5868
rect 17129 5859 17187 5865
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 25958 5896 25964 5908
rect 25919 5868 25964 5896
rect 25958 5856 25964 5868
rect 26016 5856 26022 5908
rect 28074 5896 28080 5908
rect 28035 5868 28080 5896
rect 28074 5856 28080 5868
rect 28132 5856 28138 5908
rect 35253 5899 35311 5905
rect 35253 5865 35265 5899
rect 35299 5896 35311 5899
rect 35434 5896 35440 5908
rect 35299 5868 35440 5896
rect 35299 5865 35311 5868
rect 35253 5859 35311 5865
rect 35434 5856 35440 5868
rect 35492 5856 35498 5908
rect 38286 5896 38292 5908
rect 38247 5868 38292 5896
rect 38286 5856 38292 5868
rect 38344 5856 38350 5908
rect 22465 5831 22523 5837
rect 22465 5797 22477 5831
rect 22511 5828 22523 5831
rect 25869 5831 25927 5837
rect 22511 5800 25820 5828
rect 22511 5797 22523 5800
rect 22465 5791 22523 5797
rect 20901 5763 20959 5769
rect 20901 5729 20913 5763
rect 20947 5760 20959 5763
rect 22094 5760 22100 5772
rect 20947 5732 22100 5760
rect 20947 5729 20959 5732
rect 20901 5723 20959 5729
rect 22094 5720 22100 5732
rect 22152 5720 22158 5772
rect 23842 5720 23848 5772
rect 23900 5760 23906 5772
rect 24762 5760 24768 5772
rect 23900 5732 24768 5760
rect 23900 5720 23906 5732
rect 24762 5720 24768 5732
rect 24820 5760 24826 5772
rect 25041 5763 25099 5769
rect 25041 5760 25053 5763
rect 24820 5732 25053 5760
rect 24820 5720 24826 5732
rect 25041 5729 25053 5732
rect 25087 5729 25099 5763
rect 25041 5723 25099 5729
rect 25225 5763 25283 5769
rect 25225 5729 25237 5763
rect 25271 5760 25283 5763
rect 25314 5760 25320 5772
rect 25271 5732 25320 5760
rect 25271 5729 25283 5732
rect 25225 5723 25283 5729
rect 25314 5720 25320 5732
rect 25372 5720 25378 5772
rect 25792 5760 25820 5800
rect 25869 5797 25881 5831
rect 25915 5828 25927 5831
rect 26418 5828 26424 5840
rect 25915 5800 26424 5828
rect 25915 5797 25927 5800
rect 25869 5791 25927 5797
rect 26418 5788 26424 5800
rect 26476 5788 26482 5840
rect 27246 5788 27252 5840
rect 27304 5828 27310 5840
rect 27304 5800 28672 5828
rect 27304 5788 27310 5800
rect 26050 5760 26056 5772
rect 25792 5732 25912 5760
rect 26011 5732 26056 5760
rect 15470 5692 15476 5704
rect 15431 5664 15476 5692
rect 15470 5652 15476 5664
rect 15528 5652 15534 5704
rect 16022 5692 16028 5704
rect 15983 5664 16028 5692
rect 16022 5652 16028 5664
rect 16080 5652 16086 5704
rect 18230 5692 18236 5704
rect 18191 5664 18236 5692
rect 18230 5652 18236 5664
rect 18288 5652 18294 5704
rect 18417 5695 18475 5701
rect 18417 5661 18429 5695
rect 18463 5692 18475 5695
rect 18782 5692 18788 5704
rect 18463 5664 18788 5692
rect 18463 5661 18475 5664
rect 18417 5655 18475 5661
rect 18782 5652 18788 5664
rect 18840 5652 18846 5704
rect 21174 5692 21180 5704
rect 21135 5664 21180 5692
rect 21174 5652 21180 5664
rect 21232 5652 21238 5704
rect 25777 5695 25835 5701
rect 25777 5692 25789 5695
rect 24964 5664 25789 5692
rect 24964 5568 24992 5664
rect 25777 5661 25789 5664
rect 25823 5661 25835 5695
rect 25884 5692 25912 5732
rect 26050 5720 26056 5732
rect 26108 5720 26114 5772
rect 27982 5720 27988 5772
rect 28040 5760 28046 5772
rect 28350 5760 28356 5772
rect 28040 5732 28356 5760
rect 28040 5720 28046 5732
rect 28350 5720 28356 5732
rect 28408 5760 28414 5772
rect 28644 5769 28672 5800
rect 28537 5763 28595 5769
rect 28537 5760 28549 5763
rect 28408 5732 28549 5760
rect 28408 5720 28414 5732
rect 28537 5729 28549 5732
rect 28583 5729 28595 5763
rect 28537 5723 28595 5729
rect 28629 5763 28687 5769
rect 28629 5729 28641 5763
rect 28675 5729 28687 5763
rect 28629 5723 28687 5729
rect 33042 5720 33048 5772
rect 33100 5760 33106 5772
rect 34149 5763 34207 5769
rect 34149 5760 34161 5763
rect 33100 5732 34161 5760
rect 33100 5720 33106 5732
rect 34149 5729 34161 5732
rect 34195 5729 34207 5763
rect 34149 5723 34207 5729
rect 36722 5720 36728 5772
rect 36780 5760 36786 5772
rect 36909 5763 36967 5769
rect 36909 5760 36921 5763
rect 36780 5732 36921 5760
rect 36780 5720 36786 5732
rect 36909 5729 36921 5732
rect 36955 5729 36967 5763
rect 36909 5723 36967 5729
rect 28258 5692 28264 5704
rect 25884 5664 28264 5692
rect 25777 5655 25835 5661
rect 28258 5652 28264 5664
rect 28316 5652 28322 5704
rect 28442 5692 28448 5704
rect 28403 5664 28448 5692
rect 28442 5652 28448 5664
rect 28500 5652 28506 5704
rect 30469 5695 30527 5701
rect 30469 5661 30481 5695
rect 30515 5692 30527 5695
rect 31662 5692 31668 5704
rect 30515 5664 31668 5692
rect 30515 5661 30527 5664
rect 30469 5655 30527 5661
rect 31662 5652 31668 5664
rect 31720 5652 31726 5704
rect 33965 5695 34023 5701
rect 33965 5661 33977 5695
rect 34011 5692 34023 5695
rect 34011 5664 35112 5692
rect 34011 5661 34023 5664
rect 33965 5655 34023 5661
rect 30558 5584 30564 5636
rect 30616 5624 30622 5636
rect 30714 5627 30772 5633
rect 30714 5624 30726 5627
rect 30616 5596 30726 5624
rect 30616 5584 30622 5596
rect 30714 5593 30726 5596
rect 30760 5593 30772 5627
rect 30714 5587 30772 5593
rect 33870 5584 33876 5636
rect 33928 5624 33934 5636
rect 35084 5633 35112 5664
rect 34885 5627 34943 5633
rect 34885 5624 34897 5627
rect 33928 5596 34897 5624
rect 33928 5584 33934 5596
rect 34885 5593 34897 5596
rect 34931 5593 34943 5627
rect 34885 5587 34943 5593
rect 35069 5627 35127 5633
rect 35069 5593 35081 5627
rect 35115 5624 35127 5627
rect 35342 5624 35348 5636
rect 35115 5596 35348 5624
rect 35115 5593 35127 5596
rect 35069 5587 35127 5593
rect 35342 5584 35348 5596
rect 35400 5584 35406 5636
rect 37176 5627 37234 5633
rect 37176 5593 37188 5627
rect 37222 5624 37234 5627
rect 37458 5624 37464 5636
rect 37222 5596 37464 5624
rect 37222 5593 37234 5596
rect 37176 5587 37234 5593
rect 37458 5584 37464 5596
rect 37516 5584 37522 5636
rect 18322 5556 18328 5568
rect 18283 5528 18328 5556
rect 18322 5516 18328 5528
rect 18380 5516 18386 5568
rect 24578 5556 24584 5568
rect 24539 5528 24584 5556
rect 24578 5516 24584 5528
rect 24636 5516 24642 5568
rect 24946 5556 24952 5568
rect 24907 5528 24952 5556
rect 24946 5516 24952 5528
rect 25004 5516 25010 5568
rect 30834 5516 30840 5568
rect 30892 5556 30898 5568
rect 31849 5559 31907 5565
rect 31849 5556 31861 5559
rect 30892 5528 31861 5556
rect 30892 5516 30898 5528
rect 31849 5525 31861 5528
rect 31895 5525 31907 5559
rect 31849 5519 31907 5525
rect 33597 5559 33655 5565
rect 33597 5525 33609 5559
rect 33643 5556 33655 5559
rect 33686 5556 33692 5568
rect 33643 5528 33692 5556
rect 33643 5525 33655 5528
rect 33597 5519 33655 5525
rect 33686 5516 33692 5528
rect 33744 5516 33750 5568
rect 34057 5559 34115 5565
rect 34057 5525 34069 5559
rect 34103 5556 34115 5559
rect 35710 5556 35716 5568
rect 34103 5528 35716 5556
rect 34103 5525 34115 5528
rect 34057 5519 34115 5525
rect 35710 5516 35716 5528
rect 35768 5556 35774 5568
rect 37918 5556 37924 5568
rect 35768 5528 37924 5556
rect 35768 5516 35774 5528
rect 37918 5516 37924 5528
rect 37976 5516 37982 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 21269 5355 21327 5361
rect 21269 5321 21281 5355
rect 21315 5352 21327 5355
rect 22830 5352 22836 5364
rect 21315 5324 22836 5352
rect 21315 5321 21327 5324
rect 21269 5315 21327 5321
rect 22830 5312 22836 5324
rect 22888 5312 22894 5364
rect 23474 5312 23480 5364
rect 23532 5352 23538 5364
rect 23569 5355 23627 5361
rect 23569 5352 23581 5355
rect 23532 5324 23581 5352
rect 23532 5312 23538 5324
rect 23569 5321 23581 5324
rect 23615 5352 23627 5355
rect 24670 5352 24676 5364
rect 23615 5324 24676 5352
rect 23615 5321 23627 5324
rect 23569 5315 23627 5321
rect 24670 5312 24676 5324
rect 24728 5312 24734 5364
rect 24946 5312 24952 5364
rect 25004 5352 25010 5364
rect 25409 5355 25467 5361
rect 25409 5352 25421 5355
rect 25004 5324 25421 5352
rect 25004 5312 25010 5324
rect 25409 5321 25421 5324
rect 25455 5321 25467 5355
rect 25409 5315 25467 5321
rect 30469 5355 30527 5361
rect 30469 5321 30481 5355
rect 30515 5352 30527 5355
rect 30558 5352 30564 5364
rect 30515 5324 30564 5352
rect 30515 5321 30527 5324
rect 30469 5315 30527 5321
rect 30558 5312 30564 5324
rect 30616 5312 30622 5364
rect 30834 5352 30840 5364
rect 30795 5324 30840 5352
rect 30834 5312 30840 5324
rect 30892 5312 30898 5364
rect 33689 5355 33747 5361
rect 33689 5321 33701 5355
rect 33735 5352 33747 5355
rect 33778 5352 33784 5364
rect 33735 5324 33784 5352
rect 33735 5321 33747 5324
rect 33689 5315 33747 5321
rect 33778 5312 33784 5324
rect 33836 5312 33842 5364
rect 36630 5352 36636 5364
rect 36591 5324 36636 5352
rect 36630 5312 36636 5324
rect 36688 5312 36694 5364
rect 37458 5352 37464 5364
rect 37419 5324 37464 5352
rect 37458 5312 37464 5324
rect 37516 5312 37522 5364
rect 37829 5355 37887 5361
rect 37829 5321 37841 5355
rect 37875 5352 37887 5355
rect 38286 5352 38292 5364
rect 37875 5324 38292 5352
rect 37875 5321 37887 5324
rect 37829 5315 37887 5321
rect 38286 5312 38292 5324
rect 38344 5312 38350 5364
rect 18049 5287 18107 5293
rect 18049 5253 18061 5287
rect 18095 5284 18107 5287
rect 18322 5284 18328 5296
rect 18095 5256 18328 5284
rect 18095 5253 18107 5256
rect 18049 5247 18107 5253
rect 18322 5244 18328 5256
rect 18380 5244 18386 5296
rect 23198 5284 23204 5296
rect 22204 5256 23204 5284
rect 19705 5219 19763 5225
rect 19705 5185 19717 5219
rect 19751 5216 19763 5219
rect 22094 5216 22100 5228
rect 19751 5188 22100 5216
rect 19751 5185 19763 5188
rect 19705 5179 19763 5185
rect 22094 5176 22100 5188
rect 22152 5216 22158 5228
rect 22204 5225 22232 5256
rect 23198 5244 23204 5256
rect 23256 5244 23262 5296
rect 24296 5287 24354 5293
rect 24296 5253 24308 5287
rect 24342 5284 24354 5287
rect 24578 5284 24584 5296
rect 24342 5256 24584 5284
rect 24342 5253 24354 5256
rect 24296 5247 24354 5253
rect 24578 5244 24584 5256
rect 24636 5244 24642 5296
rect 24762 5244 24768 5296
rect 24820 5284 24826 5296
rect 26329 5287 26387 5293
rect 26329 5284 26341 5287
rect 24820 5256 26341 5284
rect 24820 5244 24826 5256
rect 26329 5253 26341 5256
rect 26375 5253 26387 5287
rect 26329 5247 26387 5253
rect 28350 5244 28356 5296
rect 28408 5284 28414 5296
rect 30929 5287 30987 5293
rect 30929 5284 30941 5287
rect 28408 5256 30941 5284
rect 28408 5244 28414 5256
rect 30929 5253 30941 5256
rect 30975 5253 30987 5287
rect 37918 5284 37924 5296
rect 30929 5247 30987 5253
rect 32324 5256 33640 5284
rect 37879 5256 37924 5284
rect 22189 5219 22247 5225
rect 22189 5216 22201 5219
rect 22152 5188 22201 5216
rect 22152 5176 22158 5188
rect 22189 5185 22201 5188
rect 22235 5185 22247 5219
rect 22189 5179 22247 5185
rect 22456 5219 22514 5225
rect 22456 5185 22468 5219
rect 22502 5216 22514 5219
rect 23014 5216 23020 5228
rect 22502 5188 23020 5216
rect 22502 5185 22514 5188
rect 22456 5179 22514 5185
rect 23014 5176 23020 5188
rect 23072 5176 23078 5228
rect 26234 5216 26240 5228
rect 26147 5188 26240 5216
rect 26234 5176 26240 5188
rect 26292 5216 26298 5228
rect 26970 5216 26976 5228
rect 26292 5188 26976 5216
rect 26292 5176 26298 5188
rect 26970 5176 26976 5188
rect 27028 5176 27034 5228
rect 31754 5176 31760 5228
rect 31812 5216 31818 5228
rect 32324 5225 32352 5256
rect 32582 5225 32588 5228
rect 32309 5219 32367 5225
rect 32309 5216 32321 5219
rect 31812 5188 32321 5216
rect 31812 5176 31818 5188
rect 32309 5185 32321 5188
rect 32355 5185 32367 5219
rect 32309 5179 32367 5185
rect 32576 5179 32588 5225
rect 32640 5216 32646 5228
rect 32640 5188 32676 5216
rect 32582 5176 32588 5179
rect 32640 5176 32646 5188
rect 33612 5160 33640 5256
rect 37918 5244 37924 5256
rect 37976 5244 37982 5296
rect 35526 5225 35532 5228
rect 35520 5179 35532 5225
rect 35584 5216 35590 5228
rect 35584 5188 35620 5216
rect 35526 5176 35532 5179
rect 35584 5176 35590 5188
rect 18966 5108 18972 5160
rect 19024 5148 19030 5160
rect 19981 5151 20039 5157
rect 19981 5148 19993 5151
rect 19024 5120 19993 5148
rect 19024 5108 19030 5120
rect 19981 5117 19993 5120
rect 20027 5117 20039 5151
rect 19981 5111 20039 5117
rect 23198 5108 23204 5160
rect 23256 5148 23262 5160
rect 24026 5148 24032 5160
rect 23256 5120 24032 5148
rect 23256 5108 23262 5120
rect 24026 5108 24032 5120
rect 24084 5108 24090 5160
rect 26510 5148 26516 5160
rect 26471 5120 26516 5148
rect 26510 5108 26516 5120
rect 26568 5108 26574 5160
rect 30742 5108 30748 5160
rect 30800 5148 30806 5160
rect 31021 5151 31079 5157
rect 31021 5148 31033 5151
rect 30800 5120 31033 5148
rect 30800 5108 30806 5120
rect 31021 5117 31033 5120
rect 31067 5148 31079 5151
rect 32214 5148 32220 5160
rect 31067 5120 32220 5148
rect 31067 5117 31079 5120
rect 31021 5111 31079 5117
rect 32214 5108 32220 5120
rect 32272 5108 32278 5160
rect 33594 5108 33600 5160
rect 33652 5148 33658 5160
rect 35253 5151 35311 5157
rect 35253 5148 35265 5151
rect 33652 5120 35265 5148
rect 33652 5108 33658 5120
rect 35253 5117 35265 5120
rect 35299 5117 35311 5151
rect 38010 5148 38016 5160
rect 37971 5120 38016 5148
rect 35253 5111 35311 5117
rect 38010 5108 38016 5120
rect 38068 5108 38074 5160
rect 17954 5040 17960 5092
rect 18012 5080 18018 5092
rect 18325 5083 18383 5089
rect 18325 5080 18337 5083
rect 18012 5052 18337 5080
rect 18012 5040 18018 5052
rect 18325 5049 18337 5052
rect 18371 5049 18383 5083
rect 18325 5043 18383 5049
rect 18506 5012 18512 5024
rect 18467 4984 18512 5012
rect 18506 4972 18512 4984
rect 18564 4972 18570 5024
rect 25866 5012 25872 5024
rect 25827 4984 25872 5012
rect 25866 4972 25872 4984
rect 25924 4972 25930 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 23014 4808 23020 4820
rect 22975 4780 23020 4808
rect 23014 4768 23020 4780
rect 23072 4768 23078 4820
rect 26970 4808 26976 4820
rect 26931 4780 26976 4808
rect 26970 4768 26976 4780
rect 27028 4768 27034 4820
rect 28813 4811 28871 4817
rect 28813 4777 28825 4811
rect 28859 4808 28871 4811
rect 28994 4808 29000 4820
rect 28859 4780 29000 4808
rect 28859 4777 28871 4780
rect 28813 4771 28871 4777
rect 28994 4768 29000 4780
rect 29052 4808 29058 4820
rect 29730 4808 29736 4820
rect 29052 4780 29736 4808
rect 29052 4768 29058 4780
rect 29730 4768 29736 4780
rect 29788 4768 29794 4820
rect 30926 4768 30932 4820
rect 30984 4808 30990 4820
rect 31113 4811 31171 4817
rect 31113 4808 31125 4811
rect 30984 4780 31125 4808
rect 30984 4768 30990 4780
rect 31113 4777 31125 4780
rect 31159 4777 31171 4811
rect 32582 4808 32588 4820
rect 32543 4780 32588 4808
rect 31113 4771 31171 4777
rect 32582 4768 32588 4780
rect 32640 4768 32646 4820
rect 35526 4768 35532 4820
rect 35584 4808 35590 4820
rect 35621 4811 35679 4817
rect 35621 4808 35633 4811
rect 35584 4780 35633 4808
rect 35584 4768 35590 4780
rect 35621 4777 35633 4780
rect 35667 4777 35679 4811
rect 35621 4771 35679 4777
rect 17497 4743 17555 4749
rect 17497 4709 17509 4743
rect 17543 4740 17555 4743
rect 23658 4740 23664 4752
rect 17543 4712 23664 4740
rect 17543 4709 17555 4712
rect 17497 4703 17555 4709
rect 23658 4700 23664 4712
rect 23716 4700 23722 4752
rect 32214 4700 32220 4752
rect 32272 4740 32278 4752
rect 38010 4740 38016 4752
rect 32272 4712 38016 4740
rect 32272 4700 32278 4712
rect 16209 4675 16267 4681
rect 16209 4641 16221 4675
rect 16255 4672 16267 4675
rect 17402 4672 17408 4684
rect 16255 4644 17408 4672
rect 16255 4641 16267 4644
rect 16209 4635 16267 4641
rect 17402 4632 17408 4644
rect 17460 4632 17466 4684
rect 23566 4672 23572 4684
rect 23527 4644 23572 4672
rect 23566 4632 23572 4644
rect 23624 4632 23630 4684
rect 33042 4672 33048 4684
rect 31726 4644 33048 4672
rect 15930 4604 15936 4616
rect 15891 4576 15936 4604
rect 15930 4564 15936 4576
rect 15988 4564 15994 4616
rect 23385 4607 23443 4613
rect 23385 4573 23397 4607
rect 23431 4604 23443 4607
rect 23474 4604 23480 4616
rect 23431 4576 23480 4604
rect 23431 4573 23443 4576
rect 23385 4567 23443 4573
rect 23474 4564 23480 4576
rect 23532 4564 23538 4616
rect 24026 4564 24032 4616
rect 24084 4604 24090 4616
rect 25593 4607 25651 4613
rect 25593 4604 25605 4607
rect 24084 4576 25605 4604
rect 24084 4564 24090 4576
rect 25593 4573 25605 4576
rect 25639 4604 25651 4607
rect 27430 4604 27436 4616
rect 25639 4576 27436 4604
rect 25639 4573 25651 4576
rect 25593 4567 25651 4573
rect 27430 4564 27436 4576
rect 27488 4604 27494 4616
rect 29733 4607 29791 4613
rect 29733 4604 29745 4607
rect 27488 4576 29745 4604
rect 27488 4564 27494 4576
rect 29733 4573 29745 4576
rect 29779 4573 29791 4607
rect 29733 4567 29791 4573
rect 30282 4564 30288 4616
rect 30340 4604 30346 4616
rect 31726 4604 31754 4644
rect 33042 4632 33048 4644
rect 33100 4672 33106 4684
rect 33137 4675 33195 4681
rect 33137 4672 33149 4675
rect 33100 4644 33149 4672
rect 33100 4632 33106 4644
rect 33137 4641 33149 4644
rect 33183 4641 33195 4675
rect 33137 4635 33195 4641
rect 35894 4632 35900 4684
rect 35952 4672 35958 4684
rect 36188 4681 36216 4712
rect 38010 4700 38016 4712
rect 38068 4700 38074 4752
rect 36081 4675 36139 4681
rect 36081 4672 36093 4675
rect 35952 4644 36093 4672
rect 35952 4632 35958 4644
rect 36081 4641 36093 4644
rect 36127 4641 36139 4675
rect 36081 4635 36139 4641
rect 36173 4675 36231 4681
rect 36173 4641 36185 4675
rect 36219 4641 36231 4675
rect 38102 4672 38108 4684
rect 38063 4644 38108 4672
rect 36173 4635 36231 4641
rect 38102 4632 38108 4644
rect 38160 4632 38166 4684
rect 30340 4576 31754 4604
rect 32953 4607 33011 4613
rect 30340 4564 30346 4576
rect 32953 4573 32965 4607
rect 32999 4604 33011 4607
rect 33778 4604 33784 4616
rect 32999 4576 33784 4604
rect 32999 4573 33011 4576
rect 32953 4567 33011 4573
rect 33778 4564 33784 4576
rect 33836 4564 33842 4616
rect 35989 4607 36047 4613
rect 35989 4573 36001 4607
rect 36035 4604 36047 4607
rect 36630 4604 36636 4616
rect 36035 4576 36636 4604
rect 36035 4573 36047 4576
rect 35989 4567 36047 4573
rect 36630 4564 36636 4576
rect 36688 4564 36694 4616
rect 37829 4607 37887 4613
rect 37829 4573 37841 4607
rect 37875 4573 37887 4607
rect 37829 4567 37887 4573
rect 25866 4545 25872 4548
rect 25860 4536 25872 4545
rect 25827 4508 25872 4536
rect 25860 4499 25872 4508
rect 25866 4496 25872 4499
rect 25924 4496 25930 4548
rect 27700 4539 27758 4545
rect 27700 4505 27712 4539
rect 27746 4536 27758 4539
rect 27890 4536 27896 4548
rect 27746 4508 27896 4536
rect 27746 4505 27758 4508
rect 27700 4499 27758 4505
rect 27890 4496 27896 4508
rect 27948 4496 27954 4548
rect 30006 4545 30012 4548
rect 30000 4499 30012 4545
rect 30064 4536 30070 4548
rect 37844 4536 37872 4567
rect 30064 4508 30100 4536
rect 31726 4508 37872 4536
rect 30006 4496 30012 4499
rect 30064 4496 30070 4508
rect 23477 4471 23535 4477
rect 23477 4437 23489 4471
rect 23523 4468 23535 4471
rect 23842 4468 23848 4480
rect 23523 4440 23848 4468
rect 23523 4437 23535 4440
rect 23477 4431 23535 4437
rect 23842 4428 23848 4440
rect 23900 4428 23906 4480
rect 28166 4428 28172 4480
rect 28224 4468 28230 4480
rect 31726 4468 31754 4508
rect 28224 4440 31754 4468
rect 33045 4471 33103 4477
rect 28224 4428 28230 4440
rect 33045 4437 33057 4471
rect 33091 4468 33103 4471
rect 35894 4468 35900 4480
rect 33091 4440 35900 4468
rect 33091 4437 33103 4440
rect 33045 4431 33103 4437
rect 35894 4428 35900 4440
rect 35952 4428 35958 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 27890 4264 27896 4276
rect 27851 4236 27896 4264
rect 27890 4224 27896 4236
rect 27948 4224 27954 4276
rect 28261 4267 28319 4273
rect 28261 4233 28273 4267
rect 28307 4264 28319 4267
rect 28994 4264 29000 4276
rect 28307 4236 29000 4264
rect 28307 4233 28319 4236
rect 28261 4227 28319 4233
rect 28994 4224 29000 4236
rect 29052 4224 29058 4276
rect 29917 4267 29975 4273
rect 29917 4233 29929 4267
rect 29963 4264 29975 4267
rect 30006 4264 30012 4276
rect 29963 4236 30012 4264
rect 29963 4233 29975 4236
rect 29917 4227 29975 4233
rect 30006 4224 30012 4236
rect 30064 4224 30070 4276
rect 30285 4267 30343 4273
rect 30285 4233 30297 4267
rect 30331 4264 30343 4267
rect 30926 4264 30932 4276
rect 30331 4236 30932 4264
rect 30331 4233 30343 4236
rect 30285 4227 30343 4233
rect 30926 4224 30932 4236
rect 30984 4224 30990 4276
rect 30377 4199 30435 4205
rect 30377 4196 30389 4199
rect 28368 4168 30389 4196
rect 28368 4140 28396 4168
rect 30377 4165 30389 4168
rect 30423 4165 30435 4199
rect 30377 4159 30435 4165
rect 30466 4156 30472 4208
rect 30524 4156 30530 4208
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 18141 4131 18199 4137
rect 18141 4128 18153 4131
rect 15988 4100 18153 4128
rect 15988 4088 15994 4100
rect 18141 4097 18153 4100
rect 18187 4097 18199 4131
rect 18141 4091 18199 4097
rect 18417 4131 18475 4137
rect 18417 4097 18429 4131
rect 18463 4128 18475 4131
rect 18506 4128 18512 4140
rect 18463 4100 18512 4128
rect 18463 4097 18475 4100
rect 18417 4091 18475 4097
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 28350 4128 28356 4140
rect 28311 4100 28356 4128
rect 28350 4088 28356 4100
rect 28408 4088 28414 4140
rect 30484 4128 30512 4156
rect 33594 4128 33600 4140
rect 28460 4100 30512 4128
rect 33555 4100 33600 4128
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 19521 4063 19579 4069
rect 19521 4060 19533 4063
rect 19484 4032 19533 4060
rect 19484 4020 19490 4032
rect 19521 4029 19533 4032
rect 19567 4029 19579 4063
rect 19521 4023 19579 4029
rect 23566 4020 23572 4072
rect 23624 4060 23630 4072
rect 28460 4069 28488 4100
rect 33594 4088 33600 4100
rect 33652 4088 33658 4140
rect 33686 4088 33692 4140
rect 33744 4128 33750 4140
rect 33853 4131 33911 4137
rect 33853 4128 33865 4131
rect 33744 4100 33865 4128
rect 33744 4088 33750 4100
rect 33853 4097 33865 4100
rect 33899 4097 33911 4131
rect 33853 4091 33911 4097
rect 37829 4131 37887 4137
rect 37829 4097 37841 4131
rect 37875 4097 37887 4131
rect 38102 4128 38108 4140
rect 38063 4100 38108 4128
rect 37829 4091 37887 4097
rect 28445 4063 28503 4069
rect 28445 4060 28457 4063
rect 23624 4032 28457 4060
rect 23624 4020 23630 4032
rect 28445 4029 28457 4032
rect 28491 4029 28503 4063
rect 28445 4023 28503 4029
rect 29546 4020 29552 4072
rect 29604 4060 29610 4072
rect 30282 4060 30288 4072
rect 29604 4032 30288 4060
rect 29604 4020 29610 4032
rect 30282 4020 30288 4032
rect 30340 4060 30346 4072
rect 30469 4063 30527 4069
rect 30469 4060 30481 4063
rect 30340 4032 30481 4060
rect 30340 4020 30346 4032
rect 30469 4029 30481 4032
rect 30515 4029 30527 4063
rect 30469 4023 30527 4029
rect 37844 3992 37872 4091
rect 38102 4088 38108 4100
rect 38160 4088 38166 4140
rect 34808 3964 37872 3992
rect 29362 3884 29368 3936
rect 29420 3924 29426 3936
rect 34808 3924 34836 3964
rect 29420 3896 34836 3924
rect 34977 3927 35035 3933
rect 29420 3884 29426 3896
rect 34977 3893 34989 3927
rect 35023 3924 35035 3927
rect 35342 3924 35348 3936
rect 35023 3896 35348 3924
rect 35023 3893 35035 3896
rect 34977 3887 35035 3893
rect 35342 3884 35348 3896
rect 35400 3884 35406 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 27706 3000 27712 3052
rect 27764 3040 27770 3052
rect 37829 3043 37887 3049
rect 37829 3040 37841 3043
rect 27764 3012 37841 3040
rect 27764 3000 27770 3012
rect 37829 3009 37841 3012
rect 37875 3009 37887 3043
rect 37829 3003 37887 3009
rect 38102 2972 38108 2984
rect 38063 2944 38108 2972
rect 38102 2932 38108 2944
rect 38160 2932 38166 2984
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 27338 2388 27344 2440
rect 27396 2428 27402 2440
rect 37829 2431 37887 2437
rect 37829 2428 37841 2431
rect 27396 2400 37841 2428
rect 27396 2388 27402 2400
rect 37829 2397 37841 2400
rect 37875 2397 37887 2431
rect 37829 2391 37887 2397
rect 38102 2360 38108 2372
rect 38063 2332 38108 2360
rect 38102 2320 38108 2332
rect 38160 2320 38166 2372
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 9404 37272 9456 37324
rect 12164 37315 12216 37324
rect 12164 37281 12173 37315
rect 12173 37281 12207 37315
rect 12207 37281 12216 37315
rect 12164 37272 12216 37281
rect 26516 37315 26568 37324
rect 26516 37281 26525 37315
rect 26525 37281 26559 37315
rect 26559 37281 26568 37315
rect 26516 37272 26568 37281
rect 28080 37272 28132 37324
rect 30472 37272 30524 37324
rect 32680 37272 32732 37324
rect 1768 37204 1820 37256
rect 5080 37247 5132 37256
rect 5080 37213 5089 37247
rect 5089 37213 5123 37247
rect 5123 37213 5132 37247
rect 5080 37204 5132 37213
rect 8392 37204 8444 37256
rect 11704 37204 11756 37256
rect 15200 37247 15252 37256
rect 15200 37213 15209 37247
rect 15209 37213 15243 37247
rect 15243 37213 15252 37247
rect 15200 37204 15252 37213
rect 5540 37136 5592 37188
rect 5724 37136 5776 37188
rect 9312 37136 9364 37188
rect 9496 37179 9548 37188
rect 9496 37145 9505 37179
rect 9505 37145 9539 37179
rect 9539 37145 9548 37179
rect 9496 37136 9548 37145
rect 16028 37136 16080 37188
rect 18328 37204 18380 37256
rect 22100 37247 22152 37256
rect 22100 37213 22109 37247
rect 22109 37213 22143 37247
rect 22143 37213 22152 37247
rect 22100 37204 22152 37213
rect 24952 37204 25004 37256
rect 26240 37204 26292 37256
rect 27436 37204 27488 37256
rect 28264 37204 28316 37256
rect 31760 37204 31812 37256
rect 33784 37247 33836 37256
rect 33784 37213 33793 37247
rect 33793 37213 33827 37247
rect 33827 37213 33836 37247
rect 33784 37204 33836 37213
rect 36452 37247 36504 37256
rect 36452 37213 36461 37247
rect 36461 37213 36495 37247
rect 36495 37213 36504 37247
rect 36452 37204 36504 37213
rect 38108 37204 38160 37256
rect 18604 37179 18656 37188
rect 18604 37145 18613 37179
rect 18613 37145 18647 37179
rect 18647 37145 18656 37179
rect 18604 37136 18656 37145
rect 9128 37111 9180 37120
rect 9128 37077 9137 37111
rect 9137 37077 9171 37111
rect 9171 37077 9180 37111
rect 9128 37068 9180 37077
rect 9588 37111 9640 37120
rect 9588 37077 9597 37111
rect 9597 37077 9631 37111
rect 9631 37077 9640 37111
rect 9588 37068 9640 37077
rect 12992 37068 13044 37120
rect 24308 37136 24360 37188
rect 36728 37179 36780 37188
rect 22468 37068 22520 37120
rect 36728 37145 36737 37179
rect 36737 37145 36771 37179
rect 36771 37145 36780 37179
rect 36728 37136 36780 37145
rect 38016 37179 38068 37188
rect 38016 37145 38025 37179
rect 38025 37145 38059 37179
rect 38059 37145 38068 37179
rect 38016 37136 38068 37145
rect 28448 37068 28500 37120
rect 31024 37068 31076 37120
rect 33968 37111 34020 37120
rect 33968 37077 33977 37111
rect 33977 37077 34011 37111
rect 34011 37077 34020 37111
rect 33968 37068 34020 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 9588 36864 9640 36916
rect 9128 36796 9180 36848
rect 4528 36728 4580 36780
rect 5540 36728 5592 36780
rect 11520 36728 11572 36780
rect 12624 36728 12676 36780
rect 13360 36728 13412 36780
rect 15292 36796 15344 36848
rect 15844 36796 15896 36848
rect 16488 36728 16540 36780
rect 19524 36728 19576 36780
rect 19984 36728 20036 36780
rect 5632 36592 5684 36644
rect 7656 36660 7708 36712
rect 7932 36703 7984 36712
rect 7932 36669 7941 36703
rect 7941 36669 7975 36703
rect 7975 36669 7984 36703
rect 7932 36660 7984 36669
rect 14556 36703 14608 36712
rect 14556 36669 14565 36703
rect 14565 36669 14599 36703
rect 14599 36669 14608 36703
rect 14556 36660 14608 36669
rect 18052 36703 18104 36712
rect 18052 36669 18061 36703
rect 18061 36669 18095 36703
rect 18095 36669 18104 36703
rect 18052 36660 18104 36669
rect 20812 36660 20864 36712
rect 17684 36592 17736 36644
rect 20076 36592 20128 36644
rect 13084 36524 13136 36576
rect 16948 36567 17000 36576
rect 16948 36533 16957 36567
rect 16957 36533 16991 36567
rect 16991 36533 17000 36567
rect 16948 36524 17000 36533
rect 19892 36524 19944 36576
rect 22100 36728 22152 36780
rect 28356 36864 28408 36916
rect 38016 36864 38068 36916
rect 26424 36728 26476 36780
rect 27620 36796 27672 36848
rect 23020 36660 23072 36712
rect 24308 36660 24360 36712
rect 27068 36660 27120 36712
rect 23388 36567 23440 36576
rect 23388 36533 23397 36567
rect 23397 36533 23431 36567
rect 23431 36533 23440 36567
rect 23388 36524 23440 36533
rect 25688 36567 25740 36576
rect 25688 36533 25697 36567
rect 25697 36533 25731 36567
rect 25731 36533 25740 36567
rect 25688 36524 25740 36533
rect 28172 36728 28224 36780
rect 28632 36728 28684 36780
rect 30472 36728 30524 36780
rect 32772 36796 32824 36848
rect 33968 36796 34020 36848
rect 36820 36796 36872 36848
rect 32404 36728 32456 36780
rect 35992 36728 36044 36780
rect 37740 36728 37792 36780
rect 34244 36703 34296 36712
rect 34244 36669 34253 36703
rect 34253 36669 34287 36703
rect 34287 36669 34296 36703
rect 34244 36660 34296 36669
rect 38108 36703 38160 36712
rect 38108 36669 38117 36703
rect 38117 36669 38151 36703
rect 38151 36669 38160 36703
rect 38108 36660 38160 36669
rect 28264 36524 28316 36576
rect 29276 36524 29328 36576
rect 30104 36524 30156 36576
rect 33692 36567 33744 36576
rect 33692 36533 33701 36567
rect 33701 36533 33735 36567
rect 33735 36533 33744 36567
rect 33692 36524 33744 36533
rect 35624 36567 35676 36576
rect 35624 36533 35633 36567
rect 35633 36533 35667 36567
rect 35667 36533 35676 36567
rect 35624 36524 35676 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 12624 36363 12676 36372
rect 12624 36329 12633 36363
rect 12633 36329 12667 36363
rect 12667 36329 12676 36363
rect 12624 36320 12676 36329
rect 15292 36363 15344 36372
rect 15292 36329 15301 36363
rect 15301 36329 15335 36363
rect 15335 36329 15344 36363
rect 15292 36320 15344 36329
rect 19524 36363 19576 36372
rect 8576 36252 8628 36304
rect 9312 36252 9364 36304
rect 5632 36227 5684 36236
rect 5632 36193 5641 36227
rect 5641 36193 5675 36227
rect 5675 36193 5684 36227
rect 5632 36184 5684 36193
rect 5908 36184 5960 36236
rect 9496 36184 9548 36236
rect 11520 36252 11572 36304
rect 14004 36252 14056 36304
rect 13084 36227 13136 36236
rect 4620 36116 4672 36168
rect 7932 36116 7984 36168
rect 9680 36116 9732 36168
rect 13084 36193 13093 36227
rect 13093 36193 13127 36227
rect 13127 36193 13136 36227
rect 13084 36184 13136 36193
rect 13268 36227 13320 36236
rect 13268 36193 13277 36227
rect 13277 36193 13311 36227
rect 13311 36193 13320 36227
rect 13268 36184 13320 36193
rect 13544 36184 13596 36236
rect 19524 36329 19533 36363
rect 19533 36329 19567 36363
rect 19567 36329 19576 36363
rect 19524 36320 19576 36329
rect 27436 36363 27488 36372
rect 27436 36329 27445 36363
rect 27445 36329 27479 36363
rect 27479 36329 27488 36363
rect 27436 36320 27488 36329
rect 28172 36363 28224 36372
rect 28172 36329 28181 36363
rect 28181 36329 28215 36363
rect 28215 36329 28224 36363
rect 28172 36320 28224 36329
rect 30104 36363 30156 36372
rect 30104 36329 30113 36363
rect 30113 36329 30147 36363
rect 30147 36329 30156 36363
rect 30104 36320 30156 36329
rect 32404 36320 32456 36372
rect 32680 36363 32732 36372
rect 32680 36329 32689 36363
rect 32689 36329 32723 36363
rect 32723 36329 32732 36363
rect 32680 36320 32732 36329
rect 33784 36320 33836 36372
rect 15844 36227 15896 36236
rect 15844 36193 15853 36227
rect 15853 36193 15887 36227
rect 15887 36193 15896 36227
rect 15844 36184 15896 36193
rect 5540 36091 5592 36100
rect 5540 36057 5549 36091
rect 5549 36057 5583 36091
rect 5583 36057 5592 36091
rect 5540 36048 5592 36057
rect 7104 36048 7156 36100
rect 7840 36048 7892 36100
rect 11704 36048 11756 36100
rect 5264 35980 5316 36032
rect 7748 36023 7800 36032
rect 7748 35989 7757 36023
rect 7757 35989 7791 36023
rect 7791 35989 7800 36023
rect 7748 35980 7800 35989
rect 9588 35980 9640 36032
rect 11888 36023 11940 36032
rect 11888 35989 11897 36023
rect 11897 35989 11931 36023
rect 11931 35989 11940 36023
rect 11888 35980 11940 35989
rect 12716 36116 12768 36168
rect 12992 36159 13044 36168
rect 12992 36125 13001 36159
rect 13001 36125 13035 36159
rect 13035 36125 13044 36159
rect 12992 36116 13044 36125
rect 15200 36159 15252 36168
rect 15200 36125 15209 36159
rect 15209 36125 15243 36159
rect 15243 36125 15252 36159
rect 16488 36184 16540 36236
rect 16212 36159 16264 36168
rect 15200 36116 15252 36125
rect 16212 36125 16221 36159
rect 16221 36125 16255 36159
rect 16255 36125 16264 36159
rect 16212 36116 16264 36125
rect 18420 36159 18472 36168
rect 18420 36125 18429 36159
rect 18429 36125 18463 36159
rect 18463 36125 18472 36159
rect 18420 36116 18472 36125
rect 20628 36184 20680 36236
rect 24860 36252 24912 36304
rect 27068 36252 27120 36304
rect 32312 36252 32364 36304
rect 24952 36184 25004 36236
rect 27620 36184 27672 36236
rect 19892 36116 19944 36168
rect 20444 36116 20496 36168
rect 22928 36116 22980 36168
rect 23388 36116 23440 36168
rect 24676 36159 24728 36168
rect 24676 36125 24685 36159
rect 24685 36125 24719 36159
rect 24719 36125 24728 36159
rect 24676 36116 24728 36125
rect 26332 36159 26384 36168
rect 16948 36048 17000 36100
rect 18236 36048 18288 36100
rect 20812 36048 20864 36100
rect 20996 36048 21048 36100
rect 23756 36091 23808 36100
rect 23756 36057 23765 36091
rect 23765 36057 23799 36091
rect 23799 36057 23808 36091
rect 23756 36048 23808 36057
rect 23848 36048 23900 36100
rect 26332 36125 26341 36159
rect 26341 36125 26375 36159
rect 26375 36125 26384 36159
rect 26332 36116 26384 36125
rect 28356 36159 28408 36168
rect 28356 36125 28365 36159
rect 28365 36125 28399 36159
rect 28399 36125 28408 36159
rect 28356 36116 28408 36125
rect 30472 36184 30524 36236
rect 31208 36227 31260 36236
rect 31208 36193 31217 36227
rect 31217 36193 31251 36227
rect 31251 36193 31260 36227
rect 31208 36184 31260 36193
rect 27528 36048 27580 36100
rect 30012 36159 30064 36168
rect 30012 36125 30021 36159
rect 30021 36125 30055 36159
rect 30055 36125 30064 36159
rect 30012 36116 30064 36125
rect 34244 36184 34296 36236
rect 32588 36159 32640 36168
rect 32588 36125 32597 36159
rect 32597 36125 32631 36159
rect 32631 36125 32640 36159
rect 32588 36116 32640 36125
rect 33784 36116 33836 36168
rect 36268 36116 36320 36168
rect 29276 36048 29328 36100
rect 34520 36048 34572 36100
rect 37464 36048 37516 36100
rect 16120 35980 16172 36032
rect 18788 35980 18840 36032
rect 22468 36023 22520 36032
rect 22468 35989 22477 36023
rect 22477 35989 22511 36023
rect 22511 35989 22520 36023
rect 22468 35980 22520 35989
rect 26792 35980 26844 36032
rect 29092 35980 29144 36032
rect 36084 35980 36136 36032
rect 37832 35980 37884 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 7104 35819 7156 35828
rect 7104 35785 7113 35819
rect 7113 35785 7147 35819
rect 7147 35785 7156 35819
rect 7104 35776 7156 35785
rect 7748 35776 7800 35828
rect 11704 35819 11756 35828
rect 11704 35785 11713 35819
rect 11713 35785 11747 35819
rect 11747 35785 11756 35819
rect 11704 35776 11756 35785
rect 11888 35776 11940 35828
rect 13268 35776 13320 35828
rect 8300 35708 8352 35760
rect 9312 35708 9364 35760
rect 9956 35683 10008 35692
rect 9956 35649 9965 35683
rect 9965 35649 9999 35683
rect 9999 35649 10008 35683
rect 9956 35640 10008 35649
rect 11612 35640 11664 35692
rect 12164 35640 12216 35692
rect 13360 35683 13412 35692
rect 13360 35649 13369 35683
rect 13369 35649 13403 35683
rect 13403 35649 13412 35683
rect 13360 35640 13412 35649
rect 14740 35640 14792 35692
rect 16488 35640 16540 35692
rect 17684 35683 17736 35692
rect 17684 35649 17693 35683
rect 17693 35649 17727 35683
rect 17727 35649 17736 35683
rect 17684 35640 17736 35649
rect 18788 35683 18840 35692
rect 18788 35649 18797 35683
rect 18797 35649 18831 35683
rect 18831 35649 18840 35683
rect 18788 35640 18840 35649
rect 19892 35640 19944 35692
rect 7656 35615 7708 35624
rect 7656 35581 7665 35615
rect 7665 35581 7699 35615
rect 7699 35581 7708 35615
rect 7656 35572 7708 35581
rect 10048 35615 10100 35624
rect 10048 35581 10057 35615
rect 10057 35581 10091 35615
rect 10091 35581 10100 35615
rect 10048 35572 10100 35581
rect 13636 35615 13688 35624
rect 9404 35504 9456 35556
rect 13636 35581 13645 35615
rect 13645 35581 13679 35615
rect 13679 35581 13688 35615
rect 13636 35572 13688 35581
rect 17960 35615 18012 35624
rect 17960 35581 17969 35615
rect 17969 35581 18003 35615
rect 18003 35581 18012 35615
rect 17960 35572 18012 35581
rect 19156 35572 19208 35624
rect 13268 35504 13320 35556
rect 18420 35504 18472 35556
rect 19708 35504 19760 35556
rect 20444 35683 20496 35692
rect 20444 35649 20453 35683
rect 20453 35649 20487 35683
rect 20487 35649 20496 35683
rect 20444 35640 20496 35649
rect 22100 35776 22152 35828
rect 22928 35776 22980 35828
rect 23204 35776 23256 35828
rect 34520 35776 34572 35828
rect 36452 35776 36504 35828
rect 37464 35819 37516 35828
rect 37464 35785 37473 35819
rect 37473 35785 37507 35819
rect 37507 35785 37516 35819
rect 37464 35776 37516 35785
rect 20628 35708 20680 35760
rect 21364 35572 21416 35624
rect 22468 35640 22520 35692
rect 22928 35640 22980 35692
rect 23204 35683 23256 35692
rect 23204 35649 23213 35683
rect 23213 35649 23247 35683
rect 23247 35649 23256 35683
rect 23204 35640 23256 35649
rect 26424 35708 26476 35760
rect 32036 35708 32088 35760
rect 35624 35708 35676 35760
rect 24952 35683 25004 35692
rect 24952 35649 24961 35683
rect 24961 35649 24995 35683
rect 24995 35649 25004 35683
rect 24952 35640 25004 35649
rect 26516 35640 26568 35692
rect 27252 35683 27304 35692
rect 27252 35649 27261 35683
rect 27261 35649 27295 35683
rect 27295 35649 27304 35683
rect 27252 35640 27304 35649
rect 28632 35683 28684 35692
rect 28632 35649 28641 35683
rect 28641 35649 28675 35683
rect 28675 35649 28684 35683
rect 28632 35640 28684 35649
rect 28908 35683 28960 35692
rect 28908 35649 28942 35683
rect 28942 35649 28960 35683
rect 28908 35640 28960 35649
rect 32680 35640 32732 35692
rect 32956 35683 33008 35692
rect 32956 35649 32965 35683
rect 32965 35649 32999 35683
rect 32999 35649 33008 35683
rect 32956 35640 33008 35649
rect 33048 35683 33100 35692
rect 33048 35649 33057 35683
rect 33057 35649 33091 35683
rect 33091 35649 33100 35683
rect 33048 35640 33100 35649
rect 33784 35683 33836 35692
rect 24860 35615 24912 35624
rect 24860 35581 24869 35615
rect 24869 35581 24903 35615
rect 24903 35581 24912 35615
rect 24860 35572 24912 35581
rect 25412 35615 25464 35624
rect 25412 35581 25421 35615
rect 25421 35581 25455 35615
rect 25455 35581 25464 35615
rect 25412 35572 25464 35581
rect 26240 35572 26292 35624
rect 27528 35615 27580 35624
rect 27528 35581 27537 35615
rect 27537 35581 27571 35615
rect 27571 35581 27580 35615
rect 27528 35572 27580 35581
rect 27804 35572 27856 35624
rect 33784 35649 33793 35683
rect 33793 35649 33827 35683
rect 33827 35649 33836 35683
rect 33784 35640 33836 35649
rect 35992 35640 36044 35692
rect 37832 35683 37884 35692
rect 37832 35649 37841 35683
rect 37841 35649 37875 35683
rect 37875 35649 37884 35683
rect 37832 35640 37884 35649
rect 26332 35547 26384 35556
rect 9588 35479 9640 35488
rect 9588 35445 9597 35479
rect 9597 35445 9631 35479
rect 9631 35445 9640 35479
rect 9588 35436 9640 35445
rect 14832 35436 14884 35488
rect 16580 35436 16632 35488
rect 16948 35479 17000 35488
rect 16948 35445 16957 35479
rect 16957 35445 16991 35479
rect 16991 35445 17000 35479
rect 16948 35436 17000 35445
rect 19892 35436 19944 35488
rect 20168 35436 20220 35488
rect 20536 35436 20588 35488
rect 26332 35513 26341 35547
rect 26341 35513 26375 35547
rect 26375 35513 26384 35547
rect 26332 35504 26384 35513
rect 37740 35572 37792 35624
rect 38016 35615 38068 35624
rect 38016 35581 38025 35615
rect 38025 35581 38059 35615
rect 38059 35581 38068 35615
rect 38016 35572 38068 35581
rect 23664 35436 23716 35488
rect 24676 35436 24728 35488
rect 26424 35436 26476 35488
rect 28540 35436 28592 35488
rect 30012 35479 30064 35488
rect 30012 35445 30021 35479
rect 30021 35445 30055 35479
rect 30055 35445 30064 35479
rect 30012 35436 30064 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 10048 35232 10100 35284
rect 14740 35232 14792 35284
rect 18420 35232 18472 35284
rect 19984 35232 20036 35284
rect 23572 35275 23624 35284
rect 23572 35241 23581 35275
rect 23581 35241 23615 35275
rect 23615 35241 23624 35275
rect 23572 35232 23624 35241
rect 24860 35232 24912 35284
rect 28908 35232 28960 35284
rect 31208 35232 31260 35284
rect 32588 35232 32640 35284
rect 32864 35232 32916 35284
rect 33048 35275 33100 35284
rect 33048 35241 33057 35275
rect 33057 35241 33091 35275
rect 33091 35241 33100 35275
rect 33048 35232 33100 35241
rect 33784 35232 33836 35284
rect 11336 35207 11388 35216
rect 11336 35173 11345 35207
rect 11345 35173 11379 35207
rect 11379 35173 11388 35207
rect 11336 35164 11388 35173
rect 11888 35164 11940 35216
rect 7656 35096 7708 35148
rect 12716 35139 12768 35148
rect 12716 35105 12725 35139
rect 12725 35105 12759 35139
rect 12759 35105 12768 35139
rect 12716 35096 12768 35105
rect 9680 35028 9732 35080
rect 13084 35096 13136 35148
rect 19340 35164 19392 35216
rect 15752 35096 15804 35148
rect 19892 35096 19944 35148
rect 31668 35164 31720 35216
rect 23572 35096 23624 35148
rect 23848 35096 23900 35148
rect 29092 35139 29144 35148
rect 29092 35105 29101 35139
rect 29101 35105 29135 35139
rect 29135 35105 29144 35139
rect 29092 35096 29144 35105
rect 13544 35028 13596 35080
rect 15200 35028 15252 35080
rect 18236 35071 18288 35080
rect 18236 35037 18245 35071
rect 18245 35037 18279 35071
rect 18279 35037 18288 35071
rect 18236 35028 18288 35037
rect 19800 35071 19852 35080
rect 19800 35037 19809 35071
rect 19809 35037 19843 35071
rect 19843 35037 19852 35071
rect 19800 35028 19852 35037
rect 32128 35096 32180 35148
rect 5724 34960 5776 35012
rect 9588 34960 9640 35012
rect 11612 35003 11664 35012
rect 11612 34969 11621 35003
rect 11621 34969 11655 35003
rect 11655 34969 11664 35003
rect 11612 34960 11664 34969
rect 11796 35003 11848 35012
rect 11796 34969 11805 35003
rect 11805 34969 11839 35003
rect 11839 34969 11848 35003
rect 11796 34960 11848 34969
rect 11888 35003 11940 35012
rect 11888 34969 11897 35003
rect 11897 34969 11931 35003
rect 11931 34969 11940 35003
rect 11888 34960 11940 34969
rect 15936 34960 15988 35012
rect 16948 34960 17000 35012
rect 18420 34960 18472 35012
rect 19064 34960 19116 35012
rect 5080 34935 5132 34944
rect 5080 34901 5089 34935
rect 5089 34901 5123 34935
rect 5123 34901 5132 34935
rect 5080 34892 5132 34901
rect 5540 34935 5592 34944
rect 5540 34901 5549 34935
rect 5549 34901 5583 34935
rect 5583 34901 5592 34935
rect 5540 34892 5592 34901
rect 12716 34892 12768 34944
rect 19156 34892 19208 34944
rect 19432 34892 19484 34944
rect 19984 35003 20036 35012
rect 19984 34969 19993 35003
rect 19993 34969 20027 35003
rect 20027 34969 20036 35003
rect 20904 35028 20956 35080
rect 22008 35028 22060 35080
rect 19984 34960 20036 34969
rect 23204 35071 23256 35080
rect 23204 35037 23213 35071
rect 23213 35037 23247 35071
rect 23247 35037 23256 35071
rect 23204 35028 23256 35037
rect 24952 35028 25004 35080
rect 27160 35028 27212 35080
rect 27436 35071 27488 35080
rect 27436 35037 27446 35071
rect 27446 35037 27480 35071
rect 27480 35037 27488 35071
rect 27436 35028 27488 35037
rect 23664 34960 23716 35012
rect 25136 35003 25188 35012
rect 25136 34969 25145 35003
rect 25145 34969 25179 35003
rect 25179 34969 25188 35003
rect 25136 34960 25188 34969
rect 28908 35071 28960 35080
rect 28908 35037 28917 35071
rect 28917 35037 28951 35071
rect 28951 35037 28960 35071
rect 30656 35071 30708 35080
rect 28908 35028 28960 35037
rect 30656 35037 30665 35071
rect 30665 35037 30699 35071
rect 30699 35037 30708 35071
rect 30656 35028 30708 35037
rect 30748 35071 30800 35080
rect 30748 35037 30758 35071
rect 30758 35037 30792 35071
rect 30792 35037 30800 35071
rect 31024 35071 31076 35080
rect 30748 35028 30800 35037
rect 31024 35037 31033 35071
rect 31033 35037 31067 35071
rect 31067 35037 31076 35071
rect 31024 35028 31076 35037
rect 31668 35028 31720 35080
rect 31760 35071 31812 35080
rect 31760 35037 31769 35071
rect 31769 35037 31803 35071
rect 31803 35037 31812 35071
rect 31944 35071 31996 35080
rect 31760 35028 31812 35037
rect 31944 35037 31951 35071
rect 31951 35037 31996 35071
rect 31944 35028 31996 35037
rect 36268 35139 36320 35148
rect 36268 35105 36277 35139
rect 36277 35105 36311 35139
rect 36311 35105 36320 35139
rect 36268 35096 36320 35105
rect 29184 34960 29236 35012
rect 32312 34960 32364 35012
rect 34704 35028 34756 35080
rect 32956 34960 33008 35012
rect 36176 34960 36228 35012
rect 20444 34892 20496 34944
rect 21088 34935 21140 34944
rect 21088 34901 21097 34935
rect 21097 34901 21131 34935
rect 21131 34901 21140 34935
rect 21088 34892 21140 34901
rect 22744 34892 22796 34944
rect 24676 34892 24728 34944
rect 27712 34935 27764 34944
rect 27712 34901 27721 34935
rect 27721 34901 27755 34935
rect 27755 34901 27764 34935
rect 27712 34892 27764 34901
rect 31116 34892 31168 34944
rect 31852 34892 31904 34944
rect 32680 34892 32732 34944
rect 35440 34892 35492 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4620 34688 4672 34740
rect 5540 34688 5592 34740
rect 7012 34688 7064 34740
rect 10048 34731 10100 34740
rect 10048 34697 10057 34731
rect 10057 34697 10091 34731
rect 10091 34697 10100 34731
rect 10048 34688 10100 34697
rect 19156 34688 19208 34740
rect 20444 34731 20496 34740
rect 5080 34552 5132 34604
rect 8300 34620 8352 34672
rect 9956 34663 10008 34672
rect 9956 34629 9965 34663
rect 9965 34629 9999 34663
rect 9999 34629 10008 34663
rect 9956 34620 10008 34629
rect 16028 34620 16080 34672
rect 7748 34552 7800 34604
rect 7840 34595 7892 34604
rect 7840 34561 7849 34595
rect 7849 34561 7883 34595
rect 7883 34561 7892 34595
rect 7840 34552 7892 34561
rect 18236 34595 18288 34604
rect 5908 34416 5960 34468
rect 7748 34416 7800 34468
rect 11888 34484 11940 34536
rect 17408 34484 17460 34536
rect 18236 34561 18245 34595
rect 18245 34561 18279 34595
rect 18279 34561 18288 34595
rect 18236 34552 18288 34561
rect 19432 34620 19484 34672
rect 20076 34620 20128 34672
rect 20444 34697 20453 34731
rect 20453 34697 20487 34731
rect 20487 34697 20496 34731
rect 20444 34688 20496 34697
rect 20904 34620 20956 34672
rect 23848 34688 23900 34740
rect 30748 34688 30800 34740
rect 33692 34688 33744 34740
rect 36176 34731 36228 34740
rect 36176 34697 36185 34731
rect 36185 34697 36219 34731
rect 36219 34697 36228 34731
rect 36176 34688 36228 34697
rect 21364 34620 21416 34672
rect 17960 34484 18012 34536
rect 19064 34484 19116 34536
rect 18420 34416 18472 34468
rect 19892 34484 19944 34536
rect 21824 34552 21876 34604
rect 22008 34595 22060 34604
rect 22008 34561 22017 34595
rect 22017 34561 22051 34595
rect 22051 34561 22060 34595
rect 22008 34552 22060 34561
rect 22376 34552 22428 34604
rect 24676 34552 24728 34604
rect 25688 34552 25740 34604
rect 27160 34595 27212 34604
rect 27160 34561 27169 34595
rect 27169 34561 27203 34595
rect 27203 34561 27212 34595
rect 27160 34552 27212 34561
rect 27436 34620 27488 34672
rect 28540 34552 28592 34604
rect 29092 34595 29144 34604
rect 29092 34561 29101 34595
rect 29101 34561 29135 34595
rect 29135 34561 29144 34595
rect 29092 34552 29144 34561
rect 32956 34552 33008 34604
rect 22284 34484 22336 34536
rect 23204 34484 23256 34536
rect 23664 34527 23716 34536
rect 23664 34493 23673 34527
rect 23673 34493 23707 34527
rect 23707 34493 23716 34527
rect 23664 34484 23716 34493
rect 25872 34527 25924 34536
rect 25872 34493 25881 34527
rect 25881 34493 25915 34527
rect 25915 34493 25924 34527
rect 25872 34484 25924 34493
rect 29184 34484 29236 34536
rect 32864 34484 32916 34536
rect 34244 34552 34296 34604
rect 35440 34552 35492 34604
rect 36636 34527 36688 34536
rect 36636 34493 36645 34527
rect 36645 34493 36679 34527
rect 36679 34493 36688 34527
rect 36636 34484 36688 34493
rect 38108 34527 38160 34536
rect 20260 34416 20312 34468
rect 23572 34416 23624 34468
rect 38108 34493 38117 34527
rect 38117 34493 38151 34527
rect 38151 34493 38160 34527
rect 38108 34484 38160 34493
rect 38016 34416 38068 34468
rect 17960 34348 18012 34400
rect 18144 34391 18196 34400
rect 18144 34357 18153 34391
rect 18153 34357 18187 34391
rect 18187 34357 18196 34391
rect 18144 34348 18196 34357
rect 18236 34348 18288 34400
rect 19892 34348 19944 34400
rect 22376 34391 22428 34400
rect 22376 34357 22385 34391
rect 22385 34357 22419 34391
rect 22419 34357 22428 34391
rect 22376 34348 22428 34357
rect 22652 34391 22704 34400
rect 22652 34357 22661 34391
rect 22661 34357 22695 34391
rect 22695 34357 22704 34391
rect 22652 34348 22704 34357
rect 25136 34348 25188 34400
rect 29000 34348 29052 34400
rect 30748 34348 30800 34400
rect 35348 34348 35400 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 10232 34144 10284 34196
rect 5540 34008 5592 34060
rect 5908 34051 5960 34060
rect 5908 34017 5917 34051
rect 5917 34017 5951 34051
rect 5951 34017 5960 34051
rect 8208 34051 8260 34060
rect 5908 34008 5960 34017
rect 8208 34017 8217 34051
rect 8217 34017 8251 34051
rect 8251 34017 8260 34051
rect 8208 34008 8260 34017
rect 9680 34008 9732 34060
rect 11336 34008 11388 34060
rect 5724 33983 5776 33992
rect 5724 33949 5733 33983
rect 5733 33949 5767 33983
rect 5767 33949 5776 33983
rect 5724 33940 5776 33949
rect 7748 33983 7800 33992
rect 7748 33949 7757 33983
rect 7757 33949 7791 33983
rect 7791 33949 7800 33983
rect 7748 33940 7800 33949
rect 10600 33940 10652 33992
rect 11152 33940 11204 33992
rect 11888 33983 11940 33992
rect 11888 33949 11897 33983
rect 11897 33949 11931 33983
rect 11931 33949 11940 33983
rect 11888 33940 11940 33949
rect 12256 33940 12308 33992
rect 14648 33940 14700 33992
rect 15844 33940 15896 33992
rect 17684 34008 17736 34060
rect 20904 34144 20956 34196
rect 21732 34144 21784 34196
rect 23020 34144 23072 34196
rect 23848 34144 23900 34196
rect 25412 34144 25464 34196
rect 25780 34187 25832 34196
rect 25780 34153 25789 34187
rect 25789 34153 25823 34187
rect 25823 34153 25832 34187
rect 25780 34144 25832 34153
rect 27252 34144 27304 34196
rect 31760 34144 31812 34196
rect 31852 34187 31904 34196
rect 31852 34153 31861 34187
rect 31861 34153 31895 34187
rect 31895 34153 31904 34187
rect 31852 34144 31904 34153
rect 18604 34076 18656 34128
rect 26700 34119 26752 34128
rect 8484 33872 8536 33924
rect 9128 33915 9180 33924
rect 9128 33881 9137 33915
rect 9137 33881 9171 33915
rect 9171 33881 9180 33915
rect 9128 33872 9180 33881
rect 16580 33872 16632 33924
rect 5356 33847 5408 33856
rect 5356 33813 5365 33847
rect 5365 33813 5399 33847
rect 5399 33813 5408 33847
rect 5356 33804 5408 33813
rect 14096 33804 14148 33856
rect 15476 33804 15528 33856
rect 17592 33804 17644 33856
rect 17960 33872 18012 33924
rect 19524 34008 19576 34060
rect 19248 33940 19300 33992
rect 21548 34008 21600 34060
rect 22284 34008 22336 34060
rect 25872 34051 25924 34060
rect 20260 33983 20312 33992
rect 19064 33872 19116 33924
rect 20260 33949 20269 33983
rect 20269 33949 20303 33983
rect 20303 33949 20312 33983
rect 20260 33940 20312 33949
rect 22376 33983 22428 33992
rect 20812 33872 20864 33924
rect 19432 33804 19484 33856
rect 19984 33804 20036 33856
rect 20260 33804 20312 33856
rect 20720 33804 20772 33856
rect 21640 33915 21692 33924
rect 21640 33881 21649 33915
rect 21649 33881 21683 33915
rect 21683 33881 21692 33915
rect 22376 33949 22385 33983
rect 22385 33949 22419 33983
rect 22419 33949 22428 33983
rect 22376 33940 22428 33949
rect 21640 33872 21692 33881
rect 22192 33872 22244 33924
rect 22652 33940 22704 33992
rect 22744 33983 22796 33992
rect 22744 33949 22753 33983
rect 22753 33949 22787 33983
rect 22787 33949 22796 33983
rect 23572 33983 23624 33992
rect 22744 33940 22796 33949
rect 23572 33949 23581 33983
rect 23581 33949 23615 33983
rect 23615 33949 23624 33983
rect 23572 33940 23624 33949
rect 23848 33983 23900 33992
rect 23848 33949 23857 33983
rect 23857 33949 23891 33983
rect 23891 33949 23900 33983
rect 23848 33940 23900 33949
rect 24768 33983 24820 33992
rect 24768 33949 24777 33983
rect 24777 33949 24811 33983
rect 24811 33949 24820 33983
rect 24768 33940 24820 33949
rect 22284 33804 22336 33856
rect 23020 33872 23072 33924
rect 25044 33940 25096 33992
rect 25872 34017 25881 34051
rect 25881 34017 25915 34051
rect 25915 34017 25924 34051
rect 25872 34008 25924 34017
rect 26700 34085 26709 34119
rect 26709 34085 26743 34119
rect 26743 34085 26752 34119
rect 26700 34076 26752 34085
rect 27344 33940 27396 33992
rect 27712 33940 27764 33992
rect 25596 33872 25648 33924
rect 22744 33804 22796 33856
rect 25688 33804 25740 33856
rect 26792 33872 26844 33924
rect 27896 33915 27948 33924
rect 27896 33881 27905 33915
rect 27905 33881 27939 33915
rect 27939 33881 27948 33915
rect 27896 33872 27948 33881
rect 29000 34008 29052 34060
rect 29276 34008 29328 34060
rect 29184 33983 29236 33992
rect 29184 33949 29193 33983
rect 29193 33949 29227 33983
rect 29227 33949 29236 33983
rect 29184 33940 29236 33949
rect 29644 33940 29696 33992
rect 31944 34076 31996 34128
rect 35256 34144 35308 34196
rect 35440 34144 35492 34196
rect 33048 34076 33100 34128
rect 37832 34076 37884 34128
rect 30196 33983 30248 33992
rect 30196 33949 30210 33983
rect 30210 33949 30244 33983
rect 30244 33949 30248 33983
rect 31208 33983 31260 33992
rect 30196 33940 30248 33949
rect 31208 33949 31217 33983
rect 31217 33949 31251 33983
rect 31251 33949 31260 33983
rect 31208 33940 31260 33949
rect 31300 33983 31352 33992
rect 31300 33949 31310 33983
rect 31310 33949 31344 33983
rect 31344 33949 31352 33983
rect 36084 34008 36136 34060
rect 31668 33983 31720 33992
rect 31300 33940 31352 33949
rect 31668 33949 31682 33983
rect 31682 33949 31716 33983
rect 31716 33949 31720 33983
rect 31668 33940 31720 33949
rect 37188 33940 37240 33992
rect 30012 33915 30064 33924
rect 26516 33804 26568 33856
rect 28724 33847 28776 33856
rect 28724 33813 28733 33847
rect 28733 33813 28767 33847
rect 28767 33813 28776 33847
rect 28724 33804 28776 33813
rect 30012 33881 30021 33915
rect 30021 33881 30055 33915
rect 30055 33881 30064 33915
rect 30012 33872 30064 33881
rect 30104 33915 30156 33924
rect 30104 33881 30113 33915
rect 30113 33881 30147 33915
rect 30147 33881 30156 33915
rect 30104 33872 30156 33881
rect 31116 33872 31168 33924
rect 34520 33872 34572 33924
rect 38108 33915 38160 33924
rect 38108 33881 38117 33915
rect 38117 33881 38151 33915
rect 38151 33881 38160 33915
rect 38108 33872 38160 33881
rect 32680 33804 32732 33856
rect 35532 33804 35584 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 13636 33600 13688 33652
rect 14648 33643 14700 33652
rect 14648 33609 14657 33643
rect 14657 33609 14691 33643
rect 14691 33609 14700 33643
rect 14648 33600 14700 33609
rect 16212 33600 16264 33652
rect 17500 33600 17552 33652
rect 19340 33600 19392 33652
rect 21640 33600 21692 33652
rect 22744 33600 22796 33652
rect 24216 33600 24268 33652
rect 27344 33600 27396 33652
rect 28724 33600 28776 33652
rect 31116 33600 31168 33652
rect 32864 33600 32916 33652
rect 5172 33464 5224 33516
rect 7380 33532 7432 33584
rect 8484 33532 8536 33584
rect 9312 33532 9364 33584
rect 6552 33464 6604 33516
rect 7012 33507 7064 33516
rect 7012 33473 7021 33507
rect 7021 33473 7055 33507
rect 7055 33473 7064 33507
rect 7012 33464 7064 33473
rect 8116 33507 8168 33516
rect 8116 33473 8125 33507
rect 8125 33473 8159 33507
rect 8159 33473 8168 33507
rect 8116 33464 8168 33473
rect 8392 33464 8444 33516
rect 12072 33507 12124 33516
rect 7472 33396 7524 33448
rect 12072 33473 12081 33507
rect 12081 33473 12115 33507
rect 12115 33473 12124 33507
rect 12072 33464 12124 33473
rect 12256 33507 12308 33516
rect 12256 33473 12265 33507
rect 12265 33473 12299 33507
rect 12299 33473 12308 33507
rect 12256 33464 12308 33473
rect 11336 33396 11388 33448
rect 14188 33464 14240 33516
rect 14556 33464 14608 33516
rect 15016 33464 15068 33516
rect 15384 33507 15436 33516
rect 15384 33473 15393 33507
rect 15393 33473 15427 33507
rect 15427 33473 15436 33507
rect 15384 33464 15436 33473
rect 13544 33396 13596 33448
rect 14372 33439 14424 33448
rect 14372 33405 14381 33439
rect 14381 33405 14415 33439
rect 14415 33405 14424 33439
rect 14372 33396 14424 33405
rect 14648 33396 14700 33448
rect 17408 33507 17460 33516
rect 17408 33473 17417 33507
rect 17417 33473 17451 33507
rect 17451 33473 17460 33507
rect 17408 33464 17460 33473
rect 16948 33396 17000 33448
rect 17776 33396 17828 33448
rect 18236 33464 18288 33516
rect 15200 33328 15252 33380
rect 15844 33328 15896 33380
rect 17500 33328 17552 33380
rect 6828 33260 6880 33312
rect 9956 33260 10008 33312
rect 14096 33303 14148 33312
rect 14096 33269 14105 33303
rect 14105 33269 14139 33303
rect 14139 33269 14148 33303
rect 14096 33260 14148 33269
rect 14188 33260 14240 33312
rect 14832 33260 14884 33312
rect 15476 33303 15528 33312
rect 15476 33269 15485 33303
rect 15485 33269 15519 33303
rect 15519 33269 15528 33303
rect 15476 33260 15528 33269
rect 19156 33396 19208 33448
rect 19340 33507 19392 33516
rect 19340 33473 19349 33507
rect 19349 33473 19383 33507
rect 19383 33473 19392 33507
rect 23388 33532 23440 33584
rect 19340 33464 19392 33473
rect 19432 33396 19484 33448
rect 19800 33464 19852 33516
rect 20352 33464 20404 33516
rect 21272 33507 21324 33516
rect 21272 33473 21281 33507
rect 21281 33473 21315 33507
rect 21315 33473 21324 33507
rect 21272 33464 21324 33473
rect 22468 33507 22520 33516
rect 22468 33473 22477 33507
rect 22477 33473 22511 33507
rect 22511 33473 22520 33507
rect 22744 33507 22796 33516
rect 22468 33464 22520 33473
rect 22744 33473 22753 33507
rect 22753 33473 22787 33507
rect 22787 33473 22796 33507
rect 22744 33464 22796 33473
rect 25136 33532 25188 33584
rect 22100 33396 22152 33448
rect 24216 33507 24268 33516
rect 24216 33473 24225 33507
rect 24225 33473 24259 33507
rect 24259 33473 24268 33507
rect 24216 33464 24268 33473
rect 20352 33328 20404 33380
rect 19248 33260 19300 33312
rect 20812 33260 20864 33312
rect 20904 33260 20956 33312
rect 21456 33260 21508 33312
rect 23756 33396 23808 33448
rect 24032 33439 24084 33448
rect 24032 33405 24041 33439
rect 24041 33405 24075 33439
rect 24075 33405 24084 33439
rect 24032 33396 24084 33405
rect 24768 33464 24820 33516
rect 26240 33507 26292 33516
rect 23204 33328 23256 33380
rect 26240 33473 26249 33507
rect 26249 33473 26283 33507
rect 26283 33473 26292 33507
rect 26240 33464 26292 33473
rect 26424 33507 26476 33516
rect 26424 33473 26433 33507
rect 26433 33473 26467 33507
rect 26467 33473 26476 33507
rect 26424 33464 26476 33473
rect 30932 33532 30984 33584
rect 31392 33575 31444 33584
rect 31392 33541 31401 33575
rect 31401 33541 31435 33575
rect 31435 33541 31444 33575
rect 31392 33532 31444 33541
rect 32680 33532 32732 33584
rect 35716 33600 35768 33652
rect 36636 33600 36688 33652
rect 33692 33532 33744 33584
rect 34704 33575 34756 33584
rect 34704 33541 34709 33575
rect 34709 33541 34743 33575
rect 34743 33541 34756 33575
rect 34704 33532 34756 33541
rect 27620 33464 27672 33516
rect 31024 33507 31076 33516
rect 24860 33328 24912 33380
rect 26884 33396 26936 33448
rect 27988 33396 28040 33448
rect 27436 33328 27488 33380
rect 29092 33328 29144 33380
rect 31024 33473 31033 33507
rect 31033 33473 31067 33507
rect 31067 33473 31076 33507
rect 31024 33464 31076 33473
rect 29828 33396 29880 33448
rect 30748 33396 30800 33448
rect 31484 33507 31536 33516
rect 31484 33473 31498 33507
rect 31498 33473 31532 33507
rect 31532 33473 31536 33507
rect 32864 33507 32916 33516
rect 31484 33464 31536 33473
rect 32864 33473 32873 33507
rect 32873 33473 32907 33507
rect 32907 33473 32916 33507
rect 32864 33464 32916 33473
rect 29920 33328 29972 33380
rect 33048 33464 33100 33516
rect 34336 33464 34388 33516
rect 34428 33507 34480 33516
rect 34428 33473 34437 33507
rect 34437 33473 34471 33507
rect 34471 33473 34480 33507
rect 34428 33464 34480 33473
rect 34612 33464 34664 33516
rect 34888 33464 34940 33516
rect 35716 33507 35768 33516
rect 35256 33396 35308 33448
rect 35716 33473 35725 33507
rect 35725 33473 35759 33507
rect 35759 33473 35768 33507
rect 35716 33464 35768 33473
rect 35624 33396 35676 33448
rect 35900 33507 35952 33516
rect 35900 33473 35914 33507
rect 35914 33473 35948 33507
rect 35948 33473 35952 33507
rect 35900 33464 35952 33473
rect 36176 33464 36228 33516
rect 37832 33507 37884 33516
rect 37832 33473 37841 33507
rect 37841 33473 37875 33507
rect 37875 33473 37884 33507
rect 37832 33464 37884 33473
rect 36360 33396 36412 33448
rect 37188 33396 37240 33448
rect 38016 33439 38068 33448
rect 38016 33405 38025 33439
rect 38025 33405 38059 33439
rect 38059 33405 38068 33439
rect 38016 33396 38068 33405
rect 23756 33260 23808 33312
rect 25780 33260 25832 33312
rect 37740 33328 37792 33380
rect 37096 33260 37148 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 10232 33056 10284 33108
rect 8116 32988 8168 33040
rect 9680 32988 9732 33040
rect 13544 33056 13596 33108
rect 13728 33056 13780 33108
rect 15660 33056 15712 33108
rect 15844 33099 15896 33108
rect 15844 33065 15853 33099
rect 15853 33065 15887 33099
rect 15887 33065 15896 33099
rect 15844 33056 15896 33065
rect 15936 33056 15988 33108
rect 18052 33056 18104 33108
rect 18144 33056 18196 33108
rect 18328 33099 18380 33108
rect 18328 33065 18337 33099
rect 18337 33065 18371 33099
rect 18371 33065 18380 33099
rect 18328 33056 18380 33065
rect 20168 33056 20220 33108
rect 20352 33056 20404 33108
rect 20536 33056 20588 33108
rect 22652 33056 22704 33108
rect 25228 33099 25280 33108
rect 25228 33065 25237 33099
rect 25237 33065 25271 33099
rect 25271 33065 25280 33099
rect 25228 33056 25280 33065
rect 30656 33056 30708 33108
rect 31208 33056 31260 33108
rect 32864 33056 32916 33108
rect 35716 33056 35768 33108
rect 36360 33099 36412 33108
rect 4620 32920 4672 32972
rect 5356 32920 5408 32972
rect 5816 32920 5868 32972
rect 4528 32895 4580 32904
rect 4528 32861 4537 32895
rect 4537 32861 4571 32895
rect 4571 32861 4580 32895
rect 5172 32895 5224 32904
rect 4528 32852 4580 32861
rect 5172 32861 5181 32895
rect 5181 32861 5215 32895
rect 5215 32861 5224 32895
rect 5172 32852 5224 32861
rect 5264 32895 5316 32904
rect 5264 32861 5273 32895
rect 5273 32861 5307 32895
rect 5307 32861 5316 32895
rect 5264 32852 5316 32861
rect 7380 32895 7432 32904
rect 4712 32827 4764 32836
rect 4712 32793 4721 32827
rect 4721 32793 4755 32827
rect 4755 32793 4764 32827
rect 4712 32784 4764 32793
rect 5724 32827 5776 32836
rect 5724 32793 5733 32827
rect 5733 32793 5767 32827
rect 5767 32793 5776 32827
rect 5724 32784 5776 32793
rect 7380 32861 7389 32895
rect 7389 32861 7423 32895
rect 7423 32861 7432 32895
rect 7380 32852 7432 32861
rect 7748 32852 7800 32904
rect 8392 32920 8444 32972
rect 9772 32920 9824 32972
rect 10140 32920 10192 32972
rect 9220 32852 9272 32904
rect 9864 32895 9916 32904
rect 9864 32861 9873 32895
rect 9873 32861 9907 32895
rect 9907 32861 9916 32895
rect 9864 32852 9916 32861
rect 10232 32895 10284 32904
rect 7472 32784 7524 32836
rect 10232 32861 10241 32895
rect 10241 32861 10275 32895
rect 10275 32861 10284 32895
rect 10232 32852 10284 32861
rect 11244 32920 11296 32972
rect 11152 32895 11204 32904
rect 9588 32716 9640 32768
rect 10416 32759 10468 32768
rect 10416 32725 10425 32759
rect 10425 32725 10459 32759
rect 10459 32725 10468 32759
rect 10416 32716 10468 32725
rect 10600 32784 10652 32836
rect 11152 32861 11161 32895
rect 11161 32861 11195 32895
rect 11195 32861 11204 32895
rect 11152 32852 11204 32861
rect 13360 32920 13412 32972
rect 15384 32920 15436 32972
rect 12256 32895 12308 32904
rect 12256 32861 12265 32895
rect 12265 32861 12299 32895
rect 12299 32861 12308 32895
rect 12256 32852 12308 32861
rect 12532 32895 12584 32904
rect 11980 32784 12032 32836
rect 12532 32861 12541 32895
rect 12541 32861 12575 32895
rect 12575 32861 12584 32895
rect 12532 32852 12584 32861
rect 13544 32895 13596 32904
rect 13544 32861 13553 32895
rect 13553 32861 13587 32895
rect 13587 32861 13596 32895
rect 13544 32852 13596 32861
rect 13728 32895 13780 32904
rect 13728 32861 13737 32895
rect 13737 32861 13771 32895
rect 13771 32861 13780 32895
rect 13728 32852 13780 32861
rect 15108 32852 15160 32904
rect 20720 32988 20772 33040
rect 22744 33031 22796 33040
rect 22744 32997 22753 33031
rect 22753 32997 22787 33031
rect 22787 32997 22796 33031
rect 22744 32988 22796 32997
rect 23388 32988 23440 33040
rect 26240 32988 26292 33040
rect 17776 32920 17828 32972
rect 17592 32895 17644 32904
rect 12808 32784 12860 32836
rect 13820 32784 13872 32836
rect 15200 32784 15252 32836
rect 17592 32861 17601 32895
rect 17601 32861 17635 32895
rect 17635 32861 17644 32895
rect 17592 32852 17644 32861
rect 17868 32852 17920 32904
rect 18144 32784 18196 32836
rect 20168 32852 20220 32904
rect 20536 32895 20588 32904
rect 20536 32861 20545 32895
rect 20545 32861 20579 32895
rect 20579 32861 20588 32895
rect 20536 32852 20588 32861
rect 21640 32920 21692 32972
rect 20720 32852 20772 32904
rect 22468 32920 22520 32972
rect 20904 32827 20956 32836
rect 20904 32793 20913 32827
rect 20913 32793 20947 32827
rect 20947 32793 20956 32827
rect 22560 32852 22612 32904
rect 23020 32920 23072 32972
rect 24952 32920 25004 32972
rect 30196 32988 30248 33040
rect 23572 32852 23624 32904
rect 23848 32852 23900 32904
rect 25964 32852 26016 32904
rect 28724 32963 28776 32972
rect 28724 32929 28733 32963
rect 28733 32929 28767 32963
rect 28767 32929 28776 32963
rect 28724 32920 28776 32929
rect 26240 32852 26292 32904
rect 20904 32784 20956 32793
rect 22744 32784 22796 32836
rect 25688 32784 25740 32836
rect 27988 32852 28040 32904
rect 28172 32852 28224 32904
rect 28908 32852 28960 32904
rect 29920 32895 29972 32904
rect 29920 32861 29927 32895
rect 29927 32861 29972 32895
rect 11060 32716 11112 32768
rect 14188 32716 14240 32768
rect 15660 32716 15712 32768
rect 18420 32716 18472 32768
rect 18696 32716 18748 32768
rect 19432 32716 19484 32768
rect 19800 32759 19852 32768
rect 19800 32725 19809 32759
rect 19809 32725 19843 32759
rect 19843 32725 19852 32759
rect 19800 32716 19852 32725
rect 19984 32716 20036 32768
rect 21272 32716 21324 32768
rect 21640 32716 21692 32768
rect 22652 32716 22704 32768
rect 23112 32759 23164 32768
rect 23112 32725 23121 32759
rect 23121 32725 23155 32759
rect 23155 32725 23164 32759
rect 23112 32716 23164 32725
rect 24216 32716 24268 32768
rect 24768 32716 24820 32768
rect 26976 32716 27028 32768
rect 29920 32852 29972 32861
rect 30104 32895 30156 32904
rect 30104 32861 30113 32895
rect 30113 32861 30147 32895
rect 30147 32861 30156 32895
rect 30104 32852 30156 32861
rect 29828 32716 29880 32768
rect 30380 32852 30432 32904
rect 31484 32920 31536 32972
rect 32128 32920 32180 32972
rect 31300 32895 31352 32904
rect 31300 32861 31314 32895
rect 31314 32861 31348 32895
rect 31348 32861 31352 32895
rect 31944 32895 31996 32904
rect 31300 32852 31352 32861
rect 31944 32861 31953 32895
rect 31953 32861 31987 32895
rect 31987 32861 31996 32895
rect 31944 32852 31996 32861
rect 32312 32895 32364 32904
rect 32312 32861 32321 32895
rect 32321 32861 32355 32895
rect 32355 32861 32364 32895
rect 32312 32852 32364 32861
rect 34520 32852 34572 32904
rect 35164 32852 35216 32904
rect 35440 32852 35492 32904
rect 36360 33065 36369 33099
rect 36369 33065 36403 33099
rect 36403 33065 36412 33099
rect 36360 33056 36412 33065
rect 36268 32988 36320 33040
rect 30104 32716 30156 32768
rect 30288 32716 30340 32768
rect 31300 32716 31352 32768
rect 31760 32784 31812 32836
rect 34888 32716 34940 32768
rect 36176 32895 36228 32904
rect 36176 32861 36190 32895
rect 36190 32861 36224 32895
rect 36224 32861 36228 32895
rect 37096 32895 37148 32904
rect 36176 32852 36228 32861
rect 37096 32861 37130 32895
rect 37130 32861 37148 32895
rect 37096 32852 37148 32861
rect 36084 32827 36136 32836
rect 36084 32793 36093 32827
rect 36093 32793 36127 32827
rect 36127 32793 36136 32827
rect 36084 32784 36136 32793
rect 37832 32716 37884 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 9220 32512 9272 32564
rect 9588 32555 9640 32564
rect 9588 32521 9597 32555
rect 9597 32521 9631 32555
rect 9631 32521 9640 32555
rect 9588 32512 9640 32521
rect 10416 32512 10468 32564
rect 4712 32444 4764 32496
rect 4620 32419 4672 32428
rect 4620 32385 4629 32419
rect 4629 32385 4663 32419
rect 4663 32385 4672 32419
rect 4620 32376 4672 32385
rect 7748 32444 7800 32496
rect 8208 32487 8260 32496
rect 8208 32453 8217 32487
rect 8217 32453 8251 32487
rect 8251 32453 8260 32487
rect 8208 32444 8260 32453
rect 8392 32487 8444 32496
rect 8392 32453 8401 32487
rect 8401 32453 8435 32487
rect 8435 32453 8444 32487
rect 8392 32444 8444 32453
rect 5724 32376 5776 32428
rect 6920 32376 6972 32428
rect 9220 32376 9272 32428
rect 9496 32419 9548 32428
rect 9496 32385 9505 32419
rect 9505 32385 9539 32419
rect 9539 32385 9548 32419
rect 11888 32444 11940 32496
rect 12256 32444 12308 32496
rect 14188 32487 14240 32496
rect 14188 32453 14197 32487
rect 14197 32453 14231 32487
rect 14231 32453 14240 32487
rect 14188 32444 14240 32453
rect 14372 32512 14424 32564
rect 16304 32512 16356 32564
rect 20444 32512 20496 32564
rect 20720 32555 20772 32564
rect 20720 32521 20729 32555
rect 20729 32521 20763 32555
rect 20763 32521 20772 32555
rect 20720 32512 20772 32521
rect 20904 32512 20956 32564
rect 16856 32487 16908 32496
rect 16856 32453 16865 32487
rect 16865 32453 16899 32487
rect 16899 32453 16908 32487
rect 16856 32444 16908 32453
rect 9496 32376 9548 32385
rect 4528 32308 4580 32360
rect 5448 32240 5500 32292
rect 6460 32308 6512 32360
rect 10232 32376 10284 32428
rect 12072 32419 12124 32428
rect 12072 32385 12081 32419
rect 12081 32385 12115 32419
rect 12115 32385 12124 32419
rect 12072 32376 12124 32385
rect 11980 32308 12032 32360
rect 12164 32308 12216 32360
rect 14556 32376 14608 32428
rect 14924 32376 14976 32428
rect 12624 32308 12676 32360
rect 12900 32351 12952 32360
rect 12900 32317 12909 32351
rect 12909 32317 12943 32351
rect 12943 32317 12952 32351
rect 12900 32308 12952 32317
rect 14372 32351 14424 32360
rect 14372 32317 14381 32351
rect 14381 32317 14415 32351
rect 14415 32317 14424 32351
rect 14372 32308 14424 32317
rect 14832 32308 14884 32360
rect 15384 32351 15436 32360
rect 15384 32317 15393 32351
rect 15393 32317 15427 32351
rect 15427 32317 15436 32351
rect 15384 32308 15436 32317
rect 15476 32351 15528 32360
rect 15476 32317 15485 32351
rect 15485 32317 15519 32351
rect 15519 32317 15528 32351
rect 16304 32376 16356 32428
rect 19708 32444 19760 32496
rect 20352 32444 20404 32496
rect 20628 32444 20680 32496
rect 17316 32419 17368 32428
rect 17316 32385 17325 32419
rect 17325 32385 17359 32419
rect 17359 32385 17368 32419
rect 17316 32376 17368 32385
rect 15476 32308 15528 32317
rect 17684 32376 17736 32428
rect 18144 32419 18196 32428
rect 18144 32385 18153 32419
rect 18153 32385 18187 32419
rect 18187 32385 18196 32419
rect 18144 32376 18196 32385
rect 20904 32376 20956 32428
rect 21824 32444 21876 32496
rect 22284 32512 22336 32564
rect 25964 32555 26016 32564
rect 25964 32521 25973 32555
rect 25973 32521 26007 32555
rect 26007 32521 26016 32555
rect 25964 32512 26016 32521
rect 31024 32512 31076 32564
rect 32312 32512 32364 32564
rect 34796 32512 34848 32564
rect 35256 32512 35308 32564
rect 35440 32555 35492 32564
rect 35440 32521 35449 32555
rect 35449 32521 35483 32555
rect 35483 32521 35492 32555
rect 35440 32512 35492 32521
rect 26148 32444 26200 32496
rect 19984 32308 20036 32360
rect 21180 32308 21232 32360
rect 22836 32376 22888 32428
rect 23020 32376 23072 32428
rect 24124 32419 24176 32428
rect 24124 32385 24133 32419
rect 24133 32385 24167 32419
rect 24167 32385 24176 32419
rect 24124 32376 24176 32385
rect 24216 32419 24268 32428
rect 24216 32385 24225 32419
rect 24225 32385 24259 32419
rect 24259 32385 24268 32419
rect 24216 32376 24268 32385
rect 25044 32376 25096 32428
rect 25688 32376 25740 32428
rect 26240 32376 26292 32428
rect 27528 32444 27580 32496
rect 28448 32419 28500 32428
rect 6736 32240 6788 32292
rect 8208 32240 8260 32292
rect 10324 32240 10376 32292
rect 6644 32172 6696 32224
rect 8300 32172 8352 32224
rect 9680 32172 9732 32224
rect 11060 32172 11112 32224
rect 11520 32240 11572 32292
rect 12348 32172 12400 32224
rect 12808 32215 12860 32224
rect 12808 32181 12817 32215
rect 12817 32181 12851 32215
rect 12851 32181 12860 32215
rect 12808 32172 12860 32181
rect 14188 32215 14240 32224
rect 14188 32181 14197 32215
rect 14197 32181 14231 32215
rect 14231 32181 14240 32215
rect 14188 32172 14240 32181
rect 18420 32240 18472 32292
rect 21824 32240 21876 32292
rect 15476 32172 15528 32224
rect 16212 32215 16264 32224
rect 16212 32181 16221 32215
rect 16221 32181 16255 32215
rect 16255 32181 16264 32215
rect 16212 32172 16264 32181
rect 16948 32215 17000 32224
rect 16948 32181 16957 32215
rect 16957 32181 16991 32215
rect 16991 32181 17000 32215
rect 16948 32172 17000 32181
rect 17408 32172 17460 32224
rect 17500 32215 17552 32224
rect 17500 32181 17509 32215
rect 17509 32181 17543 32215
rect 17543 32181 17552 32215
rect 17500 32172 17552 32181
rect 18512 32172 18564 32224
rect 18788 32172 18840 32224
rect 21272 32215 21324 32224
rect 21272 32181 21281 32215
rect 21281 32181 21315 32215
rect 21315 32181 21324 32215
rect 21272 32172 21324 32181
rect 22376 32351 22428 32360
rect 22376 32317 22385 32351
rect 22385 32317 22419 32351
rect 22419 32317 22428 32351
rect 22376 32308 22428 32317
rect 28448 32385 28457 32419
rect 28457 32385 28491 32419
rect 28491 32385 28500 32419
rect 28448 32376 28500 32385
rect 28816 32419 28868 32428
rect 28816 32385 28825 32419
rect 28825 32385 28859 32419
rect 28859 32385 28868 32419
rect 28816 32376 28868 32385
rect 30104 32444 30156 32496
rect 31668 32444 31720 32496
rect 34520 32444 34572 32496
rect 34612 32444 34664 32496
rect 35164 32487 35216 32496
rect 35164 32453 35173 32487
rect 35173 32453 35207 32487
rect 35207 32453 35216 32487
rect 35164 32444 35216 32453
rect 35808 32444 35860 32496
rect 29644 32376 29696 32428
rect 30196 32419 30248 32428
rect 30196 32385 30205 32419
rect 30205 32385 30239 32419
rect 30239 32385 30248 32419
rect 30196 32376 30248 32385
rect 23020 32240 23072 32292
rect 28264 32308 28316 32360
rect 29736 32308 29788 32360
rect 30380 32376 30432 32428
rect 31208 32376 31260 32428
rect 32864 32376 32916 32428
rect 34888 32419 34940 32428
rect 34888 32385 34897 32419
rect 34897 32385 34931 32419
rect 34931 32385 34940 32419
rect 34888 32376 34940 32385
rect 35256 32419 35308 32428
rect 35256 32385 35265 32419
rect 35265 32385 35299 32419
rect 35299 32385 35308 32419
rect 35256 32376 35308 32385
rect 37832 32419 37884 32428
rect 37832 32385 37841 32419
rect 37841 32385 37875 32419
rect 37875 32385 37884 32419
rect 37832 32376 37884 32385
rect 32588 32308 32640 32360
rect 32772 32351 32824 32360
rect 32772 32317 32781 32351
rect 32781 32317 32815 32351
rect 32815 32317 32824 32351
rect 32772 32308 32824 32317
rect 35624 32308 35676 32360
rect 38108 32351 38160 32360
rect 38108 32317 38117 32351
rect 38117 32317 38151 32351
rect 38151 32317 38160 32351
rect 38108 32308 38160 32317
rect 28172 32240 28224 32292
rect 28724 32240 28776 32292
rect 32312 32240 32364 32292
rect 35716 32240 35768 32292
rect 36084 32240 36136 32292
rect 23296 32172 23348 32224
rect 25688 32172 25740 32224
rect 27160 32215 27212 32224
rect 27160 32181 27169 32215
rect 27169 32181 27203 32215
rect 27203 32181 27212 32215
rect 27160 32172 27212 32181
rect 31392 32172 31444 32224
rect 31576 32172 31628 32224
rect 34152 32215 34204 32224
rect 34152 32181 34161 32215
rect 34161 32181 34195 32215
rect 34195 32181 34204 32215
rect 34152 32172 34204 32181
rect 36176 32172 36228 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 6460 32011 6512 32020
rect 6460 31977 6469 32011
rect 6469 31977 6503 32011
rect 6503 31977 6512 32011
rect 6460 31968 6512 31977
rect 6552 31968 6604 32020
rect 4896 31900 4948 31952
rect 4712 31832 4764 31884
rect 5540 31832 5592 31884
rect 5632 31764 5684 31816
rect 5816 31764 5868 31816
rect 8300 31968 8352 32020
rect 9864 31968 9916 32020
rect 10140 32011 10192 32020
rect 10140 31977 10149 32011
rect 10149 31977 10183 32011
rect 10183 31977 10192 32011
rect 10140 31968 10192 31977
rect 11520 32011 11572 32020
rect 11520 31977 11529 32011
rect 11529 31977 11563 32011
rect 11563 31977 11572 32011
rect 11520 31968 11572 31977
rect 6828 31943 6880 31952
rect 6828 31909 6837 31943
rect 6837 31909 6871 31943
rect 6871 31909 6880 31943
rect 6828 31900 6880 31909
rect 6736 31807 6788 31816
rect 6736 31773 6745 31807
rect 6745 31773 6779 31807
rect 6779 31773 6788 31807
rect 6736 31764 6788 31773
rect 7012 31764 7064 31816
rect 6644 31628 6696 31680
rect 8208 31807 8260 31816
rect 8208 31773 8217 31807
rect 8217 31773 8251 31807
rect 8251 31773 8260 31807
rect 8208 31764 8260 31773
rect 8300 31807 8352 31816
rect 8300 31773 8309 31807
rect 8309 31773 8343 31807
rect 8343 31773 8352 31807
rect 8300 31764 8352 31773
rect 7656 31628 7708 31680
rect 10048 31832 10100 31884
rect 9772 31764 9824 31816
rect 9956 31764 10008 31816
rect 10232 31764 10284 31816
rect 10600 31807 10652 31816
rect 10600 31773 10609 31807
rect 10609 31773 10643 31807
rect 10643 31773 10652 31807
rect 10600 31764 10652 31773
rect 11704 31807 11756 31816
rect 11704 31773 11713 31807
rect 11713 31773 11747 31807
rect 11747 31773 11756 31807
rect 11704 31764 11756 31773
rect 11980 31900 12032 31952
rect 12348 31968 12400 32020
rect 14924 32011 14976 32020
rect 14924 31977 14933 32011
rect 14933 31977 14967 32011
rect 14967 31977 14976 32011
rect 14924 31968 14976 31977
rect 15108 32011 15160 32020
rect 15108 31977 15117 32011
rect 15117 31977 15151 32011
rect 15151 31977 15160 32011
rect 15108 31968 15160 31977
rect 15200 31968 15252 32020
rect 17408 31968 17460 32020
rect 17224 31900 17276 31952
rect 19064 31900 19116 31952
rect 21732 31968 21784 32020
rect 22836 31968 22888 32020
rect 11152 31696 11204 31748
rect 11520 31696 11572 31748
rect 12348 31764 12400 31816
rect 12624 31807 12676 31816
rect 12624 31773 12633 31807
rect 12633 31773 12667 31807
rect 12667 31773 12676 31807
rect 12624 31764 12676 31773
rect 12900 31764 12952 31816
rect 14832 31807 14884 31816
rect 14556 31696 14608 31748
rect 14832 31773 14841 31807
rect 14841 31773 14875 31807
rect 14875 31773 14884 31807
rect 14832 31764 14884 31773
rect 17500 31832 17552 31884
rect 15752 31764 15804 31816
rect 16948 31807 17000 31816
rect 16948 31773 16957 31807
rect 16957 31773 16991 31807
rect 16991 31773 17000 31807
rect 16948 31764 17000 31773
rect 17316 31807 17368 31816
rect 17316 31773 17325 31807
rect 17325 31773 17359 31807
rect 17359 31773 17368 31807
rect 17316 31764 17368 31773
rect 17960 31764 18012 31816
rect 18420 31764 18472 31816
rect 18788 31832 18840 31884
rect 18972 31832 19024 31884
rect 23388 31900 23440 31952
rect 23664 31968 23716 32020
rect 24124 31968 24176 32020
rect 25320 31968 25372 32020
rect 26884 31968 26936 32020
rect 28448 31968 28500 32020
rect 32864 31968 32916 32020
rect 37832 31968 37884 32020
rect 18696 31807 18748 31816
rect 18696 31773 18705 31807
rect 18705 31773 18739 31807
rect 18739 31773 18748 31807
rect 18696 31764 18748 31773
rect 15844 31696 15896 31748
rect 20444 31764 20496 31816
rect 20720 31764 20772 31816
rect 22468 31832 22520 31884
rect 9864 31628 9916 31680
rect 10600 31628 10652 31680
rect 12624 31628 12676 31680
rect 12808 31628 12860 31680
rect 15016 31628 15068 31680
rect 18972 31628 19024 31680
rect 19340 31628 19392 31680
rect 19984 31628 20036 31680
rect 21548 31807 21600 31816
rect 21548 31773 21557 31807
rect 21557 31773 21591 31807
rect 21591 31773 21600 31807
rect 21548 31764 21600 31773
rect 21916 31764 21968 31816
rect 23204 31832 23256 31884
rect 23296 31832 23348 31884
rect 25504 31832 25556 31884
rect 21732 31696 21784 31748
rect 22376 31696 22428 31748
rect 22560 31696 22612 31748
rect 23480 31764 23532 31816
rect 24860 31764 24912 31816
rect 25596 31807 25648 31816
rect 25596 31773 25605 31807
rect 25605 31773 25639 31807
rect 25639 31773 25648 31807
rect 25596 31764 25648 31773
rect 25780 31807 25832 31816
rect 25780 31773 25789 31807
rect 25789 31773 25823 31807
rect 25823 31773 25832 31807
rect 25780 31764 25832 31773
rect 26884 31807 26936 31816
rect 25412 31696 25464 31748
rect 26240 31696 26292 31748
rect 26424 31696 26476 31748
rect 25044 31628 25096 31680
rect 25872 31628 25924 31680
rect 26056 31628 26108 31680
rect 26884 31773 26893 31807
rect 26893 31773 26927 31807
rect 26927 31773 26936 31807
rect 26884 31764 26936 31773
rect 27528 31832 27580 31884
rect 27712 31764 27764 31816
rect 28816 31900 28868 31952
rect 29000 31943 29052 31952
rect 29000 31909 29009 31943
rect 29009 31909 29043 31943
rect 29043 31909 29052 31943
rect 29000 31900 29052 31909
rect 28264 31832 28316 31884
rect 35716 31900 35768 31952
rect 26792 31696 26844 31748
rect 29092 31764 29144 31816
rect 28908 31696 28960 31748
rect 32036 31739 32088 31748
rect 32036 31705 32045 31739
rect 32045 31705 32079 31739
rect 32079 31705 32088 31739
rect 32036 31696 32088 31705
rect 32496 31764 32548 31816
rect 32956 31807 33008 31816
rect 32956 31773 32965 31807
rect 32965 31773 32999 31807
rect 32999 31773 33008 31807
rect 32956 31764 33008 31773
rect 35256 31807 35308 31816
rect 35256 31773 35265 31807
rect 35265 31773 35299 31807
rect 35299 31773 35308 31807
rect 35256 31764 35308 31773
rect 32588 31696 32640 31748
rect 35440 31764 35492 31816
rect 36268 31832 36320 31884
rect 35900 31764 35952 31816
rect 37464 31764 37516 31816
rect 28632 31628 28684 31680
rect 32128 31628 32180 31680
rect 37740 31671 37792 31680
rect 37740 31637 37749 31671
rect 37749 31637 37783 31671
rect 37783 31637 37792 31671
rect 37740 31628 37792 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 11888 31424 11940 31476
rect 12900 31424 12952 31476
rect 5448 31288 5500 31340
rect 5540 31331 5592 31340
rect 5540 31297 5549 31331
rect 5549 31297 5583 31331
rect 5583 31297 5592 31331
rect 5540 31288 5592 31297
rect 6644 31288 6696 31340
rect 7840 31356 7892 31408
rect 9128 31356 9180 31408
rect 13636 31356 13688 31408
rect 7656 31331 7708 31340
rect 7656 31297 7665 31331
rect 7665 31297 7699 31331
rect 7699 31297 7708 31331
rect 7656 31288 7708 31297
rect 10324 31288 10376 31340
rect 10600 31288 10652 31340
rect 11796 31331 11848 31340
rect 11796 31297 11805 31331
rect 11805 31297 11839 31331
rect 11839 31297 11848 31331
rect 11796 31288 11848 31297
rect 8208 31220 8260 31272
rect 9588 31220 9640 31272
rect 7932 31152 7984 31204
rect 11060 31220 11112 31272
rect 12348 31288 12400 31340
rect 12440 31288 12492 31340
rect 12256 31220 12308 31272
rect 12992 31288 13044 31340
rect 14556 31331 14608 31340
rect 14556 31297 14565 31331
rect 14565 31297 14599 31331
rect 14599 31297 14608 31331
rect 14556 31288 14608 31297
rect 15384 31424 15436 31476
rect 17408 31424 17460 31476
rect 18880 31467 18932 31476
rect 18880 31433 18889 31467
rect 18889 31433 18923 31467
rect 18923 31433 18932 31467
rect 18880 31424 18932 31433
rect 16856 31399 16908 31408
rect 16856 31365 16865 31399
rect 16865 31365 16899 31399
rect 16899 31365 16908 31399
rect 16856 31356 16908 31365
rect 16948 31356 17000 31408
rect 19984 31424 20036 31476
rect 22008 31424 22060 31476
rect 23572 31424 23624 31476
rect 25596 31424 25648 31476
rect 27436 31424 27488 31476
rect 27896 31424 27948 31476
rect 28264 31424 28316 31476
rect 30748 31424 30800 31476
rect 16212 31288 16264 31340
rect 19156 31356 19208 31408
rect 19524 31356 19576 31408
rect 18512 31331 18564 31340
rect 11888 31152 11940 31204
rect 13820 31152 13872 31204
rect 15384 31220 15436 31272
rect 15476 31263 15528 31272
rect 15476 31229 15485 31263
rect 15485 31229 15519 31263
rect 15519 31229 15528 31263
rect 17224 31263 17276 31272
rect 15476 31220 15528 31229
rect 17224 31229 17233 31263
rect 17233 31229 17267 31263
rect 17267 31229 17276 31263
rect 17224 31220 17276 31229
rect 17408 31220 17460 31272
rect 18512 31297 18521 31331
rect 18521 31297 18555 31331
rect 18555 31297 18564 31331
rect 18512 31288 18564 31297
rect 18788 31288 18840 31340
rect 18972 31288 19024 31340
rect 20260 31288 20312 31340
rect 22376 31356 22428 31408
rect 21456 31331 21508 31340
rect 21456 31297 21465 31331
rect 21465 31297 21499 31331
rect 21499 31297 21508 31331
rect 21456 31288 21508 31297
rect 22284 31331 22336 31340
rect 22284 31297 22293 31331
rect 22293 31297 22327 31331
rect 22327 31297 22336 31331
rect 22284 31288 22336 31297
rect 23664 31331 23716 31340
rect 23664 31297 23673 31331
rect 23673 31297 23707 31331
rect 23707 31297 23716 31331
rect 23664 31288 23716 31297
rect 23756 31288 23808 31340
rect 5540 31084 5592 31136
rect 6092 31084 6144 31136
rect 9772 31084 9824 31136
rect 10508 31084 10560 31136
rect 11704 31084 11756 31136
rect 15844 31152 15896 31204
rect 17592 31152 17644 31204
rect 19892 31263 19944 31272
rect 19892 31229 19901 31263
rect 19901 31229 19935 31263
rect 19935 31229 19944 31263
rect 19892 31220 19944 31229
rect 21548 31220 21600 31272
rect 25412 31288 25464 31340
rect 25596 31288 25648 31340
rect 20168 31152 20220 31204
rect 23480 31152 23532 31204
rect 24308 31152 24360 31204
rect 25228 31220 25280 31272
rect 25872 31331 25924 31340
rect 25872 31297 25881 31331
rect 25881 31297 25915 31331
rect 25915 31297 25924 31331
rect 25872 31288 25924 31297
rect 29000 31356 29052 31408
rect 30564 31356 30616 31408
rect 32036 31424 32088 31476
rect 32956 31424 33008 31476
rect 35256 31424 35308 31476
rect 35348 31424 35400 31476
rect 35624 31424 35676 31476
rect 37464 31467 37516 31476
rect 37464 31433 37473 31467
rect 37473 31433 37507 31467
rect 37507 31433 37516 31467
rect 37464 31424 37516 31433
rect 37832 31424 37884 31476
rect 25964 31152 26016 31204
rect 27252 31288 27304 31340
rect 27436 31331 27488 31340
rect 27436 31297 27445 31331
rect 27445 31297 27479 31331
rect 27479 31297 27488 31331
rect 27436 31288 27488 31297
rect 26884 31220 26936 31272
rect 28632 31288 28684 31340
rect 29184 31288 29236 31340
rect 30656 31331 30708 31340
rect 27620 31220 27672 31272
rect 27896 31220 27948 31272
rect 28908 31220 28960 31272
rect 26424 31152 26476 31204
rect 30656 31297 30665 31331
rect 30665 31297 30699 31331
rect 30699 31297 30708 31331
rect 30656 31288 30708 31297
rect 30748 31331 30800 31340
rect 30748 31297 30758 31331
rect 30758 31297 30792 31331
rect 30792 31297 30800 31331
rect 30932 31331 30984 31340
rect 30748 31288 30800 31297
rect 30932 31297 30941 31331
rect 30941 31297 30975 31331
rect 30975 31297 30984 31331
rect 30932 31288 30984 31297
rect 31576 31288 31628 31340
rect 32128 31356 32180 31408
rect 34612 31356 34664 31408
rect 35532 31356 35584 31408
rect 34152 31288 34204 31340
rect 34520 31331 34572 31340
rect 34520 31297 34529 31331
rect 34529 31297 34563 31331
rect 34563 31297 34572 31331
rect 34520 31288 34572 31297
rect 34888 31331 34940 31340
rect 34888 31297 34897 31331
rect 34897 31297 34931 31331
rect 34931 31297 34940 31331
rect 34888 31288 34940 31297
rect 35440 31288 35492 31340
rect 37740 31288 37792 31340
rect 34612 31220 34664 31272
rect 38016 31263 38068 31272
rect 38016 31229 38025 31263
rect 38025 31229 38059 31263
rect 38059 31229 38068 31263
rect 38016 31220 38068 31229
rect 17500 31084 17552 31136
rect 18788 31084 18840 31136
rect 20904 31084 20956 31136
rect 22560 31084 22612 31136
rect 25412 31127 25464 31136
rect 25412 31093 25421 31127
rect 25421 31093 25455 31127
rect 25455 31093 25464 31127
rect 25412 31084 25464 31093
rect 26056 31084 26108 31136
rect 35992 31152 36044 31204
rect 32496 31127 32548 31136
rect 32496 31093 32505 31127
rect 32505 31093 32539 31127
rect 32539 31093 32548 31127
rect 32496 31084 32548 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 6552 30923 6604 30932
rect 6552 30889 6561 30923
rect 6561 30889 6595 30923
rect 6595 30889 6604 30923
rect 6552 30880 6604 30889
rect 7012 30923 7064 30932
rect 7012 30889 7021 30923
rect 7021 30889 7055 30923
rect 7055 30889 7064 30923
rect 7012 30880 7064 30889
rect 7932 30923 7984 30932
rect 7932 30889 7941 30923
rect 7941 30889 7975 30923
rect 7975 30889 7984 30923
rect 7932 30880 7984 30889
rect 9404 30880 9456 30932
rect 10232 30880 10284 30932
rect 12072 30880 12124 30932
rect 12992 30880 13044 30932
rect 14188 30880 14240 30932
rect 15016 30880 15068 30932
rect 6920 30812 6972 30864
rect 7380 30812 7432 30864
rect 6644 30787 6696 30796
rect 6644 30753 6653 30787
rect 6653 30753 6687 30787
rect 6687 30753 6696 30787
rect 6644 30744 6696 30753
rect 7196 30744 7248 30796
rect 8208 30744 8260 30796
rect 4896 30651 4948 30660
rect 4896 30617 4905 30651
rect 4905 30617 4939 30651
rect 4939 30617 4948 30651
rect 4896 30608 4948 30617
rect 5264 30651 5316 30660
rect 5264 30617 5273 30651
rect 5273 30617 5307 30651
rect 5307 30617 5316 30651
rect 5264 30608 5316 30617
rect 6092 30651 6144 30660
rect 6092 30617 6101 30651
rect 6101 30617 6135 30651
rect 6135 30617 6144 30651
rect 6092 30608 6144 30617
rect 8116 30719 8168 30728
rect 8116 30685 8125 30719
rect 8125 30685 8159 30719
rect 8159 30685 8168 30719
rect 8116 30676 8168 30685
rect 7564 30608 7616 30660
rect 7932 30608 7984 30660
rect 9220 30676 9272 30728
rect 10600 30812 10652 30864
rect 12440 30812 12492 30864
rect 11060 30744 11112 30796
rect 11704 30719 11756 30728
rect 11704 30685 11713 30719
rect 11713 30685 11747 30719
rect 11747 30685 11756 30719
rect 11704 30676 11756 30685
rect 11980 30676 12032 30728
rect 12348 30676 12400 30728
rect 13728 30744 13780 30796
rect 13360 30719 13412 30728
rect 13360 30685 13369 30719
rect 13369 30685 13403 30719
rect 13403 30685 13412 30719
rect 13360 30676 13412 30685
rect 12808 30608 12860 30660
rect 15016 30676 15068 30728
rect 15476 30812 15528 30864
rect 19340 30880 19392 30932
rect 19708 30923 19760 30932
rect 19708 30889 19717 30923
rect 19717 30889 19751 30923
rect 19751 30889 19760 30923
rect 19708 30880 19760 30889
rect 20444 30923 20496 30932
rect 20444 30889 20453 30923
rect 20453 30889 20487 30923
rect 20487 30889 20496 30923
rect 20444 30880 20496 30889
rect 20904 30880 20956 30932
rect 22008 30880 22060 30932
rect 22284 30880 22336 30932
rect 25044 30880 25096 30932
rect 29644 30880 29696 30932
rect 31116 30880 31168 30932
rect 34244 30880 34296 30932
rect 13544 30608 13596 30660
rect 15476 30719 15528 30728
rect 15476 30685 15485 30719
rect 15485 30685 15519 30719
rect 15519 30685 15528 30719
rect 15476 30676 15528 30685
rect 15844 30676 15896 30728
rect 16580 30719 16632 30728
rect 16580 30685 16589 30719
rect 16589 30685 16623 30719
rect 16623 30685 16632 30719
rect 16580 30676 16632 30685
rect 17224 30676 17276 30728
rect 17500 30608 17552 30660
rect 17592 30651 17644 30660
rect 17592 30617 17601 30651
rect 17601 30617 17635 30651
rect 17635 30617 17644 30651
rect 18696 30744 18748 30796
rect 25412 30812 25464 30864
rect 25872 30812 25924 30864
rect 20444 30744 20496 30796
rect 21456 30744 21508 30796
rect 19984 30676 20036 30728
rect 20536 30676 20588 30728
rect 22284 30719 22336 30728
rect 22284 30685 22293 30719
rect 22293 30685 22327 30719
rect 22327 30685 22336 30719
rect 22284 30676 22336 30685
rect 23020 30744 23072 30796
rect 23204 30744 23256 30796
rect 27252 30812 27304 30864
rect 28908 30855 28960 30864
rect 22744 30676 22796 30728
rect 23480 30676 23532 30728
rect 23572 30719 23624 30728
rect 23572 30685 23581 30719
rect 23581 30685 23615 30719
rect 23615 30685 23624 30719
rect 23572 30676 23624 30685
rect 23756 30676 23808 30728
rect 24860 30676 24912 30728
rect 25136 30719 25188 30728
rect 25136 30685 25145 30719
rect 25145 30685 25179 30719
rect 25179 30685 25188 30719
rect 25136 30676 25188 30685
rect 17592 30608 17644 30617
rect 9864 30540 9916 30592
rect 11152 30540 11204 30592
rect 12532 30540 12584 30592
rect 15016 30540 15068 30592
rect 15200 30540 15252 30592
rect 17868 30540 17920 30592
rect 18052 30583 18104 30592
rect 18052 30549 18061 30583
rect 18061 30549 18095 30583
rect 18095 30549 18104 30583
rect 18052 30540 18104 30549
rect 18144 30540 18196 30592
rect 22928 30608 22980 30660
rect 20904 30540 20956 30592
rect 23756 30583 23808 30592
rect 23756 30549 23765 30583
rect 23765 30549 23799 30583
rect 23799 30549 23808 30583
rect 23756 30540 23808 30549
rect 25504 30676 25556 30728
rect 25964 30676 26016 30728
rect 25688 30608 25740 30660
rect 27436 30744 27488 30796
rect 27896 30744 27948 30796
rect 28908 30821 28917 30855
rect 28917 30821 28951 30855
rect 28951 30821 28960 30855
rect 28908 30812 28960 30821
rect 32496 30812 32548 30864
rect 26516 30540 26568 30592
rect 27436 30583 27488 30592
rect 27436 30549 27445 30583
rect 27445 30549 27479 30583
rect 27479 30549 27488 30583
rect 27436 30540 27488 30549
rect 27712 30676 27764 30728
rect 29000 30676 29052 30728
rect 30748 30719 30800 30728
rect 30748 30685 30757 30719
rect 30757 30685 30791 30719
rect 30791 30685 30800 30719
rect 30748 30676 30800 30685
rect 30840 30719 30892 30728
rect 30840 30685 30850 30719
rect 30850 30685 30884 30719
rect 30884 30685 30892 30719
rect 34060 30744 34112 30796
rect 34612 30744 34664 30796
rect 30840 30676 30892 30685
rect 31576 30676 31628 30728
rect 32128 30676 32180 30728
rect 32588 30676 32640 30728
rect 35532 30744 35584 30796
rect 27988 30608 28040 30660
rect 30196 30608 30248 30660
rect 30932 30608 30984 30660
rect 28172 30540 28224 30592
rect 28632 30540 28684 30592
rect 31116 30651 31168 30660
rect 31116 30617 31125 30651
rect 31125 30617 31159 30651
rect 31159 30617 31168 30651
rect 31116 30608 31168 30617
rect 31392 30540 31444 30592
rect 31852 30608 31904 30660
rect 35440 30719 35492 30728
rect 35440 30685 35449 30719
rect 35449 30685 35483 30719
rect 35483 30685 35492 30719
rect 36728 30719 36780 30728
rect 35440 30676 35492 30685
rect 36728 30685 36737 30719
rect 36737 30685 36771 30719
rect 36771 30685 36780 30719
rect 36728 30676 36780 30685
rect 34796 30608 34848 30660
rect 37004 30651 37056 30660
rect 37004 30617 37013 30651
rect 37013 30617 37047 30651
rect 37047 30617 37056 30651
rect 37004 30608 37056 30617
rect 37280 30608 37332 30660
rect 35532 30540 35584 30592
rect 35808 30540 35860 30592
rect 38016 30583 38068 30592
rect 38016 30549 38025 30583
rect 38025 30549 38059 30583
rect 38059 30549 38068 30583
rect 38016 30540 38068 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4896 30336 4948 30388
rect 6552 30336 6604 30388
rect 7472 30336 7524 30388
rect 7932 30336 7984 30388
rect 9680 30336 9732 30388
rect 10324 30336 10376 30388
rect 11796 30336 11848 30388
rect 2780 30200 2832 30252
rect 9588 30268 9640 30320
rect 3976 30200 4028 30252
rect 5540 30200 5592 30252
rect 6368 30200 6420 30252
rect 6920 30200 6972 30252
rect 8668 30243 8720 30252
rect 8668 30209 8677 30243
rect 8677 30209 8711 30243
rect 8711 30209 8720 30243
rect 8668 30200 8720 30209
rect 9036 30243 9088 30252
rect 9036 30209 9045 30243
rect 9045 30209 9079 30243
rect 9079 30209 9088 30243
rect 9036 30200 9088 30209
rect 9312 30200 9364 30252
rect 6276 30132 6328 30184
rect 6552 30175 6604 30184
rect 6552 30141 6561 30175
rect 6561 30141 6595 30175
rect 6595 30141 6604 30175
rect 6552 30132 6604 30141
rect 7104 30132 7156 30184
rect 8116 30132 8168 30184
rect 11980 30268 12032 30320
rect 10048 30200 10100 30252
rect 10140 30243 10192 30252
rect 10140 30209 10149 30243
rect 10149 30209 10183 30243
rect 10183 30209 10192 30243
rect 10140 30200 10192 30209
rect 11980 30132 12032 30184
rect 13912 30200 13964 30252
rect 14188 30268 14240 30320
rect 14464 30336 14516 30388
rect 15752 30336 15804 30388
rect 16580 30336 16632 30388
rect 23204 30336 23256 30388
rect 23572 30336 23624 30388
rect 26240 30336 26292 30388
rect 30656 30336 30708 30388
rect 30840 30336 30892 30388
rect 18144 30268 18196 30320
rect 20260 30311 20312 30320
rect 20260 30277 20269 30311
rect 20269 30277 20303 30311
rect 20303 30277 20312 30311
rect 20260 30268 20312 30277
rect 14464 30200 14516 30252
rect 13176 30175 13228 30184
rect 13176 30141 13185 30175
rect 13185 30141 13219 30175
rect 13219 30141 13228 30175
rect 13176 30132 13228 30141
rect 13268 30132 13320 30184
rect 15200 30243 15252 30252
rect 15200 30209 15209 30243
rect 15209 30209 15243 30243
rect 15243 30209 15252 30243
rect 15200 30200 15252 30209
rect 16028 30200 16080 30252
rect 18052 30200 18104 30252
rect 15752 30175 15804 30184
rect 5448 30064 5500 30116
rect 4620 29996 4672 30048
rect 12808 30064 12860 30116
rect 8208 30039 8260 30048
rect 8208 30005 8217 30039
rect 8217 30005 8251 30039
rect 8251 30005 8260 30039
rect 8208 29996 8260 30005
rect 13820 30039 13872 30048
rect 13820 30005 13829 30039
rect 13829 30005 13863 30039
rect 13863 30005 13872 30039
rect 13820 29996 13872 30005
rect 14648 30064 14700 30116
rect 15752 30141 15761 30175
rect 15761 30141 15795 30175
rect 15795 30141 15804 30175
rect 15752 30132 15804 30141
rect 17500 30175 17552 30184
rect 17500 30141 17509 30175
rect 17509 30141 17543 30175
rect 17543 30141 17552 30175
rect 17500 30132 17552 30141
rect 16304 30064 16356 30116
rect 16856 30064 16908 30116
rect 17960 30132 18012 30184
rect 18604 30200 18656 30252
rect 19156 30200 19208 30252
rect 19984 30200 20036 30252
rect 20444 30243 20496 30252
rect 20444 30209 20453 30243
rect 20453 30209 20487 30243
rect 20487 30209 20496 30243
rect 20444 30200 20496 30209
rect 22100 30200 22152 30252
rect 22744 30200 22796 30252
rect 22836 30200 22888 30252
rect 23020 30175 23072 30184
rect 17684 30064 17736 30116
rect 23020 30141 23029 30175
rect 23029 30141 23063 30175
rect 23063 30141 23072 30175
rect 23020 30132 23072 30141
rect 23204 30175 23256 30184
rect 23204 30141 23213 30175
rect 23213 30141 23247 30175
rect 23247 30141 23256 30175
rect 23204 30132 23256 30141
rect 23664 30268 23716 30320
rect 24768 30268 24820 30320
rect 24216 30200 24268 30252
rect 24860 30200 24912 30252
rect 25780 30200 25832 30252
rect 26240 30200 26292 30252
rect 26516 30243 26568 30252
rect 26516 30209 26525 30243
rect 26525 30209 26559 30243
rect 26559 30209 26568 30243
rect 26516 30200 26568 30209
rect 25228 30132 25280 30184
rect 14924 29996 14976 30048
rect 15568 29996 15620 30048
rect 15660 30039 15712 30048
rect 15660 30005 15669 30039
rect 15669 30005 15703 30039
rect 15703 30005 15712 30039
rect 15660 29996 15712 30005
rect 15936 29996 15988 30048
rect 17408 30039 17460 30048
rect 17408 30005 17417 30039
rect 17417 30005 17451 30039
rect 17451 30005 17460 30039
rect 17408 29996 17460 30005
rect 18236 30039 18288 30048
rect 18236 30005 18245 30039
rect 18245 30005 18279 30039
rect 18279 30005 18288 30039
rect 18236 29996 18288 30005
rect 20628 30039 20680 30048
rect 20628 30005 20637 30039
rect 20637 30005 20671 30039
rect 20671 30005 20680 30039
rect 20628 29996 20680 30005
rect 22560 30064 22612 30116
rect 22928 30107 22980 30116
rect 22928 30073 22937 30107
rect 22937 30073 22971 30107
rect 22971 30073 22980 30107
rect 22928 30064 22980 30073
rect 23296 30064 23348 30116
rect 27712 30175 27764 30184
rect 27712 30141 27721 30175
rect 27721 30141 27755 30175
rect 27755 30141 27764 30175
rect 27712 30132 27764 30141
rect 28172 30268 28224 30320
rect 28356 30243 28408 30252
rect 28356 30209 28365 30243
rect 28365 30209 28399 30243
rect 28399 30209 28408 30243
rect 28356 30200 28408 30209
rect 28908 30200 28960 30252
rect 29644 30200 29696 30252
rect 31024 30268 31076 30320
rect 31392 30311 31444 30320
rect 31392 30277 31401 30311
rect 31401 30277 31435 30311
rect 31435 30277 31444 30311
rect 34060 30311 34112 30320
rect 31392 30268 31444 30277
rect 34060 30277 34094 30311
rect 34094 30277 34112 30311
rect 34060 30268 34112 30277
rect 30012 30243 30064 30252
rect 30012 30209 30021 30243
rect 30021 30209 30055 30243
rect 30055 30209 30064 30243
rect 30012 30200 30064 30209
rect 28724 30175 28776 30184
rect 28724 30141 28733 30175
rect 28733 30141 28767 30175
rect 28767 30141 28776 30175
rect 28724 30132 28776 30141
rect 29368 30064 29420 30116
rect 30288 30200 30340 30252
rect 30472 30200 30524 30252
rect 31116 30243 31168 30252
rect 31116 30209 31125 30243
rect 31125 30209 31159 30243
rect 31159 30209 31168 30243
rect 31116 30200 31168 30209
rect 31300 30243 31352 30252
rect 31300 30209 31307 30243
rect 31307 30209 31352 30243
rect 31300 30200 31352 30209
rect 31024 30132 31076 30184
rect 31576 30243 31628 30252
rect 31576 30209 31590 30243
rect 31590 30209 31624 30243
rect 31624 30209 31628 30243
rect 31576 30200 31628 30209
rect 32220 30132 32272 30184
rect 32772 30132 32824 30184
rect 30380 30064 30432 30116
rect 31852 30064 31904 30116
rect 35900 30336 35952 30388
rect 36176 30311 36228 30320
rect 36176 30277 36185 30311
rect 36185 30277 36219 30311
rect 36219 30277 36228 30311
rect 36176 30268 36228 30277
rect 37832 30379 37884 30388
rect 37832 30345 37841 30379
rect 37841 30345 37875 30379
rect 37875 30345 37884 30379
rect 37832 30336 37884 30345
rect 36728 30268 36780 30320
rect 35808 30243 35860 30252
rect 35808 30209 35817 30243
rect 35817 30209 35851 30243
rect 35851 30209 35860 30243
rect 35808 30200 35860 30209
rect 35900 30243 35952 30252
rect 35900 30209 35910 30243
rect 35910 30209 35944 30243
rect 35944 30209 35952 30243
rect 35900 30200 35952 30209
rect 36084 30243 36136 30252
rect 36084 30209 36093 30243
rect 36093 30209 36127 30243
rect 36127 30209 36136 30243
rect 36084 30200 36136 30209
rect 36268 30243 36320 30252
rect 36268 30209 36282 30243
rect 36282 30209 36316 30243
rect 36316 30209 36320 30243
rect 36268 30200 36320 30209
rect 38016 30175 38068 30184
rect 38016 30141 38025 30175
rect 38025 30141 38059 30175
rect 38059 30141 38068 30175
rect 38016 30132 38068 30141
rect 36084 30064 36136 30116
rect 24308 29996 24360 30048
rect 24676 29996 24728 30048
rect 25504 30039 25556 30048
rect 25504 30005 25513 30039
rect 25513 30005 25547 30039
rect 25547 30005 25556 30039
rect 25504 29996 25556 30005
rect 28632 30039 28684 30048
rect 28632 30005 28641 30039
rect 28641 30005 28675 30039
rect 28675 30005 28684 30039
rect 28632 29996 28684 30005
rect 29460 29996 29512 30048
rect 31392 29996 31444 30048
rect 31576 29996 31628 30048
rect 32404 29996 32456 30048
rect 37464 30039 37516 30048
rect 37464 30005 37473 30039
rect 37473 30005 37507 30039
rect 37507 30005 37516 30039
rect 37464 29996 37516 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 3976 29835 4028 29844
rect 3976 29801 3985 29835
rect 3985 29801 4019 29835
rect 4019 29801 4028 29835
rect 3976 29792 4028 29801
rect 6368 29792 6420 29844
rect 8760 29792 8812 29844
rect 9036 29792 9088 29844
rect 10508 29792 10560 29844
rect 11796 29835 11848 29844
rect 5264 29724 5316 29776
rect 4160 29656 4212 29708
rect 5080 29656 5132 29708
rect 6276 29724 6328 29776
rect 6552 29724 6604 29776
rect 11796 29801 11805 29835
rect 11805 29801 11839 29835
rect 11839 29801 11848 29835
rect 11796 29792 11848 29801
rect 12256 29792 12308 29844
rect 5632 29699 5684 29708
rect 4620 29588 4672 29640
rect 5632 29665 5641 29699
rect 5641 29665 5675 29699
rect 5675 29665 5684 29699
rect 5632 29656 5684 29665
rect 6000 29656 6052 29708
rect 5356 29631 5408 29640
rect 5356 29597 5365 29631
rect 5365 29597 5399 29631
rect 5399 29597 5408 29631
rect 5356 29588 5408 29597
rect 5448 29588 5500 29640
rect 6736 29656 6788 29708
rect 5264 29520 5316 29572
rect 6644 29588 6696 29640
rect 7012 29631 7064 29640
rect 7012 29597 7021 29631
rect 7021 29597 7055 29631
rect 7055 29597 7064 29631
rect 7012 29588 7064 29597
rect 7104 29588 7156 29640
rect 7656 29656 7708 29708
rect 12072 29724 12124 29776
rect 15476 29792 15528 29844
rect 17776 29835 17828 29844
rect 6368 29520 6420 29572
rect 8116 29588 8168 29640
rect 7840 29520 7892 29572
rect 9220 29588 9272 29640
rect 9956 29588 10008 29640
rect 11980 29588 12032 29640
rect 12532 29631 12584 29640
rect 12532 29597 12541 29631
rect 12541 29597 12575 29631
rect 12575 29597 12584 29631
rect 14464 29724 14516 29776
rect 15660 29724 15712 29776
rect 17776 29801 17785 29835
rect 17785 29801 17819 29835
rect 17819 29801 17828 29835
rect 17776 29792 17828 29801
rect 22100 29792 22152 29844
rect 22192 29792 22244 29844
rect 23388 29835 23440 29844
rect 23388 29801 23397 29835
rect 23397 29801 23431 29835
rect 23431 29801 23440 29835
rect 23388 29792 23440 29801
rect 26056 29792 26108 29844
rect 26424 29792 26476 29844
rect 26516 29792 26568 29844
rect 20720 29724 20772 29776
rect 22652 29724 22704 29776
rect 28356 29724 28408 29776
rect 30748 29792 30800 29844
rect 30656 29724 30708 29776
rect 14280 29656 14332 29708
rect 15384 29656 15436 29708
rect 18236 29656 18288 29708
rect 19984 29656 20036 29708
rect 12532 29588 12584 29597
rect 11704 29520 11756 29572
rect 13360 29588 13412 29640
rect 13912 29588 13964 29640
rect 15752 29588 15804 29640
rect 16488 29588 16540 29640
rect 13176 29520 13228 29572
rect 16028 29520 16080 29572
rect 16856 29588 16908 29640
rect 17776 29588 17828 29640
rect 20260 29588 20312 29640
rect 20628 29631 20680 29640
rect 20628 29597 20637 29631
rect 20637 29597 20671 29631
rect 20671 29597 20680 29631
rect 20628 29588 20680 29597
rect 21364 29656 21416 29708
rect 22008 29656 22060 29708
rect 21180 29631 21232 29640
rect 21180 29597 21189 29631
rect 21189 29597 21223 29631
rect 21223 29597 21232 29631
rect 21180 29588 21232 29597
rect 24124 29656 24176 29708
rect 22560 29588 22612 29640
rect 23020 29588 23072 29640
rect 23388 29588 23440 29640
rect 23664 29588 23716 29640
rect 17316 29563 17368 29572
rect 17316 29529 17325 29563
rect 17325 29529 17359 29563
rect 17359 29529 17368 29563
rect 17316 29520 17368 29529
rect 18328 29520 18380 29572
rect 19248 29520 19300 29572
rect 20536 29520 20588 29572
rect 27712 29656 27764 29708
rect 25044 29588 25096 29640
rect 25504 29588 25556 29640
rect 26884 29631 26936 29640
rect 26884 29597 26893 29631
rect 26893 29597 26927 29631
rect 26927 29597 26936 29631
rect 26884 29588 26936 29597
rect 27528 29588 27580 29640
rect 29644 29588 29696 29640
rect 30012 29631 30064 29640
rect 30012 29597 30019 29631
rect 30019 29597 30064 29631
rect 30012 29588 30064 29597
rect 30104 29631 30156 29640
rect 30104 29597 30113 29631
rect 30113 29597 30147 29631
rect 30147 29597 30156 29631
rect 30104 29588 30156 29597
rect 30380 29588 30432 29640
rect 32220 29656 32272 29708
rect 32588 29724 32640 29776
rect 32404 29631 32456 29640
rect 3332 29495 3384 29504
rect 3332 29461 3341 29495
rect 3341 29461 3375 29495
rect 3375 29461 3384 29495
rect 3332 29452 3384 29461
rect 6184 29495 6236 29504
rect 6184 29461 6193 29495
rect 6193 29461 6227 29495
rect 6227 29461 6236 29495
rect 6184 29452 6236 29461
rect 6828 29452 6880 29504
rect 7288 29495 7340 29504
rect 7288 29461 7297 29495
rect 7297 29461 7331 29495
rect 7331 29461 7340 29495
rect 7288 29452 7340 29461
rect 8668 29452 8720 29504
rect 11980 29452 12032 29504
rect 15936 29452 15988 29504
rect 16212 29452 16264 29504
rect 16764 29452 16816 29504
rect 18972 29452 19024 29504
rect 19156 29452 19208 29504
rect 19432 29452 19484 29504
rect 20720 29452 20772 29504
rect 24676 29495 24728 29504
rect 24676 29461 24685 29495
rect 24685 29461 24719 29495
rect 24719 29461 24728 29495
rect 24676 29452 24728 29461
rect 24768 29452 24820 29504
rect 27896 29520 27948 29572
rect 29552 29520 29604 29572
rect 32404 29597 32413 29631
rect 32413 29597 32447 29631
rect 32447 29597 32456 29631
rect 32404 29588 32456 29597
rect 32496 29588 32548 29640
rect 34796 29588 34848 29640
rect 37832 29792 37884 29844
rect 35440 29656 35492 29708
rect 35532 29631 35584 29640
rect 35532 29597 35541 29631
rect 35541 29597 35575 29631
rect 35575 29597 35584 29631
rect 35532 29588 35584 29597
rect 36360 29656 36412 29708
rect 36820 29699 36872 29708
rect 36820 29665 36829 29699
rect 36829 29665 36863 29699
rect 36863 29665 36872 29699
rect 36820 29656 36872 29665
rect 37464 29588 37516 29640
rect 31024 29563 31076 29572
rect 31024 29529 31033 29563
rect 31033 29529 31067 29563
rect 31067 29529 31076 29563
rect 31024 29520 31076 29529
rect 35440 29563 35492 29572
rect 35440 29529 35449 29563
rect 35449 29529 35483 29563
rect 35483 29529 35492 29563
rect 35440 29520 35492 29529
rect 25964 29495 26016 29504
rect 25964 29461 25989 29495
rect 25989 29461 26016 29495
rect 25964 29452 26016 29461
rect 26608 29452 26660 29504
rect 30656 29452 30708 29504
rect 31760 29452 31812 29504
rect 32772 29452 32824 29504
rect 33232 29495 33284 29504
rect 33232 29461 33241 29495
rect 33241 29461 33275 29495
rect 33275 29461 33284 29495
rect 33232 29452 33284 29461
rect 35716 29452 35768 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 5172 29248 5224 29300
rect 3332 29180 3384 29232
rect 4804 29180 4856 29232
rect 5448 29180 5500 29232
rect 7012 29180 7064 29232
rect 7472 29180 7524 29232
rect 10140 29248 10192 29300
rect 11796 29291 11848 29300
rect 11796 29257 11805 29291
rect 11805 29257 11839 29291
rect 11839 29257 11848 29291
rect 11796 29248 11848 29257
rect 15660 29248 15712 29300
rect 17868 29248 17920 29300
rect 16212 29180 16264 29232
rect 4068 29155 4120 29164
rect 4068 29121 4077 29155
rect 4077 29121 4111 29155
rect 4111 29121 4120 29155
rect 4068 29112 4120 29121
rect 4896 29112 4948 29164
rect 5264 29155 5316 29164
rect 5264 29121 5273 29155
rect 5273 29121 5307 29155
rect 5307 29121 5316 29155
rect 5264 29112 5316 29121
rect 7564 29112 7616 29164
rect 8760 29112 8812 29164
rect 9588 29112 9640 29164
rect 9864 29112 9916 29164
rect 10232 29112 10284 29164
rect 11520 29112 11572 29164
rect 11612 29112 11664 29164
rect 11888 29155 11940 29164
rect 11888 29121 11897 29155
rect 11897 29121 11931 29155
rect 11931 29121 11940 29155
rect 11888 29112 11940 29121
rect 12808 29155 12860 29164
rect 12808 29121 12817 29155
rect 12817 29121 12851 29155
rect 12851 29121 12860 29155
rect 12808 29112 12860 29121
rect 13636 29155 13688 29164
rect 13636 29121 13645 29155
rect 13645 29121 13679 29155
rect 13679 29121 13688 29155
rect 13636 29112 13688 29121
rect 16948 29112 17000 29164
rect 19432 29248 19484 29300
rect 22284 29248 22336 29300
rect 22928 29248 22980 29300
rect 23388 29291 23440 29300
rect 23388 29257 23397 29291
rect 23397 29257 23431 29291
rect 23431 29257 23440 29291
rect 23388 29248 23440 29257
rect 23572 29248 23624 29300
rect 24032 29248 24084 29300
rect 24952 29291 25004 29300
rect 24952 29257 24961 29291
rect 24961 29257 24995 29291
rect 24995 29257 25004 29291
rect 24952 29248 25004 29257
rect 5356 29044 5408 29096
rect 9220 29044 9272 29096
rect 9772 29044 9824 29096
rect 10140 29087 10192 29096
rect 10140 29053 10149 29087
rect 10149 29053 10183 29087
rect 10183 29053 10192 29087
rect 10140 29044 10192 29053
rect 4620 29019 4672 29028
rect 4620 28985 4629 29019
rect 4629 28985 4663 29019
rect 4663 28985 4672 29019
rect 4620 28976 4672 28985
rect 4896 28976 4948 29028
rect 7104 28976 7156 29028
rect 11152 28976 11204 29028
rect 14188 29044 14240 29096
rect 14924 29044 14976 29096
rect 13084 28976 13136 29028
rect 14648 28976 14700 29028
rect 16304 29087 16356 29096
rect 16304 29053 16313 29087
rect 16313 29053 16347 29087
rect 16347 29053 16356 29087
rect 16304 29044 16356 29053
rect 16488 29044 16540 29096
rect 21916 29180 21968 29232
rect 18144 29112 18196 29164
rect 17408 29087 17460 29096
rect 17408 29053 17417 29087
rect 17417 29053 17451 29087
rect 17451 29053 17460 29087
rect 17408 29044 17460 29053
rect 18512 29087 18564 29096
rect 18512 29053 18521 29087
rect 18521 29053 18555 29087
rect 18555 29053 18564 29087
rect 18512 29044 18564 29053
rect 18788 29087 18840 29096
rect 18788 29053 18797 29087
rect 18797 29053 18831 29087
rect 18831 29053 18840 29087
rect 18788 29044 18840 29053
rect 19248 29112 19300 29164
rect 19432 29112 19484 29164
rect 20260 29155 20312 29164
rect 20260 29121 20269 29155
rect 20269 29121 20303 29155
rect 20303 29121 20312 29155
rect 20260 29112 20312 29121
rect 20720 29155 20772 29164
rect 19616 29044 19668 29096
rect 19984 29044 20036 29096
rect 20720 29121 20729 29155
rect 20729 29121 20763 29155
rect 20763 29121 20772 29155
rect 20720 29112 20772 29121
rect 22008 29112 22060 29164
rect 23388 29112 23440 29164
rect 23572 29155 23624 29164
rect 23572 29121 23581 29155
rect 23581 29121 23615 29155
rect 23615 29121 23624 29155
rect 23572 29112 23624 29121
rect 23756 29155 23808 29164
rect 23756 29121 23765 29155
rect 23765 29121 23799 29155
rect 23799 29121 23808 29155
rect 23756 29112 23808 29121
rect 24768 29112 24820 29164
rect 25964 29248 26016 29300
rect 25228 29180 25280 29232
rect 26884 29180 26936 29232
rect 27712 29223 27764 29232
rect 27712 29189 27721 29223
rect 27721 29189 27755 29223
rect 27755 29189 27764 29223
rect 27712 29180 27764 29189
rect 25412 29155 25464 29164
rect 25412 29121 25421 29155
rect 25421 29121 25455 29155
rect 25455 29121 25464 29155
rect 25964 29155 26016 29164
rect 25412 29112 25464 29121
rect 25964 29121 25973 29155
rect 25973 29121 26007 29155
rect 26007 29121 26016 29155
rect 25964 29112 26016 29121
rect 21456 29044 21508 29096
rect 22652 29044 22704 29096
rect 23664 29087 23716 29096
rect 23664 29053 23673 29087
rect 23673 29053 23707 29087
rect 23707 29053 23716 29087
rect 23664 29044 23716 29053
rect 19064 28976 19116 29028
rect 20260 28976 20312 29028
rect 22560 28976 22612 29028
rect 23204 28976 23256 29028
rect 3976 28908 4028 28960
rect 4160 28908 4212 28960
rect 4712 28908 4764 28960
rect 6736 28908 6788 28960
rect 9128 28908 9180 28960
rect 9220 28908 9272 28960
rect 12440 28908 12492 28960
rect 15844 28908 15896 28960
rect 16304 28908 16356 28960
rect 19340 28908 19392 28960
rect 20812 28908 20864 28960
rect 21732 28908 21784 28960
rect 22284 28908 22336 28960
rect 23296 28908 23348 28960
rect 25228 29087 25280 29096
rect 25228 29053 25237 29087
rect 25237 29053 25271 29087
rect 25271 29053 25280 29087
rect 25228 29044 25280 29053
rect 25872 29044 25924 29096
rect 27620 29112 27672 29164
rect 28172 29155 28224 29164
rect 28172 29121 28181 29155
rect 28181 29121 28215 29155
rect 28215 29121 28224 29155
rect 28172 29112 28224 29121
rect 30564 29248 30616 29300
rect 32404 29248 32456 29300
rect 32588 29248 32640 29300
rect 29368 29223 29420 29232
rect 29368 29189 29377 29223
rect 29377 29189 29411 29223
rect 29411 29189 29420 29223
rect 29368 29180 29420 29189
rect 29644 29155 29696 29164
rect 27988 29044 28040 29096
rect 27068 28976 27120 29028
rect 27528 28976 27580 29028
rect 28356 28976 28408 29028
rect 29644 29121 29653 29155
rect 29653 29121 29687 29155
rect 29687 29121 29696 29155
rect 29644 29112 29696 29121
rect 30472 29180 30524 29232
rect 30748 29180 30800 29232
rect 32772 29180 32824 29232
rect 33232 29180 33284 29232
rect 36084 29223 36136 29232
rect 36084 29189 36093 29223
rect 36093 29189 36127 29223
rect 36127 29189 36136 29223
rect 36084 29180 36136 29189
rect 28724 29019 28776 29028
rect 28724 28985 28733 29019
rect 28733 28985 28767 29019
rect 28767 28985 28776 29019
rect 28724 28976 28776 28985
rect 31300 29112 31352 29164
rect 31760 29112 31812 29164
rect 35716 29155 35768 29164
rect 31576 29044 31628 29096
rect 33048 29044 33100 29096
rect 35716 29121 35725 29155
rect 35725 29121 35759 29155
rect 35759 29121 35768 29155
rect 35716 29112 35768 29121
rect 35808 29155 35860 29164
rect 35808 29121 35818 29155
rect 35818 29121 35852 29155
rect 35852 29121 35860 29155
rect 35808 29112 35860 29121
rect 35992 29155 36044 29164
rect 35992 29121 36001 29155
rect 36001 29121 36035 29155
rect 36035 29121 36044 29155
rect 35992 29112 36044 29121
rect 36268 29112 36320 29164
rect 37924 29112 37976 29164
rect 37740 29087 37792 29096
rect 37740 29053 37749 29087
rect 37749 29053 37783 29087
rect 37783 29053 37792 29087
rect 37740 29044 37792 29053
rect 36636 28976 36688 29028
rect 25320 28908 25372 28960
rect 26240 28908 26292 28960
rect 29368 28951 29420 28960
rect 29368 28917 29377 28951
rect 29377 28917 29411 28951
rect 29411 28917 29420 28951
rect 29368 28908 29420 28917
rect 32496 28951 32548 28960
rect 32496 28917 32505 28951
rect 32505 28917 32539 28951
rect 32539 28917 32548 28951
rect 32496 28908 32548 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 4804 28704 4856 28756
rect 4712 28500 4764 28552
rect 6184 28704 6236 28756
rect 7380 28704 7432 28756
rect 9220 28704 9272 28756
rect 11060 28747 11112 28756
rect 11060 28713 11069 28747
rect 11069 28713 11103 28747
rect 11103 28713 11112 28747
rect 11060 28704 11112 28713
rect 11888 28704 11940 28756
rect 11980 28747 12032 28756
rect 11980 28713 11989 28747
rect 11989 28713 12023 28747
rect 12023 28713 12032 28747
rect 11980 28704 12032 28713
rect 14004 28704 14056 28756
rect 14832 28747 14884 28756
rect 14832 28713 14841 28747
rect 14841 28713 14875 28747
rect 14875 28713 14884 28747
rect 14832 28704 14884 28713
rect 15568 28704 15620 28756
rect 5540 28636 5592 28688
rect 5356 28543 5408 28552
rect 5356 28509 5365 28543
rect 5365 28509 5399 28543
rect 5399 28509 5408 28543
rect 5356 28500 5408 28509
rect 6920 28500 6972 28552
rect 8576 28568 8628 28620
rect 8300 28543 8352 28552
rect 5448 28475 5500 28484
rect 5448 28441 5457 28475
rect 5457 28441 5491 28475
rect 5491 28441 5500 28475
rect 5448 28432 5500 28441
rect 6460 28432 6512 28484
rect 6736 28432 6788 28484
rect 7012 28475 7064 28484
rect 7012 28441 7021 28475
rect 7021 28441 7055 28475
rect 7055 28441 7064 28475
rect 7012 28432 7064 28441
rect 5724 28407 5776 28416
rect 5724 28373 5733 28407
rect 5733 28373 5767 28407
rect 5767 28373 5776 28407
rect 5724 28364 5776 28373
rect 8300 28509 8309 28543
rect 8309 28509 8343 28543
rect 8343 28509 8352 28543
rect 8300 28500 8352 28509
rect 9128 28543 9180 28552
rect 8116 28432 8168 28484
rect 9128 28509 9137 28543
rect 9137 28509 9171 28543
rect 9171 28509 9180 28543
rect 9128 28500 9180 28509
rect 13544 28636 13596 28688
rect 15200 28636 15252 28688
rect 16856 28704 16908 28756
rect 17316 28704 17368 28756
rect 18512 28704 18564 28756
rect 11152 28568 11204 28620
rect 13360 28568 13412 28620
rect 14372 28568 14424 28620
rect 16764 28636 16816 28688
rect 17684 28636 17736 28688
rect 8484 28432 8536 28484
rect 10416 28432 10468 28484
rect 10968 28432 11020 28484
rect 8024 28364 8076 28416
rect 9128 28364 9180 28416
rect 11612 28364 11664 28416
rect 14280 28543 14332 28552
rect 14280 28509 14289 28543
rect 14289 28509 14323 28543
rect 14323 28509 14332 28543
rect 14280 28500 14332 28509
rect 14464 28543 14516 28552
rect 14464 28509 14473 28543
rect 14473 28509 14507 28543
rect 14507 28509 14516 28543
rect 14464 28500 14516 28509
rect 14648 28543 14700 28552
rect 14648 28509 14657 28543
rect 14657 28509 14691 28543
rect 14691 28509 14700 28543
rect 14648 28500 14700 28509
rect 16304 28543 16356 28552
rect 16304 28509 16313 28543
rect 16313 28509 16347 28543
rect 16347 28509 16356 28543
rect 16304 28500 16356 28509
rect 16764 28543 16816 28552
rect 11796 28475 11848 28484
rect 11796 28441 11805 28475
rect 11805 28441 11839 28475
rect 11839 28441 11848 28475
rect 11796 28432 11848 28441
rect 16212 28432 16264 28484
rect 16764 28509 16773 28543
rect 16773 28509 16807 28543
rect 16807 28509 16816 28543
rect 16764 28500 16816 28509
rect 19340 28636 19392 28688
rect 20444 28636 20496 28688
rect 17868 28500 17920 28552
rect 17040 28432 17092 28484
rect 18880 28500 18932 28552
rect 19432 28500 19484 28552
rect 19616 28500 19668 28552
rect 20628 28568 20680 28620
rect 21548 28704 21600 28756
rect 23480 28704 23532 28756
rect 24860 28704 24912 28756
rect 25964 28704 26016 28756
rect 27252 28704 27304 28756
rect 27988 28704 28040 28756
rect 30196 28704 30248 28756
rect 32588 28704 32640 28756
rect 35348 28704 35400 28756
rect 35716 28704 35768 28756
rect 26240 28636 26292 28688
rect 28448 28636 28500 28688
rect 28908 28636 28960 28688
rect 20536 28500 20588 28552
rect 21364 28500 21416 28552
rect 21640 28500 21692 28552
rect 21824 28500 21876 28552
rect 25872 28568 25924 28620
rect 12716 28364 12768 28416
rect 13268 28364 13320 28416
rect 15016 28364 15068 28416
rect 22652 28432 22704 28484
rect 22100 28364 22152 28416
rect 22928 28364 22980 28416
rect 24676 28500 24728 28552
rect 30012 28568 30064 28620
rect 28356 28543 28408 28552
rect 28356 28509 28365 28543
rect 28365 28509 28399 28543
rect 28399 28509 28408 28543
rect 28356 28500 28408 28509
rect 28816 28500 28868 28552
rect 31668 28636 31720 28688
rect 30472 28611 30524 28620
rect 30472 28577 30481 28611
rect 30481 28577 30515 28611
rect 30515 28577 30524 28611
rect 30472 28568 30524 28577
rect 30380 28500 30432 28552
rect 30564 28500 30616 28552
rect 31300 28543 31352 28552
rect 31300 28509 31309 28543
rect 31309 28509 31343 28543
rect 31343 28509 31352 28543
rect 31300 28500 31352 28509
rect 31392 28543 31444 28552
rect 31392 28509 31402 28543
rect 31402 28509 31436 28543
rect 31436 28509 31444 28543
rect 31392 28500 31444 28509
rect 31576 28543 31628 28552
rect 31576 28509 31585 28543
rect 31585 28509 31619 28543
rect 31619 28509 31628 28543
rect 32496 28636 32548 28688
rect 33140 28611 33192 28620
rect 33140 28577 33149 28611
rect 33149 28577 33183 28611
rect 33183 28577 33192 28611
rect 33140 28568 33192 28577
rect 36820 28611 36872 28620
rect 36820 28577 36829 28611
rect 36829 28577 36863 28611
rect 36863 28577 36872 28611
rect 36820 28568 36872 28577
rect 31576 28500 31628 28509
rect 32772 28543 32824 28552
rect 32772 28509 32781 28543
rect 32781 28509 32815 28543
rect 32815 28509 32824 28543
rect 32772 28500 32824 28509
rect 24124 28432 24176 28484
rect 28264 28475 28316 28484
rect 28264 28441 28273 28475
rect 28273 28441 28307 28475
rect 28307 28441 28316 28475
rect 28264 28432 28316 28441
rect 30932 28432 30984 28484
rect 32220 28432 32272 28484
rect 35348 28432 35400 28484
rect 37464 28432 37516 28484
rect 23296 28364 23348 28416
rect 24952 28364 25004 28416
rect 27252 28364 27304 28416
rect 27620 28364 27672 28416
rect 30012 28364 30064 28416
rect 35808 28364 35860 28416
rect 38200 28407 38252 28416
rect 38200 28373 38209 28407
rect 38209 28373 38243 28407
rect 38243 28373 38252 28407
rect 38200 28364 38252 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4804 28024 4856 28076
rect 7104 28160 7156 28212
rect 8484 28160 8536 28212
rect 11060 28203 11112 28212
rect 7380 28092 7432 28144
rect 11060 28169 11069 28203
rect 11069 28169 11103 28203
rect 11103 28169 11112 28203
rect 11060 28160 11112 28169
rect 11796 28160 11848 28212
rect 16948 28203 17000 28212
rect 7564 28024 7616 28076
rect 8300 28067 8352 28076
rect 8300 28033 8309 28067
rect 8309 28033 8343 28067
rect 8343 28033 8352 28067
rect 8300 28024 8352 28033
rect 9036 28024 9088 28076
rect 9312 28092 9364 28144
rect 9588 28092 9640 28144
rect 9404 28067 9456 28076
rect 9404 28033 9413 28067
rect 9413 28033 9447 28067
rect 9447 28033 9456 28067
rect 9404 28024 9456 28033
rect 10232 28067 10284 28076
rect 5264 27956 5316 28008
rect 6368 27956 6420 28008
rect 7840 27956 7892 28008
rect 7104 27888 7156 27940
rect 7564 27888 7616 27940
rect 4988 27863 5040 27872
rect 4988 27829 4997 27863
rect 4997 27829 5031 27863
rect 5031 27829 5040 27863
rect 4988 27820 5040 27829
rect 5080 27820 5132 27872
rect 6736 27820 6788 27872
rect 8300 27820 8352 27872
rect 9864 27956 9916 28008
rect 10232 28033 10241 28067
rect 10241 28033 10275 28067
rect 10275 28033 10284 28067
rect 10232 28024 10284 28033
rect 12716 28067 12768 28076
rect 10140 27999 10192 28008
rect 10140 27965 10149 27999
rect 10149 27965 10183 27999
rect 10183 27965 10192 27999
rect 10140 27956 10192 27965
rect 12716 28033 12725 28067
rect 12725 28033 12759 28067
rect 12759 28033 12768 28067
rect 12716 28024 12768 28033
rect 13268 28092 13320 28144
rect 13728 28024 13780 28076
rect 12072 27956 12124 28008
rect 11428 27888 11480 27940
rect 14372 28067 14424 28076
rect 14372 28033 14381 28067
rect 14381 28033 14415 28067
rect 14415 28033 14424 28067
rect 14372 28024 14424 28033
rect 16948 28169 16957 28203
rect 16957 28169 16991 28203
rect 16991 28169 17000 28203
rect 16948 28160 17000 28169
rect 17592 28160 17644 28212
rect 16764 28092 16816 28144
rect 18788 28092 18840 28144
rect 20444 28092 20496 28144
rect 21548 28092 21600 28144
rect 22560 28135 22612 28144
rect 22560 28101 22569 28135
rect 22569 28101 22603 28135
rect 22603 28101 22612 28135
rect 22560 28092 22612 28101
rect 24308 28092 24360 28144
rect 17040 28067 17092 28076
rect 17040 28033 17049 28067
rect 17049 28033 17083 28067
rect 17083 28033 17092 28067
rect 17040 28024 17092 28033
rect 18604 28024 18656 28076
rect 18880 28067 18932 28076
rect 18880 28033 18889 28067
rect 18889 28033 18923 28067
rect 18923 28033 18932 28067
rect 18880 28024 18932 28033
rect 18972 28024 19024 28076
rect 19984 28024 20036 28076
rect 22100 28067 22152 28076
rect 22100 28033 22109 28067
rect 22109 28033 22143 28067
rect 22143 28033 22152 28067
rect 22100 28024 22152 28033
rect 23112 28024 23164 28076
rect 25780 28160 25832 28212
rect 26516 28160 26568 28212
rect 24860 28092 24912 28144
rect 25228 28092 25280 28144
rect 27160 28135 27212 28144
rect 24676 28024 24728 28076
rect 25504 28067 25556 28076
rect 25504 28033 25513 28067
rect 25513 28033 25547 28067
rect 25547 28033 25556 28067
rect 25504 28024 25556 28033
rect 27160 28101 27169 28135
rect 27169 28101 27203 28135
rect 27203 28101 27212 28135
rect 27160 28092 27212 28101
rect 27988 28092 28040 28144
rect 28448 28135 28500 28144
rect 28448 28101 28457 28135
rect 28457 28101 28491 28135
rect 28491 28101 28500 28135
rect 28448 28092 28500 28101
rect 28908 28160 28960 28212
rect 30104 28160 30156 28212
rect 31116 28160 31168 28212
rect 36268 28203 36320 28212
rect 36268 28169 36277 28203
rect 36277 28169 36311 28203
rect 36311 28169 36320 28203
rect 36268 28160 36320 28169
rect 37464 28203 37516 28212
rect 37464 28169 37473 28203
rect 37473 28169 37507 28203
rect 37507 28169 37516 28203
rect 37464 28160 37516 28169
rect 37924 28203 37976 28212
rect 37924 28169 37933 28203
rect 37933 28169 37967 28203
rect 37967 28169 37976 28203
rect 37924 28160 37976 28169
rect 26700 28024 26752 28076
rect 20168 27999 20220 28008
rect 15660 27888 15712 27940
rect 18420 27888 18472 27940
rect 20168 27965 20177 27999
rect 20177 27965 20211 27999
rect 20211 27965 20220 27999
rect 20168 27956 20220 27965
rect 20720 27956 20772 28008
rect 20996 27956 21048 28008
rect 22284 27956 22336 28008
rect 10324 27820 10376 27872
rect 14556 27863 14608 27872
rect 14556 27829 14565 27863
rect 14565 27829 14599 27863
rect 14599 27829 14608 27863
rect 14556 27820 14608 27829
rect 20076 27863 20128 27872
rect 20076 27829 20085 27863
rect 20085 27829 20119 27863
rect 20119 27829 20128 27863
rect 20076 27820 20128 27829
rect 22008 27820 22060 27872
rect 24032 27931 24084 27940
rect 24032 27897 24041 27931
rect 24041 27897 24075 27931
rect 24075 27897 24084 27931
rect 24032 27888 24084 27897
rect 24676 27888 24728 27940
rect 28816 28024 28868 28076
rect 29920 28092 29972 28144
rect 33140 28092 33192 28144
rect 35808 28092 35860 28144
rect 38200 28092 38252 28144
rect 29644 28024 29696 28076
rect 30012 28024 30064 28076
rect 30196 28067 30248 28076
rect 30196 28033 30206 28067
rect 30206 28033 30240 28067
rect 30240 28033 30248 28067
rect 30196 28024 30248 28033
rect 30564 28067 30616 28076
rect 30564 28033 30578 28067
rect 30578 28033 30612 28067
rect 30612 28033 30616 28067
rect 30564 28024 30616 28033
rect 31208 28024 31260 28076
rect 32680 28024 32732 28076
rect 33048 28024 33100 28076
rect 36084 28067 36136 28076
rect 36084 28033 36093 28067
rect 36093 28033 36127 28067
rect 36127 28033 36136 28067
rect 36084 28024 36136 28033
rect 30380 27956 30432 28008
rect 38016 27999 38068 28008
rect 38016 27965 38025 27999
rect 38025 27965 38059 27999
rect 38059 27965 38068 27999
rect 38016 27956 38068 27965
rect 25964 27888 26016 27940
rect 27344 27888 27396 27940
rect 27528 27888 27580 27940
rect 31392 27888 31444 27940
rect 26148 27820 26200 27872
rect 27436 27863 27488 27872
rect 27436 27829 27445 27863
rect 27445 27829 27479 27863
rect 27479 27829 27488 27863
rect 27436 27820 27488 27829
rect 27804 27863 27856 27872
rect 27804 27829 27813 27863
rect 27813 27829 27847 27863
rect 27847 27829 27856 27863
rect 27804 27820 27856 27829
rect 28816 27863 28868 27872
rect 28816 27829 28825 27863
rect 28825 27829 28859 27863
rect 28859 27829 28868 27863
rect 28816 27820 28868 27829
rect 28908 27820 28960 27872
rect 31944 27820 31996 27872
rect 33232 27820 33284 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 3976 27616 4028 27668
rect 4436 27616 4488 27668
rect 4620 27548 4672 27600
rect 4804 27616 4856 27668
rect 8116 27616 8168 27668
rect 13268 27659 13320 27668
rect 5632 27548 5684 27600
rect 6920 27548 6972 27600
rect 7380 27548 7432 27600
rect 9956 27591 10008 27600
rect 4712 27480 4764 27532
rect 8024 27523 8076 27532
rect 8024 27489 8033 27523
rect 8033 27489 8067 27523
rect 8067 27489 8076 27523
rect 8024 27480 8076 27489
rect 9956 27557 9965 27591
rect 9965 27557 9999 27591
rect 9999 27557 10008 27591
rect 9956 27548 10008 27557
rect 13268 27625 13277 27659
rect 13277 27625 13311 27659
rect 13311 27625 13320 27659
rect 13268 27616 13320 27625
rect 14004 27616 14056 27668
rect 20720 27616 20772 27668
rect 4436 27455 4488 27464
rect 4436 27421 4445 27455
rect 4445 27421 4479 27455
rect 4479 27421 4488 27455
rect 4436 27412 4488 27421
rect 4620 27455 4672 27464
rect 4620 27421 4629 27455
rect 4629 27421 4663 27455
rect 4663 27421 4672 27455
rect 4620 27412 4672 27421
rect 5080 27455 5132 27464
rect 5080 27421 5089 27455
rect 5089 27421 5123 27455
rect 5123 27421 5132 27455
rect 5080 27412 5132 27421
rect 5264 27455 5316 27464
rect 5264 27421 5273 27455
rect 5273 27421 5307 27455
rect 5307 27421 5316 27455
rect 5264 27412 5316 27421
rect 5448 27455 5500 27464
rect 5448 27421 5457 27455
rect 5457 27421 5491 27455
rect 5491 27421 5500 27455
rect 5448 27412 5500 27421
rect 5724 27344 5776 27396
rect 6092 27412 6144 27464
rect 7012 27455 7064 27464
rect 7012 27421 7021 27455
rect 7021 27421 7055 27455
rect 7055 27421 7064 27455
rect 7012 27412 7064 27421
rect 9404 27480 9456 27532
rect 9220 27412 9272 27464
rect 13820 27548 13872 27600
rect 15660 27591 15712 27600
rect 15660 27557 15669 27591
rect 15669 27557 15703 27591
rect 15703 27557 15712 27591
rect 15660 27548 15712 27557
rect 17040 27548 17092 27600
rect 21640 27616 21692 27668
rect 23296 27616 23348 27668
rect 26792 27616 26844 27668
rect 27160 27616 27212 27668
rect 18972 27480 19024 27532
rect 3976 27319 4028 27328
rect 3976 27285 3985 27319
rect 3985 27285 4019 27319
rect 4019 27285 4028 27319
rect 3976 27276 4028 27285
rect 4528 27276 4580 27328
rect 7840 27319 7892 27328
rect 7840 27285 7849 27319
rect 7849 27285 7883 27319
rect 7883 27285 7892 27319
rect 7840 27276 7892 27285
rect 8116 27344 8168 27396
rect 9036 27344 9088 27396
rect 9588 27387 9640 27396
rect 9588 27353 9597 27387
rect 9597 27353 9631 27387
rect 9631 27353 9640 27387
rect 9588 27344 9640 27353
rect 9864 27344 9916 27396
rect 11428 27412 11480 27464
rect 11796 27344 11848 27396
rect 14188 27412 14240 27464
rect 14556 27455 14608 27464
rect 14556 27421 14590 27455
rect 14590 27421 14608 27455
rect 14556 27412 14608 27421
rect 17684 27412 17736 27464
rect 18880 27412 18932 27464
rect 19064 27412 19116 27464
rect 10140 27276 10192 27328
rect 10600 27319 10652 27328
rect 10600 27285 10609 27319
rect 10609 27285 10643 27319
rect 10643 27285 10652 27319
rect 10600 27276 10652 27285
rect 11244 27319 11296 27328
rect 11244 27285 11253 27319
rect 11253 27285 11287 27319
rect 11287 27285 11296 27319
rect 11244 27276 11296 27285
rect 18328 27344 18380 27396
rect 19156 27344 19208 27396
rect 21916 27548 21968 27600
rect 25872 27548 25924 27600
rect 20076 27412 20128 27464
rect 21916 27344 21968 27396
rect 24124 27480 24176 27532
rect 25596 27480 25648 27532
rect 22744 27455 22796 27464
rect 22744 27421 22753 27455
rect 22753 27421 22787 27455
rect 22787 27421 22796 27455
rect 22744 27412 22796 27421
rect 23480 27455 23532 27464
rect 23480 27421 23489 27455
rect 23489 27421 23523 27455
rect 23523 27421 23532 27455
rect 23480 27412 23532 27421
rect 25504 27412 25556 27464
rect 26424 27412 26476 27464
rect 24492 27344 24544 27396
rect 26608 27415 26614 27430
rect 26614 27415 26648 27430
rect 26648 27415 26660 27430
rect 26608 27378 26660 27415
rect 26700 27455 26752 27464
rect 26700 27421 26709 27455
rect 26709 27421 26743 27455
rect 26743 27421 26752 27455
rect 26700 27412 26752 27421
rect 26884 27455 26936 27464
rect 26884 27421 26893 27455
rect 26893 27421 26927 27455
rect 26927 27421 26936 27455
rect 26884 27412 26936 27421
rect 18420 27276 18472 27328
rect 18512 27276 18564 27328
rect 25780 27276 25832 27328
rect 27252 27276 27304 27328
rect 27620 27455 27672 27464
rect 27620 27421 27629 27455
rect 27629 27421 27663 27455
rect 27663 27421 27672 27455
rect 27620 27412 27672 27421
rect 31300 27616 31352 27668
rect 30380 27548 30432 27600
rect 35532 27548 35584 27600
rect 29276 27480 29328 27532
rect 30104 27480 30156 27532
rect 28448 27412 28500 27464
rect 28908 27412 28960 27464
rect 29092 27344 29144 27396
rect 30472 27412 30524 27464
rect 30288 27387 30340 27396
rect 30288 27353 30297 27387
rect 30297 27353 30331 27387
rect 30331 27353 30340 27387
rect 30288 27344 30340 27353
rect 28448 27276 28500 27328
rect 29368 27276 29420 27328
rect 29736 27319 29788 27328
rect 29736 27285 29745 27319
rect 29745 27285 29779 27319
rect 29779 27285 29788 27319
rect 29736 27276 29788 27285
rect 30012 27276 30064 27328
rect 30932 27455 30984 27464
rect 30932 27421 30942 27455
rect 30942 27421 30976 27455
rect 30976 27421 30984 27455
rect 31208 27480 31260 27532
rect 30932 27412 30984 27421
rect 34796 27480 34848 27532
rect 35808 27480 35860 27532
rect 31208 27387 31260 27396
rect 31208 27353 31217 27387
rect 31217 27353 31251 27387
rect 31251 27353 31260 27387
rect 31208 27344 31260 27353
rect 30932 27276 30984 27328
rect 32864 27412 32916 27464
rect 36912 27455 36964 27464
rect 32036 27344 32088 27396
rect 32220 27387 32272 27396
rect 32220 27353 32229 27387
rect 32229 27353 32263 27387
rect 32263 27353 32272 27387
rect 32220 27344 32272 27353
rect 32772 27344 32824 27396
rect 36912 27421 36921 27455
rect 36921 27421 36955 27455
rect 36955 27421 36964 27455
rect 36912 27412 36964 27421
rect 37096 27412 37148 27464
rect 37188 27387 37240 27396
rect 37188 27353 37197 27387
rect 37197 27353 37231 27387
rect 37231 27353 37240 27387
rect 37188 27344 37240 27353
rect 38108 27387 38160 27396
rect 38108 27353 38117 27387
rect 38117 27353 38151 27387
rect 38151 27353 38160 27387
rect 38108 27344 38160 27353
rect 32496 27319 32548 27328
rect 32496 27285 32505 27319
rect 32505 27285 32539 27319
rect 32539 27285 32548 27319
rect 32496 27276 32548 27285
rect 32956 27276 33008 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 4436 27072 4488 27124
rect 16580 27072 16632 27124
rect 20168 27072 20220 27124
rect 24676 27072 24728 27124
rect 3976 27004 4028 27056
rect 4528 27004 4580 27056
rect 5172 27004 5224 27056
rect 2780 26979 2832 26988
rect 2780 26945 2789 26979
rect 2789 26945 2823 26979
rect 2823 26945 2832 26979
rect 2780 26936 2832 26945
rect 5724 26936 5776 26988
rect 6460 26936 6512 26988
rect 5356 26911 5408 26920
rect 5356 26877 5365 26911
rect 5365 26877 5399 26911
rect 5399 26877 5408 26911
rect 6828 26911 6880 26920
rect 5356 26868 5408 26877
rect 4988 26800 5040 26852
rect 6828 26877 6837 26911
rect 6837 26877 6871 26911
rect 6871 26877 6880 26911
rect 6828 26868 6880 26877
rect 8116 26936 8168 26988
rect 8484 26979 8536 26988
rect 8484 26945 8493 26979
rect 8493 26945 8527 26979
rect 8527 26945 8536 26979
rect 8484 26936 8536 26945
rect 9956 26936 10008 26988
rect 11980 26936 12032 26988
rect 13268 26936 13320 26988
rect 9128 26868 9180 26920
rect 10968 26911 11020 26920
rect 10968 26877 10977 26911
rect 10977 26877 11011 26911
rect 11011 26877 11020 26911
rect 14464 26936 14516 26988
rect 16396 26936 16448 26988
rect 17040 26979 17092 26988
rect 17040 26945 17049 26979
rect 17049 26945 17083 26979
rect 17083 26945 17092 26979
rect 17040 26936 17092 26945
rect 17316 26979 17368 26988
rect 17316 26945 17325 26979
rect 17325 26945 17359 26979
rect 17359 26945 17368 26979
rect 17316 26936 17368 26945
rect 17684 26936 17736 26988
rect 20996 27004 21048 27056
rect 22008 27047 22060 27056
rect 22008 27013 22017 27047
rect 22017 27013 22051 27047
rect 22051 27013 22060 27047
rect 22008 27004 22060 27013
rect 19156 26936 19208 26988
rect 19984 26979 20036 26988
rect 10968 26868 11020 26877
rect 14280 26868 14332 26920
rect 14648 26911 14700 26920
rect 14648 26877 14657 26911
rect 14657 26877 14691 26911
rect 14691 26877 14700 26911
rect 14648 26868 14700 26877
rect 17224 26911 17276 26920
rect 17224 26877 17233 26911
rect 17233 26877 17267 26911
rect 17267 26877 17276 26911
rect 17224 26868 17276 26877
rect 8668 26843 8720 26852
rect 8668 26809 8677 26843
rect 8677 26809 8711 26843
rect 8711 26809 8720 26843
rect 8668 26800 8720 26809
rect 9588 26800 9640 26852
rect 9864 26800 9916 26852
rect 10784 26800 10836 26852
rect 11888 26800 11940 26852
rect 17132 26843 17184 26852
rect 17132 26809 17141 26843
rect 17141 26809 17175 26843
rect 17175 26809 17184 26843
rect 18696 26868 18748 26920
rect 18972 26868 19024 26920
rect 19984 26945 19993 26979
rect 19993 26945 20027 26979
rect 20027 26945 20036 26979
rect 19984 26936 20036 26945
rect 20168 26979 20220 26988
rect 20168 26945 20177 26979
rect 20177 26945 20211 26979
rect 20211 26945 20220 26979
rect 20168 26936 20220 26945
rect 20812 26979 20864 26988
rect 20812 26945 20821 26979
rect 20821 26945 20855 26979
rect 20855 26945 20864 26979
rect 20812 26936 20864 26945
rect 22376 27004 22428 27056
rect 23388 27004 23440 27056
rect 23480 27004 23532 27056
rect 24032 27004 24084 27056
rect 20904 26911 20956 26920
rect 20904 26877 20913 26911
rect 20913 26877 20947 26911
rect 20947 26877 20956 26911
rect 20904 26868 20956 26877
rect 17132 26800 17184 26809
rect 17500 26800 17552 26852
rect 22560 26936 22612 26988
rect 22744 26936 22796 26988
rect 22192 26868 22244 26920
rect 23112 26868 23164 26920
rect 24308 26936 24360 26988
rect 25596 27072 25648 27124
rect 25780 27004 25832 27056
rect 27804 27072 27856 27124
rect 29092 27115 29144 27124
rect 29092 27081 29101 27115
rect 29101 27081 29135 27115
rect 29135 27081 29144 27115
rect 29092 27072 29144 27081
rect 31668 27072 31720 27124
rect 25412 26936 25464 26988
rect 26700 26936 26752 26988
rect 28448 27004 28500 27056
rect 28632 27004 28684 27056
rect 25964 26868 26016 26920
rect 26148 26868 26200 26920
rect 29000 26936 29052 26988
rect 27712 26868 27764 26920
rect 30656 26936 30708 26988
rect 30380 26868 30432 26920
rect 31208 26936 31260 26988
rect 32036 27004 32088 27056
rect 31392 26979 31444 26988
rect 31392 26945 31401 26979
rect 31401 26945 31435 26979
rect 31435 26945 31444 26979
rect 32680 26979 32732 26988
rect 31392 26936 31444 26945
rect 32680 26945 32689 26979
rect 32689 26945 32723 26979
rect 32723 26945 32732 26979
rect 32680 26936 32732 26945
rect 32956 27047 33008 27056
rect 32956 27013 32990 27047
rect 32990 27013 33008 27047
rect 32956 27004 33008 27013
rect 35992 27072 36044 27124
rect 36912 27072 36964 27124
rect 37832 27047 37884 27056
rect 34796 26936 34848 26988
rect 37832 27013 37841 27047
rect 37841 27013 37875 27047
rect 37875 27013 37884 27047
rect 37832 27004 37884 27013
rect 5540 26775 5592 26784
rect 5540 26741 5549 26775
rect 5549 26741 5583 26775
rect 5583 26741 5592 26775
rect 5540 26732 5592 26741
rect 6828 26732 6880 26784
rect 7380 26732 7432 26784
rect 9220 26775 9272 26784
rect 9220 26741 9229 26775
rect 9229 26741 9263 26775
rect 9263 26741 9272 26775
rect 9220 26732 9272 26741
rect 10876 26732 10928 26784
rect 13176 26775 13228 26784
rect 13176 26741 13185 26775
rect 13185 26741 13219 26775
rect 13219 26741 13228 26775
rect 13176 26732 13228 26741
rect 15568 26732 15620 26784
rect 19064 26775 19116 26784
rect 19064 26741 19073 26775
rect 19073 26741 19107 26775
rect 19107 26741 19116 26775
rect 19064 26732 19116 26741
rect 21916 26732 21968 26784
rect 22376 26732 22428 26784
rect 32128 26800 32180 26852
rect 33876 26800 33928 26852
rect 34612 26800 34664 26852
rect 35808 26936 35860 26988
rect 36360 26979 36412 26988
rect 36360 26945 36369 26979
rect 36369 26945 36403 26979
rect 36403 26945 36412 26979
rect 36360 26936 36412 26945
rect 36636 26979 36688 26988
rect 36636 26945 36645 26979
rect 36645 26945 36679 26979
rect 36679 26945 36688 26979
rect 36636 26936 36688 26945
rect 38016 26911 38068 26920
rect 38016 26877 38025 26911
rect 38025 26877 38059 26911
rect 38059 26877 38068 26911
rect 38016 26868 38068 26877
rect 23296 26732 23348 26784
rect 24584 26732 24636 26784
rect 26884 26732 26936 26784
rect 30748 26732 30800 26784
rect 33416 26732 33468 26784
rect 35808 26732 35860 26784
rect 36544 26775 36596 26784
rect 36544 26741 36553 26775
rect 36553 26741 36587 26775
rect 36587 26741 36596 26775
rect 36544 26732 36596 26741
rect 37464 26775 37516 26784
rect 37464 26741 37473 26775
rect 37473 26741 37507 26775
rect 37507 26741 37516 26775
rect 37464 26732 37516 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 4528 26528 4580 26580
rect 4804 26528 4856 26580
rect 5172 26528 5224 26580
rect 5540 26528 5592 26580
rect 9128 26571 9180 26580
rect 9128 26537 9137 26571
rect 9137 26537 9171 26571
rect 9171 26537 9180 26571
rect 9128 26528 9180 26537
rect 4436 26460 4488 26512
rect 4804 26392 4856 26444
rect 5264 26460 5316 26512
rect 6276 26460 6328 26512
rect 7656 26460 7708 26512
rect 5172 26367 5224 26376
rect 5172 26333 5181 26367
rect 5181 26333 5215 26367
rect 5215 26333 5224 26367
rect 5172 26324 5224 26333
rect 5540 26324 5592 26376
rect 7012 26392 7064 26444
rect 6276 26367 6328 26376
rect 6276 26333 6285 26367
rect 6285 26333 6319 26367
rect 6319 26333 6328 26367
rect 6736 26367 6788 26376
rect 6276 26324 6328 26333
rect 6736 26333 6745 26367
rect 6745 26333 6779 26367
rect 6779 26333 6788 26367
rect 6736 26324 6788 26333
rect 7196 26324 7248 26376
rect 11244 26528 11296 26580
rect 11980 26571 12032 26580
rect 11980 26537 11989 26571
rect 11989 26537 12023 26571
rect 12023 26537 12032 26571
rect 13268 26571 13320 26580
rect 11980 26528 12032 26537
rect 9680 26460 9732 26512
rect 9772 26460 9824 26512
rect 10140 26460 10192 26512
rect 13268 26537 13277 26571
rect 13277 26537 13311 26571
rect 13311 26537 13320 26571
rect 13268 26528 13320 26537
rect 16672 26528 16724 26580
rect 17592 26528 17644 26580
rect 18420 26528 18472 26580
rect 21824 26528 21876 26580
rect 22008 26528 22060 26580
rect 22744 26571 22796 26580
rect 22744 26537 22753 26571
rect 22753 26537 22787 26571
rect 22787 26537 22796 26571
rect 22744 26528 22796 26537
rect 28908 26528 28960 26580
rect 30196 26528 30248 26580
rect 34796 26528 34848 26580
rect 36360 26528 36412 26580
rect 37832 26528 37884 26580
rect 17316 26460 17368 26512
rect 20260 26460 20312 26512
rect 10508 26392 10560 26444
rect 11796 26392 11848 26444
rect 12256 26392 12308 26444
rect 8484 26256 8536 26308
rect 9496 26333 9505 26354
rect 9505 26333 9539 26354
rect 9539 26333 9548 26354
rect 9496 26302 9548 26333
rect 9864 26324 9916 26376
rect 10876 26367 10928 26376
rect 10876 26333 10910 26367
rect 10910 26333 10928 26367
rect 10876 26324 10928 26333
rect 13544 26324 13596 26376
rect 14648 26324 14700 26376
rect 15568 26367 15620 26376
rect 15568 26333 15577 26367
rect 15577 26333 15611 26367
rect 15611 26333 15620 26367
rect 15568 26324 15620 26333
rect 9588 26299 9640 26308
rect 9588 26265 9623 26299
rect 9623 26265 9640 26299
rect 9588 26256 9640 26265
rect 4712 26188 4764 26240
rect 5172 26188 5224 26240
rect 5264 26188 5316 26240
rect 8392 26188 8444 26240
rect 15016 26256 15068 26308
rect 15108 26256 15160 26308
rect 16028 26367 16080 26376
rect 16028 26333 16037 26367
rect 16037 26333 16071 26367
rect 16071 26333 16080 26367
rect 16028 26324 16080 26333
rect 16948 26324 17000 26376
rect 17132 26367 17184 26376
rect 17132 26333 17141 26367
rect 17141 26333 17175 26367
rect 17175 26333 17184 26367
rect 17132 26324 17184 26333
rect 17224 26324 17276 26376
rect 18144 26392 18196 26444
rect 17592 26324 17644 26376
rect 20628 26367 20680 26376
rect 20628 26333 20637 26367
rect 20637 26333 20671 26367
rect 20671 26333 20680 26367
rect 20628 26324 20680 26333
rect 20720 26324 20772 26376
rect 21272 26460 21324 26512
rect 22008 26392 22060 26444
rect 17868 26188 17920 26240
rect 21548 26324 21600 26376
rect 28080 26460 28132 26512
rect 28632 26460 28684 26512
rect 32772 26460 32824 26512
rect 22836 26392 22888 26444
rect 22376 26324 22428 26376
rect 23020 26324 23072 26376
rect 23388 26367 23440 26376
rect 23388 26333 23397 26367
rect 23397 26333 23431 26367
rect 23431 26333 23440 26367
rect 23388 26324 23440 26333
rect 24676 26392 24728 26444
rect 24584 26367 24636 26376
rect 24584 26333 24593 26367
rect 24593 26333 24627 26367
rect 24627 26333 24636 26367
rect 24584 26324 24636 26333
rect 24952 26367 25004 26376
rect 24952 26333 24961 26367
rect 24961 26333 24995 26367
rect 24995 26333 25004 26367
rect 24952 26324 25004 26333
rect 25136 26367 25188 26376
rect 25136 26333 25145 26367
rect 25145 26333 25179 26367
rect 25179 26333 25188 26367
rect 27620 26392 27672 26444
rect 28540 26435 28592 26444
rect 28540 26401 28549 26435
rect 28549 26401 28583 26435
rect 28583 26401 28592 26435
rect 28540 26392 28592 26401
rect 32404 26392 32456 26444
rect 32496 26392 32548 26444
rect 25136 26324 25188 26333
rect 26332 26324 26384 26376
rect 28080 26324 28132 26376
rect 32128 26324 32180 26376
rect 33140 26367 33192 26376
rect 33140 26333 33149 26367
rect 33149 26333 33183 26367
rect 33183 26333 33192 26367
rect 33140 26324 33192 26333
rect 33232 26367 33284 26376
rect 33232 26333 33241 26367
rect 33241 26333 33275 26367
rect 33275 26333 33284 26367
rect 33416 26367 33468 26376
rect 33232 26324 33284 26333
rect 33416 26333 33425 26367
rect 33425 26333 33459 26367
rect 33459 26333 33468 26367
rect 33416 26324 33468 26333
rect 33600 26392 33652 26444
rect 33968 26367 34020 26376
rect 33968 26333 33977 26367
rect 33977 26333 34011 26367
rect 34011 26333 34020 26367
rect 33968 26324 34020 26333
rect 34152 26367 34204 26376
rect 34152 26333 34161 26367
rect 34161 26333 34195 26367
rect 34195 26333 34204 26367
rect 34152 26324 34204 26333
rect 35440 26367 35492 26376
rect 35440 26333 35449 26367
rect 35449 26333 35483 26367
rect 35483 26333 35492 26367
rect 35440 26324 35492 26333
rect 35532 26367 35584 26376
rect 35532 26333 35541 26367
rect 35541 26333 35575 26367
rect 35575 26333 35584 26367
rect 35532 26324 35584 26333
rect 35808 26367 35860 26376
rect 35808 26333 35817 26367
rect 35817 26333 35851 26367
rect 35851 26333 35860 26367
rect 35808 26324 35860 26333
rect 36820 26324 36872 26376
rect 37464 26324 37516 26376
rect 25780 26299 25832 26308
rect 21640 26231 21692 26240
rect 21640 26197 21649 26231
rect 21649 26197 21683 26231
rect 21683 26197 21692 26231
rect 21640 26188 21692 26197
rect 24032 26188 24084 26240
rect 25320 26231 25372 26240
rect 25320 26197 25329 26231
rect 25329 26197 25363 26231
rect 25363 26197 25372 26231
rect 25320 26188 25372 26197
rect 25780 26265 25789 26299
rect 25789 26265 25823 26299
rect 25823 26265 25832 26299
rect 25780 26256 25832 26265
rect 25964 26299 26016 26308
rect 25964 26265 25973 26299
rect 25973 26265 26007 26299
rect 26007 26265 26016 26299
rect 25964 26256 26016 26265
rect 26424 26256 26476 26308
rect 37096 26256 37148 26308
rect 26148 26231 26200 26240
rect 26148 26197 26157 26231
rect 26157 26197 26191 26231
rect 26191 26197 26200 26231
rect 26148 26188 26200 26197
rect 28448 26231 28500 26240
rect 28448 26197 28457 26231
rect 28457 26197 28491 26231
rect 28491 26197 28500 26231
rect 28448 26188 28500 26197
rect 30564 26231 30616 26240
rect 30564 26197 30573 26231
rect 30573 26197 30607 26231
rect 30607 26197 30616 26231
rect 30564 26188 30616 26197
rect 30932 26231 30984 26240
rect 30932 26197 30941 26231
rect 30941 26197 30975 26231
rect 30975 26197 30984 26231
rect 30932 26188 30984 26197
rect 31300 26188 31352 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 5080 25984 5132 26036
rect 6368 25916 6420 25968
rect 6736 25891 6788 25900
rect 4896 25780 4948 25832
rect 6736 25857 6745 25891
rect 6745 25857 6779 25891
rect 6779 25857 6788 25891
rect 6736 25848 6788 25857
rect 7932 25984 7984 26036
rect 8208 26027 8260 26036
rect 8208 25993 8217 26027
rect 8217 25993 8251 26027
rect 8251 25993 8260 26027
rect 8208 25984 8260 25993
rect 9864 25984 9916 26036
rect 15108 25984 15160 26036
rect 16948 25984 17000 26036
rect 18144 26027 18196 26036
rect 18144 25993 18153 26027
rect 18153 25993 18187 26027
rect 18187 25993 18196 26027
rect 18144 25984 18196 25993
rect 9404 25916 9456 25968
rect 13176 25916 13228 25968
rect 8484 25848 8536 25900
rect 9220 25848 9272 25900
rect 9956 25848 10008 25900
rect 10600 25848 10652 25900
rect 10876 25848 10928 25900
rect 17040 25848 17092 25900
rect 17684 25848 17736 25900
rect 19984 25916 20036 25968
rect 18604 25891 18656 25900
rect 18604 25857 18613 25891
rect 18613 25857 18647 25891
rect 18647 25857 18656 25891
rect 18604 25848 18656 25857
rect 20352 25848 20404 25900
rect 13176 25823 13228 25832
rect 13176 25789 13185 25823
rect 13185 25789 13219 25823
rect 13219 25789 13228 25823
rect 13176 25780 13228 25789
rect 21640 25984 21692 26036
rect 22468 25984 22520 26036
rect 23848 25984 23900 26036
rect 24584 25984 24636 26036
rect 32128 25984 32180 26036
rect 32864 25984 32916 26036
rect 23020 25916 23072 25968
rect 20720 25848 20772 25900
rect 20904 25848 20956 25900
rect 21456 25848 21508 25900
rect 4436 25712 4488 25764
rect 7472 25712 7524 25764
rect 19340 25712 19392 25764
rect 20996 25780 21048 25832
rect 23572 25848 23624 25900
rect 24492 25848 24544 25900
rect 25044 25916 25096 25968
rect 31024 25916 31076 25968
rect 35348 25916 35400 25968
rect 26148 25848 26200 25900
rect 27528 25891 27580 25900
rect 27528 25857 27537 25891
rect 27537 25857 27571 25891
rect 27571 25857 27580 25891
rect 27528 25848 27580 25857
rect 20076 25712 20128 25764
rect 20444 25712 20496 25764
rect 20628 25712 20680 25764
rect 25412 25780 25464 25832
rect 26700 25780 26752 25832
rect 27160 25780 27212 25832
rect 27988 25780 28040 25832
rect 28448 25848 28500 25900
rect 33140 25891 33192 25900
rect 33140 25857 33149 25891
rect 33149 25857 33183 25891
rect 33183 25857 33192 25891
rect 33140 25848 33192 25857
rect 34152 25848 34204 25900
rect 37924 25848 37976 25900
rect 24584 25712 24636 25764
rect 24860 25755 24912 25764
rect 24860 25721 24869 25755
rect 24869 25721 24903 25755
rect 24903 25721 24912 25755
rect 24860 25712 24912 25721
rect 26240 25712 26292 25764
rect 28356 25780 28408 25832
rect 28816 25780 28868 25832
rect 29000 25823 29052 25832
rect 29000 25789 29009 25823
rect 29009 25789 29043 25823
rect 29043 25789 29052 25823
rect 29000 25780 29052 25789
rect 31760 25780 31812 25832
rect 32680 25780 32732 25832
rect 33968 25780 34020 25832
rect 38108 25823 38160 25832
rect 38108 25789 38117 25823
rect 38117 25789 38151 25823
rect 38151 25789 38160 25823
rect 38108 25780 38160 25789
rect 4896 25644 4948 25696
rect 5172 25687 5224 25696
rect 5172 25653 5181 25687
rect 5181 25653 5215 25687
rect 5215 25653 5224 25687
rect 5172 25644 5224 25653
rect 6460 25644 6512 25696
rect 8116 25644 8168 25696
rect 9312 25644 9364 25696
rect 10600 25644 10652 25696
rect 17224 25687 17276 25696
rect 17224 25653 17233 25687
rect 17233 25653 17267 25687
rect 17267 25653 17276 25687
rect 17224 25644 17276 25653
rect 28172 25644 28224 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 5632 25440 5684 25492
rect 8392 25440 8444 25492
rect 10324 25440 10376 25492
rect 5172 25372 5224 25424
rect 8024 25372 8076 25424
rect 4712 25304 4764 25356
rect 4896 25347 4948 25356
rect 4896 25313 4905 25347
rect 4905 25313 4939 25347
rect 4939 25313 4948 25347
rect 4896 25304 4948 25313
rect 5448 25304 5500 25356
rect 6460 25347 6512 25356
rect 6460 25313 6469 25347
rect 6469 25313 6503 25347
rect 6503 25313 6512 25347
rect 6460 25304 6512 25313
rect 6920 25304 6972 25356
rect 4160 25279 4212 25288
rect 4160 25245 4169 25279
rect 4169 25245 4203 25279
rect 4203 25245 4212 25279
rect 4160 25236 4212 25245
rect 4436 25279 4488 25288
rect 4436 25245 4445 25279
rect 4445 25245 4479 25279
rect 4479 25245 4488 25279
rect 5356 25279 5408 25288
rect 4436 25236 4488 25245
rect 5356 25245 5365 25279
rect 5365 25245 5399 25279
rect 5399 25245 5408 25279
rect 5356 25236 5408 25245
rect 9680 25304 9732 25356
rect 8116 25279 8168 25288
rect 8116 25245 8125 25279
rect 8125 25245 8159 25279
rect 8159 25245 8168 25279
rect 8392 25279 8444 25288
rect 8116 25236 8168 25245
rect 8392 25245 8401 25279
rect 8401 25245 8435 25279
rect 8435 25245 8444 25279
rect 8392 25236 8444 25245
rect 3976 25143 4028 25152
rect 3976 25109 3985 25143
rect 3985 25109 4019 25143
rect 4019 25109 4028 25143
rect 3976 25100 4028 25109
rect 5540 25143 5592 25152
rect 5540 25109 5549 25143
rect 5549 25109 5583 25143
rect 5583 25109 5592 25143
rect 5540 25100 5592 25109
rect 7472 25100 7524 25152
rect 10600 25236 10652 25288
rect 19156 25440 19208 25492
rect 21364 25440 21416 25492
rect 26240 25440 26292 25492
rect 28080 25440 28132 25492
rect 16580 25415 16632 25424
rect 16580 25381 16589 25415
rect 16589 25381 16623 25415
rect 16623 25381 16632 25415
rect 16580 25372 16632 25381
rect 13728 25304 13780 25356
rect 10876 25279 10928 25288
rect 10876 25245 10885 25279
rect 10885 25245 10919 25279
rect 10919 25245 10928 25279
rect 10876 25236 10928 25245
rect 13176 25236 13228 25288
rect 14188 25236 14240 25288
rect 14648 25279 14700 25288
rect 14648 25245 14657 25279
rect 14657 25245 14691 25279
rect 14691 25245 14700 25279
rect 14648 25236 14700 25245
rect 9220 25100 9272 25152
rect 9496 25143 9548 25152
rect 9496 25109 9505 25143
rect 9505 25109 9539 25143
rect 9539 25109 9548 25143
rect 9496 25100 9548 25109
rect 13544 25168 13596 25220
rect 15660 25168 15712 25220
rect 14832 25143 14884 25152
rect 14832 25109 14841 25143
rect 14841 25109 14875 25143
rect 14875 25109 14884 25143
rect 14832 25100 14884 25109
rect 18512 25372 18564 25424
rect 18788 25372 18840 25424
rect 19248 25372 19300 25424
rect 18328 25347 18380 25356
rect 18328 25313 18337 25347
rect 18337 25313 18371 25347
rect 18371 25313 18380 25347
rect 18328 25304 18380 25313
rect 17684 25236 17736 25288
rect 18604 25236 18656 25288
rect 18880 25279 18932 25288
rect 18880 25245 18889 25279
rect 18889 25245 18923 25279
rect 18923 25245 18932 25279
rect 18880 25236 18932 25245
rect 19432 25236 19484 25288
rect 20996 25279 21048 25288
rect 17868 25168 17920 25220
rect 20996 25245 21005 25279
rect 21005 25245 21039 25279
rect 21039 25245 21048 25279
rect 20996 25236 21048 25245
rect 21640 25279 21692 25288
rect 21640 25245 21649 25279
rect 21649 25245 21683 25279
rect 21683 25245 21692 25279
rect 21640 25236 21692 25245
rect 21824 25279 21876 25288
rect 21824 25245 21833 25279
rect 21833 25245 21867 25279
rect 21867 25245 21876 25279
rect 21824 25236 21876 25245
rect 24768 25372 24820 25424
rect 24860 25372 24912 25424
rect 29920 25440 29972 25492
rect 28908 25372 28960 25424
rect 33140 25372 33192 25424
rect 25412 25304 25464 25356
rect 25688 25304 25740 25356
rect 25872 25304 25924 25356
rect 24952 25279 25004 25288
rect 20720 25168 20772 25220
rect 24952 25245 24961 25279
rect 24961 25245 24995 25279
rect 24995 25245 25004 25279
rect 24952 25236 25004 25245
rect 25228 25236 25280 25288
rect 26148 25236 26200 25288
rect 26332 25236 26384 25288
rect 25504 25168 25556 25220
rect 26056 25168 26108 25220
rect 26884 25236 26936 25288
rect 28448 25279 28500 25288
rect 28448 25245 28457 25279
rect 28457 25245 28491 25279
rect 28491 25245 28500 25279
rect 28448 25236 28500 25245
rect 28632 25236 28684 25288
rect 29000 25236 29052 25288
rect 33876 25304 33928 25356
rect 34060 25347 34112 25356
rect 34060 25313 34069 25347
rect 34069 25313 34103 25347
rect 34103 25313 34112 25347
rect 34060 25304 34112 25313
rect 31760 25236 31812 25288
rect 27712 25168 27764 25220
rect 29644 25168 29696 25220
rect 30564 25168 30616 25220
rect 17316 25100 17368 25152
rect 17776 25100 17828 25152
rect 18972 25100 19024 25152
rect 19432 25100 19484 25152
rect 20536 25143 20588 25152
rect 20536 25109 20545 25143
rect 20545 25109 20579 25143
rect 20579 25109 20588 25143
rect 20536 25100 20588 25109
rect 23020 25143 23072 25152
rect 23020 25109 23029 25143
rect 23029 25109 23063 25143
rect 23063 25109 23072 25143
rect 23020 25100 23072 25109
rect 24584 25100 24636 25152
rect 28264 25143 28316 25152
rect 28264 25109 28273 25143
rect 28273 25109 28307 25143
rect 28307 25109 28316 25143
rect 28264 25100 28316 25109
rect 31300 25100 31352 25152
rect 32772 25236 32824 25288
rect 32956 25279 33008 25288
rect 32956 25245 32965 25279
rect 32965 25245 32999 25279
rect 32999 25245 33008 25279
rect 32956 25236 33008 25245
rect 33692 25236 33744 25288
rect 36820 25279 36872 25288
rect 36820 25245 36829 25279
rect 36829 25245 36863 25279
rect 36863 25245 36872 25279
rect 36820 25236 36872 25245
rect 37464 25168 37516 25220
rect 32496 25100 32548 25152
rect 34612 25100 34664 25152
rect 36268 25143 36320 25152
rect 36268 25109 36277 25143
rect 36277 25109 36311 25143
rect 36311 25109 36320 25143
rect 36268 25100 36320 25109
rect 37832 25100 37884 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 4160 24896 4212 24948
rect 5448 24896 5500 24948
rect 8392 24896 8444 24948
rect 3976 24828 4028 24880
rect 2780 24760 2832 24812
rect 4804 24760 4856 24812
rect 5080 24828 5132 24880
rect 5632 24760 5684 24812
rect 6736 24803 6788 24812
rect 6736 24769 6745 24803
rect 6745 24769 6779 24803
rect 6779 24769 6788 24803
rect 6736 24760 6788 24769
rect 6920 24803 6972 24812
rect 6920 24769 6929 24803
rect 6929 24769 6963 24803
rect 6963 24769 6972 24803
rect 6920 24760 6972 24769
rect 7196 24760 7248 24812
rect 8208 24828 8260 24880
rect 7748 24760 7800 24812
rect 9312 24760 9364 24812
rect 9772 24760 9824 24812
rect 18880 24896 18932 24948
rect 19248 24828 19300 24880
rect 6644 24692 6696 24744
rect 8576 24692 8628 24744
rect 9680 24735 9732 24744
rect 9680 24701 9689 24735
rect 9689 24701 9723 24735
rect 9723 24701 9732 24735
rect 9680 24692 9732 24701
rect 10600 24760 10652 24812
rect 7748 24624 7800 24676
rect 10232 24692 10284 24744
rect 10876 24803 10928 24812
rect 10876 24769 10885 24803
rect 10885 24769 10919 24803
rect 10919 24769 10928 24803
rect 10876 24760 10928 24769
rect 11152 24760 11204 24812
rect 14832 24760 14884 24812
rect 16856 24803 16908 24812
rect 16856 24769 16865 24803
rect 16865 24769 16899 24803
rect 16899 24769 16908 24803
rect 16856 24760 16908 24769
rect 17684 24803 17736 24812
rect 17684 24769 17693 24803
rect 17693 24769 17727 24803
rect 17727 24769 17736 24803
rect 17684 24760 17736 24769
rect 17868 24803 17920 24812
rect 17868 24769 17877 24803
rect 17877 24769 17911 24803
rect 17911 24769 17920 24803
rect 17868 24760 17920 24769
rect 18512 24803 18564 24812
rect 18512 24769 18521 24803
rect 18521 24769 18555 24803
rect 18555 24769 18564 24803
rect 18512 24760 18564 24769
rect 19156 24803 19208 24812
rect 19156 24769 19165 24803
rect 19165 24769 19199 24803
rect 19199 24769 19208 24803
rect 19156 24760 19208 24769
rect 12072 24692 12124 24744
rect 14280 24692 14332 24744
rect 15568 24692 15620 24744
rect 20076 24760 20128 24812
rect 21088 24828 21140 24880
rect 22652 24896 22704 24948
rect 25320 24896 25372 24948
rect 26424 24896 26476 24948
rect 32220 24896 32272 24948
rect 32956 24939 33008 24948
rect 24124 24828 24176 24880
rect 19984 24692 20036 24744
rect 23480 24760 23532 24812
rect 23940 24803 23992 24812
rect 23940 24769 23967 24803
rect 23967 24769 23992 24803
rect 23940 24760 23992 24769
rect 25596 24828 25648 24880
rect 25228 24803 25280 24812
rect 4436 24556 4488 24608
rect 5172 24556 5224 24608
rect 7656 24599 7708 24608
rect 7656 24565 7665 24599
rect 7665 24565 7699 24599
rect 7699 24565 7708 24599
rect 7656 24556 7708 24565
rect 9312 24556 9364 24608
rect 9864 24599 9916 24608
rect 9864 24565 9873 24599
rect 9873 24565 9907 24599
rect 9907 24565 9916 24599
rect 9864 24556 9916 24565
rect 10140 24556 10192 24608
rect 10968 24556 11020 24608
rect 19064 24624 19116 24676
rect 19248 24667 19300 24676
rect 19248 24633 19257 24667
rect 19257 24633 19291 24667
rect 19291 24633 19300 24667
rect 19248 24624 19300 24633
rect 19892 24624 19944 24676
rect 20444 24624 20496 24676
rect 23112 24692 23164 24744
rect 23572 24735 23624 24744
rect 23572 24701 23581 24735
rect 23581 24701 23615 24735
rect 23615 24701 23624 24735
rect 23572 24692 23624 24701
rect 25228 24769 25237 24803
rect 25237 24769 25271 24803
rect 25271 24769 25280 24803
rect 25228 24760 25280 24769
rect 25504 24803 25556 24812
rect 25504 24769 25513 24803
rect 25513 24769 25547 24803
rect 25547 24769 25556 24803
rect 25504 24760 25556 24769
rect 27988 24828 28040 24880
rect 31668 24828 31720 24880
rect 32956 24905 32965 24939
rect 32965 24905 32999 24939
rect 32999 24905 33008 24939
rect 32956 24896 33008 24905
rect 33968 24896 34020 24948
rect 37464 24939 37516 24948
rect 37464 24905 37473 24939
rect 37473 24905 37507 24939
rect 37507 24905 37516 24939
rect 37464 24896 37516 24905
rect 37832 24939 37884 24948
rect 37832 24905 37841 24939
rect 37841 24905 37875 24939
rect 37875 24905 37884 24939
rect 37832 24896 37884 24905
rect 25688 24735 25740 24744
rect 25688 24701 25697 24735
rect 25697 24701 25731 24735
rect 25731 24701 25740 24735
rect 25688 24692 25740 24701
rect 26792 24692 26844 24744
rect 27896 24760 27948 24812
rect 14372 24556 14424 24608
rect 15660 24599 15712 24608
rect 15660 24565 15669 24599
rect 15669 24565 15703 24599
rect 15703 24565 15712 24599
rect 15660 24556 15712 24565
rect 16764 24556 16816 24608
rect 18144 24556 18196 24608
rect 20260 24556 20312 24608
rect 22560 24599 22612 24608
rect 22560 24565 22569 24599
rect 22569 24565 22603 24599
rect 22603 24565 22612 24599
rect 22560 24556 22612 24565
rect 22744 24556 22796 24608
rect 28540 24692 28592 24744
rect 29276 24803 29328 24812
rect 29276 24769 29285 24803
rect 29285 24769 29319 24803
rect 29319 24769 29328 24803
rect 29276 24760 29328 24769
rect 29644 24760 29696 24812
rect 30012 24803 30064 24812
rect 30012 24769 30021 24803
rect 30021 24769 30055 24803
rect 30055 24769 30064 24803
rect 30012 24760 30064 24769
rect 28264 24624 28316 24676
rect 29000 24667 29052 24676
rect 29000 24633 29009 24667
rect 29009 24633 29043 24667
rect 29043 24633 29052 24667
rect 29000 24624 29052 24633
rect 29828 24667 29880 24676
rect 29828 24633 29837 24667
rect 29837 24633 29871 24667
rect 29871 24633 29880 24667
rect 29828 24624 29880 24633
rect 32036 24624 32088 24676
rect 32405 24803 32457 24812
rect 32405 24769 32414 24803
rect 32414 24769 32448 24803
rect 32448 24769 32457 24803
rect 32405 24760 32457 24769
rect 32680 24803 32732 24846
rect 32680 24794 32686 24803
rect 32686 24794 32720 24803
rect 32720 24794 32732 24803
rect 33232 24828 33284 24880
rect 34060 24828 34112 24880
rect 36820 24828 36872 24880
rect 33692 24803 33744 24812
rect 32680 24624 32732 24676
rect 29736 24556 29788 24608
rect 30472 24556 30524 24608
rect 33692 24769 33701 24803
rect 33701 24769 33735 24803
rect 33735 24769 33744 24803
rect 33692 24760 33744 24769
rect 34336 24803 34388 24812
rect 34336 24769 34345 24803
rect 34345 24769 34379 24803
rect 34379 24769 34388 24803
rect 34336 24760 34388 24769
rect 34520 24803 34572 24812
rect 34520 24769 34529 24803
rect 34529 24769 34563 24803
rect 34563 24769 34572 24803
rect 34520 24760 34572 24769
rect 34612 24803 34664 24812
rect 34612 24769 34621 24803
rect 34621 24769 34655 24803
rect 34655 24769 34664 24803
rect 34612 24760 34664 24769
rect 35348 24760 35400 24812
rect 37924 24735 37976 24744
rect 37924 24701 37933 24735
rect 37933 24701 37967 24735
rect 37967 24701 37976 24735
rect 37924 24692 37976 24701
rect 38016 24735 38068 24744
rect 38016 24701 38025 24735
rect 38025 24701 38059 24735
rect 38059 24701 38068 24735
rect 38016 24692 38068 24701
rect 34060 24624 34112 24676
rect 34520 24624 34572 24676
rect 36268 24624 36320 24676
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 8392 24352 8444 24404
rect 9404 24352 9456 24404
rect 7196 24284 7248 24336
rect 7932 24327 7984 24336
rect 7932 24293 7941 24327
rect 7941 24293 7975 24327
rect 7975 24293 7984 24327
rect 7932 24284 7984 24293
rect 10416 24352 10468 24404
rect 12072 24395 12124 24404
rect 12072 24361 12081 24395
rect 12081 24361 12115 24395
rect 12115 24361 12124 24395
rect 12072 24352 12124 24361
rect 19248 24352 19300 24404
rect 17684 24284 17736 24336
rect 19892 24284 19944 24336
rect 20352 24284 20404 24336
rect 20536 24284 20588 24336
rect 22376 24352 22428 24404
rect 23388 24352 23440 24404
rect 23940 24352 23992 24404
rect 24584 24352 24636 24404
rect 26516 24352 26568 24404
rect 27896 24395 27948 24404
rect 27896 24361 27905 24395
rect 27905 24361 27939 24395
rect 27939 24361 27948 24395
rect 27896 24352 27948 24361
rect 23572 24284 23624 24336
rect 26148 24284 26200 24336
rect 31300 24352 31352 24404
rect 34336 24352 34388 24404
rect 10508 24216 10560 24268
rect 16764 24259 16816 24268
rect 16764 24225 16773 24259
rect 16773 24225 16807 24259
rect 16807 24225 16816 24259
rect 16764 24216 16816 24225
rect 4160 24080 4212 24132
rect 6828 24080 6880 24132
rect 8208 24123 8260 24132
rect 8208 24089 8217 24123
rect 8217 24089 8251 24123
rect 8251 24089 8260 24123
rect 8208 24080 8260 24089
rect 4804 24012 4856 24064
rect 8300 24055 8352 24064
rect 8300 24021 8309 24055
rect 8309 24021 8343 24055
rect 8343 24021 8352 24055
rect 8300 24012 8352 24021
rect 8760 24148 8812 24200
rect 9220 24148 9272 24200
rect 10968 24191 11020 24200
rect 9312 24123 9364 24132
rect 9312 24089 9321 24123
rect 9321 24089 9355 24123
rect 9355 24089 9364 24123
rect 9312 24080 9364 24089
rect 10968 24157 11002 24191
rect 11002 24157 11020 24191
rect 10968 24148 11020 24157
rect 14280 24191 14332 24200
rect 14280 24157 14289 24191
rect 14289 24157 14323 24191
rect 14323 24157 14332 24191
rect 14280 24148 14332 24157
rect 14372 24148 14424 24200
rect 17224 24216 17276 24268
rect 22376 24216 22428 24268
rect 17316 24191 17368 24200
rect 17316 24157 17325 24191
rect 17325 24157 17359 24191
rect 17359 24157 17368 24191
rect 17316 24148 17368 24157
rect 17592 24148 17644 24200
rect 19156 24148 19208 24200
rect 19892 24080 19944 24132
rect 20260 24191 20312 24200
rect 20260 24157 20269 24191
rect 20269 24157 20303 24191
rect 20303 24157 20312 24191
rect 20260 24148 20312 24157
rect 21824 24148 21876 24200
rect 22744 24148 22796 24200
rect 23020 24191 23072 24200
rect 23020 24157 23029 24191
rect 23029 24157 23063 24191
rect 23063 24157 23072 24191
rect 23020 24148 23072 24157
rect 23296 24191 23348 24200
rect 23296 24157 23305 24191
rect 23305 24157 23339 24191
rect 23339 24157 23348 24191
rect 23296 24148 23348 24157
rect 23388 24148 23440 24200
rect 24032 24191 24084 24200
rect 24032 24157 24041 24191
rect 24041 24157 24075 24191
rect 24075 24157 24084 24191
rect 24032 24148 24084 24157
rect 21364 24080 21416 24132
rect 24768 24191 24820 24200
rect 24768 24157 24777 24191
rect 24777 24157 24811 24191
rect 24811 24157 24820 24191
rect 25964 24191 26016 24200
rect 24768 24148 24820 24157
rect 25964 24157 25973 24191
rect 25973 24157 26007 24191
rect 26007 24157 26016 24191
rect 25964 24148 26016 24157
rect 26332 24191 26384 24200
rect 26332 24157 26341 24191
rect 26341 24157 26375 24191
rect 26375 24157 26384 24191
rect 26332 24148 26384 24157
rect 26516 24216 26568 24268
rect 29828 24216 29880 24268
rect 26700 24148 26752 24200
rect 27160 24148 27212 24200
rect 27436 24191 27488 24200
rect 27436 24157 27443 24191
rect 27443 24157 27488 24191
rect 27436 24148 27488 24157
rect 27804 24148 27856 24200
rect 27896 24148 27948 24200
rect 29276 24148 29328 24200
rect 30564 24216 30616 24268
rect 31668 24216 31720 24268
rect 35256 24284 35308 24336
rect 24952 24080 25004 24132
rect 26424 24080 26476 24132
rect 27528 24123 27580 24132
rect 27528 24089 27537 24123
rect 27537 24089 27571 24123
rect 27571 24089 27580 24123
rect 27528 24080 27580 24089
rect 28080 24080 28132 24132
rect 28356 24080 28408 24132
rect 30012 24080 30064 24132
rect 31944 24191 31996 24200
rect 31944 24157 31954 24191
rect 31954 24157 31988 24191
rect 31988 24157 31996 24191
rect 31944 24148 31996 24157
rect 32128 24191 32180 24200
rect 32128 24157 32137 24191
rect 32137 24157 32171 24191
rect 32171 24157 32180 24191
rect 32588 24216 32640 24268
rect 32128 24148 32180 24157
rect 32680 24148 32732 24200
rect 33140 24191 33192 24200
rect 33140 24157 33147 24191
rect 33147 24157 33192 24191
rect 33140 24148 33192 24157
rect 37832 24191 37884 24200
rect 37832 24157 37841 24191
rect 37841 24157 37875 24191
rect 37875 24157 37884 24191
rect 37832 24148 37884 24157
rect 10232 24012 10284 24064
rect 17592 24012 17644 24064
rect 18144 24055 18196 24064
rect 18144 24021 18153 24055
rect 18153 24021 18187 24055
rect 18187 24021 18196 24055
rect 18144 24012 18196 24021
rect 18788 24055 18840 24064
rect 18788 24021 18797 24055
rect 18797 24021 18831 24055
rect 18831 24021 18840 24055
rect 18788 24012 18840 24021
rect 20996 24012 21048 24064
rect 21088 24055 21140 24064
rect 21088 24021 21097 24055
rect 21097 24021 21131 24055
rect 21131 24021 21140 24055
rect 22652 24055 22704 24064
rect 21088 24012 21140 24021
rect 22652 24021 22661 24055
rect 22661 24021 22695 24055
rect 22695 24021 22704 24055
rect 22652 24012 22704 24021
rect 25504 24012 25556 24064
rect 33232 24123 33284 24132
rect 33232 24089 33241 24123
rect 33241 24089 33275 24123
rect 33275 24089 33284 24123
rect 33232 24080 33284 24089
rect 33324 24123 33376 24132
rect 33324 24089 33333 24123
rect 33333 24089 33367 24123
rect 33367 24089 33376 24123
rect 38108 24123 38160 24132
rect 33324 24080 33376 24089
rect 38108 24089 38117 24123
rect 38117 24089 38151 24123
rect 38151 24089 38160 24123
rect 38108 24080 38160 24089
rect 28540 24012 28592 24064
rect 29184 24012 29236 24064
rect 29552 24012 29604 24064
rect 31944 24012 31996 24064
rect 32404 24012 32456 24064
rect 32588 24012 32640 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4160 23808 4212 23860
rect 4620 23740 4672 23792
rect 2780 23672 2832 23724
rect 3976 23672 4028 23724
rect 4712 23715 4764 23724
rect 4712 23681 4721 23715
rect 4721 23681 4755 23715
rect 4755 23681 4764 23715
rect 4712 23672 4764 23681
rect 5540 23808 5592 23860
rect 5172 23740 5224 23792
rect 16856 23808 16908 23860
rect 18788 23808 18840 23860
rect 21180 23808 21232 23860
rect 23296 23808 23348 23860
rect 23388 23808 23440 23860
rect 5816 23672 5868 23724
rect 7012 23740 7064 23792
rect 7196 23740 7248 23792
rect 6828 23672 6880 23724
rect 7104 23715 7156 23724
rect 7104 23681 7113 23715
rect 7113 23681 7147 23715
rect 7147 23681 7156 23715
rect 7104 23672 7156 23681
rect 6644 23604 6696 23656
rect 7472 23740 7524 23792
rect 8116 23672 8168 23724
rect 8392 23715 8444 23724
rect 8392 23681 8401 23715
rect 8401 23681 8435 23715
rect 8435 23681 8444 23715
rect 8392 23672 8444 23681
rect 15844 23740 15896 23792
rect 16028 23740 16080 23792
rect 21272 23740 21324 23792
rect 9680 23672 9732 23724
rect 11152 23672 11204 23724
rect 14464 23672 14516 23724
rect 18052 23672 18104 23724
rect 8668 23604 8720 23656
rect 8208 23536 8260 23588
rect 9312 23536 9364 23588
rect 22836 23672 22888 23724
rect 21364 23604 21416 23656
rect 24032 23740 24084 23792
rect 23296 23672 23348 23724
rect 23756 23715 23808 23724
rect 23756 23681 23765 23715
rect 23765 23681 23799 23715
rect 23799 23681 23808 23715
rect 23756 23672 23808 23681
rect 24952 23672 25004 23724
rect 25688 23808 25740 23860
rect 26608 23808 26660 23860
rect 26792 23740 26844 23792
rect 27160 23783 27212 23792
rect 27160 23749 27169 23783
rect 27169 23749 27203 23783
rect 27203 23749 27212 23783
rect 27160 23740 27212 23749
rect 27712 23808 27764 23860
rect 26332 23672 26384 23724
rect 26976 23672 27028 23724
rect 27344 23715 27396 23724
rect 27344 23681 27353 23715
rect 27353 23681 27387 23715
rect 27387 23681 27396 23715
rect 27896 23740 27948 23792
rect 27344 23672 27396 23681
rect 28816 23808 28868 23860
rect 29460 23808 29512 23860
rect 31300 23808 31352 23860
rect 31944 23808 31996 23860
rect 33048 23808 33100 23860
rect 33140 23808 33192 23860
rect 28632 23783 28684 23792
rect 28632 23749 28641 23783
rect 28641 23749 28675 23783
rect 28675 23749 28684 23783
rect 28632 23740 28684 23749
rect 31392 23740 31444 23792
rect 32128 23740 32180 23792
rect 32772 23740 32824 23792
rect 29920 23715 29972 23724
rect 23664 23579 23716 23588
rect 23664 23545 23673 23579
rect 23673 23545 23707 23579
rect 23707 23545 23716 23579
rect 23664 23536 23716 23545
rect 27068 23604 27120 23656
rect 29920 23681 29929 23715
rect 29929 23681 29963 23715
rect 29963 23681 29972 23715
rect 29920 23672 29972 23681
rect 32588 23715 32640 23724
rect 29644 23604 29696 23656
rect 29828 23604 29880 23656
rect 32588 23681 32597 23715
rect 32597 23681 32631 23715
rect 32631 23681 32640 23715
rect 32588 23672 32640 23681
rect 34428 23740 34480 23792
rect 37740 23808 37792 23860
rect 37832 23808 37884 23860
rect 34796 23715 34848 23724
rect 30656 23604 30708 23656
rect 34796 23681 34805 23715
rect 34805 23681 34839 23715
rect 34839 23681 34848 23715
rect 34796 23672 34848 23681
rect 34888 23715 34940 23724
rect 34888 23681 34898 23715
rect 34898 23681 34932 23715
rect 34932 23681 34940 23715
rect 35256 23715 35308 23724
rect 34888 23672 34940 23681
rect 35256 23681 35270 23715
rect 35270 23681 35304 23715
rect 35304 23681 35308 23715
rect 35256 23672 35308 23681
rect 27896 23536 27948 23588
rect 30012 23579 30064 23588
rect 4620 23468 4672 23520
rect 5356 23468 5408 23520
rect 5908 23511 5960 23520
rect 5908 23477 5917 23511
rect 5917 23477 5951 23511
rect 5951 23477 5960 23511
rect 5908 23468 5960 23477
rect 6920 23511 6972 23520
rect 6920 23477 6929 23511
rect 6929 23477 6963 23511
rect 6963 23477 6972 23511
rect 6920 23468 6972 23477
rect 8576 23468 8628 23520
rect 10600 23511 10652 23520
rect 10600 23477 10609 23511
rect 10609 23477 10643 23511
rect 10643 23477 10652 23511
rect 10600 23468 10652 23477
rect 10692 23468 10744 23520
rect 12440 23468 12492 23520
rect 16304 23468 16356 23520
rect 16488 23468 16540 23520
rect 19892 23468 19944 23520
rect 20076 23511 20128 23520
rect 20076 23477 20085 23511
rect 20085 23477 20119 23511
rect 20119 23477 20128 23511
rect 20076 23468 20128 23477
rect 20536 23468 20588 23520
rect 26240 23468 26292 23520
rect 28356 23468 28408 23520
rect 28632 23468 28684 23520
rect 30012 23545 30021 23579
rect 30021 23545 30055 23579
rect 30055 23545 30064 23579
rect 30012 23536 30064 23545
rect 36176 23715 36228 23724
rect 36176 23681 36185 23715
rect 36185 23681 36219 23715
rect 36219 23681 36228 23715
rect 36176 23672 36228 23681
rect 36544 23604 36596 23656
rect 28954 23468 29006 23520
rect 32956 23468 33008 23520
rect 35624 23536 35676 23588
rect 36268 23536 36320 23588
rect 37740 23672 37792 23724
rect 38016 23647 38068 23656
rect 38016 23613 38025 23647
rect 38025 23613 38059 23647
rect 38059 23613 38068 23647
rect 38016 23604 38068 23613
rect 37924 23536 37976 23588
rect 37004 23468 37056 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 3976 23307 4028 23316
rect 3976 23273 3985 23307
rect 3985 23273 4019 23307
rect 4019 23273 4028 23307
rect 3976 23264 4028 23273
rect 5908 23264 5960 23316
rect 6920 23239 6972 23248
rect 6920 23205 6929 23239
rect 6929 23205 6963 23239
rect 6963 23205 6972 23239
rect 6920 23196 6972 23205
rect 4804 23128 4856 23180
rect 6000 23128 6052 23180
rect 7196 23128 7248 23180
rect 4160 23060 4212 23112
rect 4620 23060 4672 23112
rect 4896 23060 4948 23112
rect 6644 23060 6696 23112
rect 6736 23103 6788 23112
rect 6736 23069 6745 23103
rect 6745 23069 6779 23103
rect 6779 23069 6788 23103
rect 6736 23060 6788 23069
rect 6920 23060 6972 23112
rect 10692 23264 10744 23316
rect 15660 23264 15712 23316
rect 20720 23264 20772 23316
rect 21272 23307 21324 23316
rect 21272 23273 21281 23307
rect 21281 23273 21315 23307
rect 21315 23273 21324 23307
rect 21272 23264 21324 23273
rect 22560 23307 22612 23316
rect 22560 23273 22569 23307
rect 22569 23273 22603 23307
rect 22603 23273 22612 23307
rect 22560 23264 22612 23273
rect 36176 23264 36228 23316
rect 37740 23264 37792 23316
rect 15200 23196 15252 23248
rect 14280 23128 14332 23180
rect 8668 23060 8720 23112
rect 9128 23103 9180 23112
rect 9128 23069 9137 23103
rect 9137 23069 9171 23103
rect 9171 23069 9180 23103
rect 9128 23060 9180 23069
rect 7196 22924 7248 22976
rect 7564 22967 7616 22976
rect 7564 22933 7573 22967
rect 7573 22933 7607 22967
rect 7607 22933 7616 22967
rect 7564 22924 7616 22933
rect 8944 22992 8996 23044
rect 12348 23035 12400 23044
rect 12348 23001 12382 23035
rect 12382 23001 12400 23035
rect 12348 22992 12400 23001
rect 9864 22924 9916 22976
rect 12072 22924 12124 22976
rect 15384 23060 15436 23112
rect 15660 23060 15712 23112
rect 15752 23060 15804 23112
rect 18420 23060 18472 23112
rect 16028 22924 16080 22976
rect 17224 23035 17276 23044
rect 17224 23001 17258 23035
rect 17258 23001 17276 23035
rect 31944 23196 31996 23248
rect 32956 23196 33008 23248
rect 36544 23196 36596 23248
rect 20536 23171 20588 23180
rect 20536 23137 20545 23171
rect 20545 23137 20579 23171
rect 20579 23137 20588 23171
rect 20536 23128 20588 23137
rect 20628 23171 20680 23180
rect 20628 23137 20637 23171
rect 20637 23137 20671 23171
rect 20671 23137 20680 23171
rect 20628 23128 20680 23137
rect 20904 23128 20956 23180
rect 20996 23128 21048 23180
rect 18972 23060 19024 23112
rect 23204 23128 23256 23180
rect 25412 23128 25464 23180
rect 17224 22992 17276 23001
rect 18328 22967 18380 22976
rect 18328 22933 18337 22967
rect 18337 22933 18371 22967
rect 18371 22933 18380 22967
rect 18328 22924 18380 22933
rect 24768 23060 24820 23112
rect 26240 23060 26292 23112
rect 27344 23128 27396 23180
rect 27896 23128 27948 23180
rect 29644 23128 29696 23180
rect 29920 23128 29972 23180
rect 26792 23060 26844 23112
rect 27712 23060 27764 23112
rect 27988 23103 28040 23112
rect 27988 23069 27997 23103
rect 27997 23069 28031 23103
rect 28031 23069 28040 23103
rect 27988 23060 28040 23069
rect 28632 23103 28684 23112
rect 28632 23069 28639 23103
rect 28639 23069 28684 23103
rect 28632 23060 28684 23069
rect 28724 23103 28776 23112
rect 28724 23069 28733 23103
rect 28733 23069 28767 23103
rect 28767 23069 28776 23103
rect 28724 23060 28776 23069
rect 28908 23103 28960 23112
rect 28908 23069 28922 23103
rect 28922 23069 28956 23103
rect 28956 23069 28960 23103
rect 28908 23060 28960 23069
rect 29276 23060 29328 23112
rect 29828 23103 29880 23112
rect 29828 23069 29837 23103
rect 29837 23069 29871 23103
rect 29871 23069 29880 23103
rect 29828 23060 29880 23069
rect 30012 23060 30064 23112
rect 31300 23128 31352 23180
rect 35808 23128 35860 23180
rect 34520 23060 34572 23112
rect 35532 23103 35584 23112
rect 31852 22992 31904 23044
rect 20444 22967 20496 22976
rect 20444 22933 20453 22967
rect 20453 22933 20487 22967
rect 20487 22933 20496 22967
rect 20444 22924 20496 22933
rect 21640 22967 21692 22976
rect 21640 22933 21649 22967
rect 21649 22933 21683 22967
rect 21683 22933 21692 22967
rect 21640 22924 21692 22933
rect 24492 22924 24544 22976
rect 29460 22924 29512 22976
rect 29920 22924 29972 22976
rect 30932 22967 30984 22976
rect 30932 22933 30941 22967
rect 30941 22933 30975 22967
rect 30975 22933 30984 22967
rect 35532 23069 35541 23103
rect 35541 23069 35575 23103
rect 35575 23069 35584 23103
rect 35532 23060 35584 23069
rect 36820 23060 36872 23112
rect 37004 23103 37056 23112
rect 37004 23069 37038 23103
rect 37038 23069 37056 23103
rect 37004 23060 37056 23069
rect 30932 22924 30984 22933
rect 35440 22924 35492 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 4712 22720 4764 22772
rect 6644 22720 6696 22772
rect 7104 22720 7156 22772
rect 8944 22763 8996 22772
rect 8944 22729 8953 22763
rect 8953 22729 8987 22763
rect 8987 22729 8996 22763
rect 8944 22720 8996 22729
rect 12348 22763 12400 22772
rect 12348 22729 12357 22763
rect 12357 22729 12391 22763
rect 12391 22729 12400 22763
rect 12348 22720 12400 22729
rect 15660 22763 15712 22772
rect 15660 22729 15669 22763
rect 15669 22729 15703 22763
rect 15703 22729 15712 22763
rect 15660 22720 15712 22729
rect 5080 22652 5132 22704
rect 7840 22652 7892 22704
rect 10416 22652 10468 22704
rect 4896 22627 4948 22636
rect 4896 22593 4905 22627
rect 4905 22593 4939 22627
rect 4939 22593 4948 22627
rect 4896 22584 4948 22593
rect 7472 22627 7524 22636
rect 7472 22593 7481 22627
rect 7481 22593 7515 22627
rect 7515 22593 7524 22627
rect 7472 22584 7524 22593
rect 8668 22584 8720 22636
rect 10600 22584 10652 22636
rect 11704 22652 11756 22704
rect 12072 22695 12124 22704
rect 12072 22661 12081 22695
rect 12081 22661 12115 22695
rect 12115 22661 12124 22695
rect 12072 22652 12124 22661
rect 14280 22652 14332 22704
rect 11152 22627 11204 22636
rect 7288 22559 7340 22568
rect 7288 22525 7297 22559
rect 7297 22525 7331 22559
rect 7331 22525 7340 22559
rect 7288 22516 7340 22525
rect 8024 22516 8076 22568
rect 9312 22559 9364 22568
rect 9312 22525 9321 22559
rect 9321 22525 9355 22559
rect 9355 22525 9364 22559
rect 11152 22593 11161 22627
rect 11161 22593 11195 22627
rect 11195 22593 11204 22627
rect 11152 22584 11204 22593
rect 11796 22627 11848 22636
rect 11796 22593 11805 22627
rect 11805 22593 11839 22627
rect 11839 22593 11848 22627
rect 11796 22584 11848 22593
rect 12256 22584 12308 22636
rect 14372 22627 14424 22636
rect 14372 22593 14381 22627
rect 14381 22593 14415 22627
rect 14415 22593 14424 22627
rect 14372 22584 14424 22593
rect 14556 22627 14608 22636
rect 14556 22593 14565 22627
rect 14565 22593 14599 22627
rect 14599 22593 14608 22627
rect 14556 22584 14608 22593
rect 15292 22652 15344 22704
rect 16856 22695 16908 22704
rect 15108 22584 15160 22636
rect 9312 22516 9364 22525
rect 5908 22448 5960 22500
rect 15292 22448 15344 22500
rect 7196 22423 7248 22432
rect 7196 22389 7205 22423
rect 7205 22389 7239 22423
rect 7239 22389 7248 22423
rect 7196 22380 7248 22389
rect 8116 22380 8168 22432
rect 10600 22380 10652 22432
rect 14464 22423 14516 22432
rect 14464 22389 14473 22423
rect 14473 22389 14507 22423
rect 14507 22389 14516 22423
rect 14464 22380 14516 22389
rect 15476 22380 15528 22432
rect 16029 22627 16081 22636
rect 16029 22593 16038 22627
rect 16038 22593 16072 22627
rect 16072 22593 16081 22627
rect 16856 22661 16865 22695
rect 16865 22661 16899 22695
rect 16899 22661 16908 22695
rect 21088 22720 21140 22772
rect 21640 22720 21692 22772
rect 16856 22652 16908 22661
rect 20076 22695 20128 22704
rect 16029 22584 16081 22593
rect 16580 22584 16632 22636
rect 17132 22584 17184 22636
rect 17500 22584 17552 22636
rect 18328 22627 18380 22636
rect 18328 22593 18337 22627
rect 18337 22593 18371 22627
rect 18371 22593 18380 22627
rect 18328 22584 18380 22593
rect 18420 22584 18472 22636
rect 20076 22661 20110 22695
rect 20110 22661 20128 22695
rect 20076 22652 20128 22661
rect 21824 22652 21876 22704
rect 21548 22584 21600 22636
rect 22652 22627 22704 22636
rect 22652 22593 22661 22627
rect 22661 22593 22695 22627
rect 22695 22593 22704 22627
rect 22652 22584 22704 22593
rect 22928 22627 22980 22636
rect 22928 22593 22937 22627
rect 22937 22593 22971 22627
rect 22971 22593 22980 22627
rect 22928 22584 22980 22593
rect 23664 22584 23716 22636
rect 16488 22516 16540 22568
rect 17408 22559 17460 22568
rect 17408 22525 17417 22559
rect 17417 22525 17451 22559
rect 17451 22525 17460 22559
rect 17408 22516 17460 22525
rect 18512 22559 18564 22568
rect 18512 22525 18521 22559
rect 18521 22525 18555 22559
rect 18555 22525 18564 22559
rect 18512 22516 18564 22525
rect 23388 22559 23440 22568
rect 23388 22525 23397 22559
rect 23397 22525 23431 22559
rect 23431 22525 23440 22559
rect 23388 22516 23440 22525
rect 24400 22652 24452 22704
rect 24492 22627 24544 22636
rect 24492 22593 24501 22627
rect 24501 22593 24535 22627
rect 24535 22593 24544 22627
rect 24492 22584 24544 22593
rect 25320 22652 25372 22704
rect 26424 22652 26476 22704
rect 25596 22584 25648 22636
rect 16212 22448 16264 22500
rect 19800 22448 19852 22500
rect 16856 22380 16908 22432
rect 20168 22380 20220 22432
rect 25780 22516 25832 22568
rect 26148 22516 26200 22568
rect 27620 22720 27672 22772
rect 28540 22720 28592 22772
rect 29828 22720 29880 22772
rect 30104 22720 30156 22772
rect 30748 22720 30800 22772
rect 27344 22652 27396 22704
rect 30840 22652 30892 22704
rect 33692 22720 33744 22772
rect 32496 22652 32548 22704
rect 35808 22695 35860 22704
rect 35808 22661 35817 22695
rect 35817 22661 35851 22695
rect 35851 22661 35860 22695
rect 35808 22652 35860 22661
rect 27620 22627 27672 22636
rect 27620 22593 27629 22627
rect 27629 22593 27663 22627
rect 27663 22593 27672 22627
rect 27620 22584 27672 22593
rect 27712 22627 27764 22636
rect 27712 22593 27722 22627
rect 27722 22593 27756 22627
rect 27756 22593 27764 22627
rect 27896 22627 27948 22636
rect 27712 22584 27764 22593
rect 27896 22593 27905 22627
rect 27905 22593 27939 22627
rect 27939 22593 27948 22627
rect 27896 22584 27948 22593
rect 28264 22584 28316 22636
rect 28908 22584 28960 22636
rect 29368 22627 29420 22636
rect 29368 22593 29377 22627
rect 29377 22593 29411 22627
rect 29411 22593 29420 22627
rect 29368 22584 29420 22593
rect 29736 22627 29788 22636
rect 29736 22593 29745 22627
rect 29745 22593 29779 22627
rect 29779 22593 29788 22627
rect 29736 22584 29788 22593
rect 30472 22584 30524 22636
rect 31208 22627 31260 22636
rect 31208 22593 31217 22627
rect 31217 22593 31251 22627
rect 31251 22593 31260 22627
rect 31208 22584 31260 22593
rect 31576 22627 31628 22636
rect 31576 22593 31585 22627
rect 31585 22593 31619 22627
rect 31619 22593 31628 22627
rect 31576 22584 31628 22593
rect 33140 22627 33192 22636
rect 33140 22593 33149 22627
rect 33149 22593 33183 22627
rect 33183 22593 33192 22627
rect 33140 22584 33192 22593
rect 33968 22584 34020 22636
rect 35440 22627 35492 22636
rect 35440 22593 35449 22627
rect 35449 22593 35483 22627
rect 35483 22593 35492 22627
rect 35440 22584 35492 22593
rect 35532 22584 35584 22636
rect 35716 22627 35768 22636
rect 35716 22593 35725 22627
rect 35725 22593 35759 22627
rect 35759 22593 35768 22627
rect 35716 22584 35768 22593
rect 37740 22584 37792 22636
rect 29460 22516 29512 22568
rect 30748 22559 30800 22568
rect 30748 22525 30757 22559
rect 30757 22525 30791 22559
rect 30791 22525 30800 22559
rect 30748 22516 30800 22525
rect 34612 22516 34664 22568
rect 38108 22559 38160 22568
rect 38108 22525 38117 22559
rect 38117 22525 38151 22559
rect 38151 22525 38160 22559
rect 38108 22516 38160 22525
rect 31484 22448 31536 22500
rect 29000 22380 29052 22432
rect 36360 22380 36412 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 7472 22176 7524 22228
rect 11704 22176 11756 22228
rect 11888 22219 11940 22228
rect 11888 22185 11897 22219
rect 11897 22185 11931 22219
rect 11931 22185 11940 22219
rect 11888 22176 11940 22185
rect 14372 22176 14424 22228
rect 16488 22176 16540 22228
rect 19800 22176 19852 22228
rect 20444 22176 20496 22228
rect 20720 22176 20772 22228
rect 21824 22176 21876 22228
rect 9312 22108 9364 22160
rect 4620 22083 4672 22092
rect 4620 22049 4629 22083
rect 4629 22049 4663 22083
rect 4663 22049 4672 22083
rect 4620 22040 4672 22049
rect 4712 21972 4764 22024
rect 7104 21972 7156 22024
rect 7472 22015 7524 22024
rect 7472 21981 7481 22015
rect 7481 21981 7515 22015
rect 7515 21981 7524 22015
rect 7472 21972 7524 21981
rect 7840 22015 7892 22024
rect 6736 21904 6788 21956
rect 7196 21904 7248 21956
rect 7840 21981 7849 22015
rect 7849 21981 7883 22015
rect 7883 21981 7892 22015
rect 7840 21972 7892 21981
rect 7932 21972 7984 22024
rect 8392 21972 8444 22024
rect 9220 22015 9272 22024
rect 9220 21981 9229 22015
rect 9229 21981 9263 22015
rect 9263 21981 9272 22015
rect 9220 21972 9272 21981
rect 12164 21972 12216 22024
rect 15200 22040 15252 22092
rect 14464 22015 14516 22024
rect 14464 21981 14473 22015
rect 14473 21981 14507 22015
rect 14507 21981 14516 22015
rect 14464 21972 14516 21981
rect 15384 22040 15436 22092
rect 15936 22108 15988 22160
rect 17408 22108 17460 22160
rect 22192 22176 22244 22228
rect 22468 22176 22520 22228
rect 27620 22176 27672 22228
rect 31208 22176 31260 22228
rect 33048 22176 33100 22228
rect 24308 22108 24360 22160
rect 16580 22040 16632 22092
rect 23020 22083 23072 22092
rect 23020 22049 23029 22083
rect 23029 22049 23063 22083
rect 23063 22049 23072 22083
rect 23020 22040 23072 22049
rect 26056 22108 26108 22160
rect 27712 22108 27764 22160
rect 25780 22083 25832 22092
rect 15476 22015 15528 22024
rect 15476 21981 15485 22015
rect 15485 21981 15519 22015
rect 15519 21981 15528 22015
rect 15476 21972 15528 21981
rect 16212 22015 16264 22024
rect 16212 21981 16221 22015
rect 16221 21981 16255 22015
rect 16255 21981 16264 22015
rect 16212 21972 16264 21981
rect 16764 21972 16816 22024
rect 22928 22015 22980 22024
rect 22928 21981 22937 22015
rect 22937 21981 22971 22015
rect 22971 21981 22980 22015
rect 22928 21972 22980 21981
rect 24124 21972 24176 22024
rect 24952 21972 25004 22024
rect 25136 21972 25188 22024
rect 25228 21972 25280 22024
rect 25780 22049 25789 22083
rect 25789 22049 25823 22083
rect 25823 22049 25832 22083
rect 25780 22040 25832 22049
rect 28540 22040 28592 22092
rect 28816 22040 28868 22092
rect 29460 22040 29512 22092
rect 31760 22108 31812 22160
rect 31300 22083 31352 22092
rect 31300 22049 31309 22083
rect 31309 22049 31343 22083
rect 31343 22049 31352 22083
rect 31300 22040 31352 22049
rect 26792 22015 26844 22024
rect 26792 21981 26801 22015
rect 26801 21981 26835 22015
rect 26835 21981 26844 22015
rect 26792 21972 26844 21981
rect 27712 21972 27764 22024
rect 27896 22015 27948 22024
rect 27896 21981 27905 22015
rect 27905 21981 27939 22015
rect 27939 21981 27948 22015
rect 27896 21972 27948 21981
rect 27988 21972 28040 22024
rect 28356 21972 28408 22024
rect 28448 21972 28500 22024
rect 30932 22015 30984 22024
rect 30932 21981 30941 22015
rect 30941 21981 30975 22015
rect 30975 21981 30984 22015
rect 30932 21972 30984 21981
rect 31116 21972 31168 22024
rect 32496 21972 32548 22024
rect 32680 22108 32732 22160
rect 33140 22108 33192 22160
rect 35532 22176 35584 22228
rect 33692 22040 33744 22092
rect 33048 22015 33100 22024
rect 33048 21981 33062 22015
rect 33062 21981 33096 22015
rect 33096 21981 33100 22015
rect 33048 21972 33100 21981
rect 33968 21972 34020 22024
rect 9680 21904 9732 21956
rect 10048 21904 10100 21956
rect 10600 21904 10652 21956
rect 3976 21879 4028 21888
rect 3976 21845 3985 21879
rect 3985 21845 4019 21879
rect 4019 21845 4028 21879
rect 3976 21836 4028 21845
rect 4344 21879 4396 21888
rect 4344 21845 4353 21879
rect 4353 21845 4387 21879
rect 4387 21845 4396 21879
rect 4344 21836 4396 21845
rect 6644 21836 6696 21888
rect 7564 21836 7616 21888
rect 8576 21836 8628 21888
rect 14648 21947 14700 21956
rect 14648 21913 14657 21947
rect 14657 21913 14691 21947
rect 14691 21913 14700 21947
rect 14648 21904 14700 21913
rect 13728 21879 13780 21888
rect 13728 21845 13737 21879
rect 13737 21845 13771 21879
rect 13771 21845 13780 21879
rect 13728 21836 13780 21845
rect 15936 21904 15988 21956
rect 17224 21904 17276 21956
rect 26700 21904 26752 21956
rect 16028 21836 16080 21888
rect 16580 21879 16632 21888
rect 16580 21845 16589 21879
rect 16589 21845 16623 21879
rect 16623 21845 16632 21879
rect 16580 21836 16632 21845
rect 24676 21836 24728 21888
rect 24952 21836 25004 21888
rect 25780 21836 25832 21888
rect 27068 21947 27120 21956
rect 27068 21913 27077 21947
rect 27077 21913 27111 21947
rect 27111 21913 27120 21947
rect 27068 21904 27120 21913
rect 32128 21904 32180 21956
rect 32864 21947 32916 21956
rect 32864 21913 32873 21947
rect 32873 21913 32907 21947
rect 32907 21913 32916 21947
rect 32864 21904 32916 21913
rect 36820 21972 36872 22024
rect 27252 21836 27304 21888
rect 27528 21836 27580 21888
rect 27988 21836 28040 21888
rect 28632 21836 28684 21888
rect 30656 21879 30708 21888
rect 30656 21845 30665 21879
rect 30665 21845 30699 21879
rect 30699 21845 30708 21879
rect 30656 21836 30708 21845
rect 31392 21836 31444 21888
rect 31760 21836 31812 21888
rect 32220 21836 32272 21888
rect 37464 21904 37516 21956
rect 33232 21879 33284 21888
rect 33232 21845 33241 21879
rect 33241 21845 33275 21879
rect 33275 21845 33284 21879
rect 33232 21836 33284 21845
rect 35532 21836 35584 21888
rect 36636 21836 36688 21888
rect 38292 21879 38344 21888
rect 38292 21845 38301 21879
rect 38301 21845 38335 21879
rect 38335 21845 38344 21879
rect 38292 21836 38344 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 5908 21632 5960 21684
rect 3976 21564 4028 21616
rect 2780 21539 2832 21548
rect 2780 21505 2789 21539
rect 2789 21505 2823 21539
rect 2823 21505 2832 21539
rect 2780 21496 2832 21505
rect 5816 21496 5868 21548
rect 6644 21564 6696 21616
rect 7472 21632 7524 21684
rect 9404 21632 9456 21684
rect 12440 21632 12492 21684
rect 6736 21539 6788 21548
rect 6736 21505 6745 21539
rect 6745 21505 6779 21539
rect 6779 21505 6788 21539
rect 6736 21496 6788 21505
rect 6920 21539 6972 21548
rect 6920 21505 6929 21539
rect 6929 21505 6963 21539
rect 6963 21505 6972 21539
rect 6920 21496 6972 21505
rect 8208 21496 8260 21548
rect 4620 21428 4672 21480
rect 7932 21471 7984 21480
rect 7932 21437 7941 21471
rect 7941 21437 7975 21471
rect 7975 21437 7984 21471
rect 7932 21428 7984 21437
rect 4344 21360 4396 21412
rect 6000 21292 6052 21344
rect 7656 21335 7708 21344
rect 7656 21301 7665 21335
rect 7665 21301 7699 21335
rect 7699 21301 7708 21335
rect 7656 21292 7708 21301
rect 7840 21360 7892 21412
rect 8116 21471 8168 21480
rect 8116 21437 8125 21471
rect 8125 21437 8159 21471
rect 8159 21437 8168 21471
rect 8116 21428 8168 21437
rect 11888 21564 11940 21616
rect 15752 21564 15804 21616
rect 9772 21496 9824 21548
rect 13820 21496 13872 21548
rect 15660 21496 15712 21548
rect 9220 21428 9272 21480
rect 11888 21428 11940 21480
rect 14556 21428 14608 21480
rect 14924 21471 14976 21480
rect 14924 21437 14933 21471
rect 14933 21437 14967 21471
rect 14967 21437 14976 21471
rect 14924 21428 14976 21437
rect 16948 21564 17000 21616
rect 16672 21496 16724 21548
rect 19432 21496 19484 21548
rect 16212 21471 16264 21480
rect 16212 21437 16221 21471
rect 16221 21437 16255 21471
rect 16255 21437 16264 21471
rect 16212 21428 16264 21437
rect 18420 21428 18472 21480
rect 22100 21632 22152 21684
rect 24584 21632 24636 21684
rect 26884 21632 26936 21684
rect 27252 21632 27304 21684
rect 27068 21564 27120 21616
rect 27436 21607 27488 21616
rect 27436 21573 27445 21607
rect 27445 21573 27479 21607
rect 27479 21573 27488 21607
rect 27436 21564 27488 21573
rect 22192 21539 22244 21548
rect 22192 21505 22201 21539
rect 22201 21505 22235 21539
rect 22235 21505 22244 21539
rect 22192 21496 22244 21505
rect 22376 21539 22428 21548
rect 22376 21505 22390 21539
rect 22390 21505 22424 21539
rect 22424 21505 22428 21539
rect 22376 21496 22428 21505
rect 24676 21496 24728 21548
rect 26332 21539 26384 21548
rect 26332 21505 26341 21539
rect 26341 21505 26375 21539
rect 26375 21505 26384 21539
rect 26332 21496 26384 21505
rect 26608 21539 26660 21548
rect 26608 21505 26617 21539
rect 26617 21505 26651 21539
rect 26651 21505 26660 21539
rect 26608 21496 26660 21505
rect 26700 21496 26752 21548
rect 27620 21564 27672 21616
rect 28632 21607 28684 21616
rect 28632 21573 28641 21607
rect 28641 21573 28675 21607
rect 28675 21573 28684 21607
rect 28632 21564 28684 21573
rect 28540 21539 28592 21548
rect 28540 21505 28547 21539
rect 28547 21505 28592 21539
rect 9220 21335 9272 21344
rect 9220 21301 9229 21335
rect 9229 21301 9263 21335
rect 9263 21301 9272 21335
rect 9220 21292 9272 21301
rect 9588 21292 9640 21344
rect 10968 21360 11020 21412
rect 13544 21360 13596 21412
rect 13636 21360 13688 21412
rect 21824 21360 21876 21412
rect 27252 21428 27304 21480
rect 28540 21496 28592 21505
rect 35532 21632 35584 21684
rect 37464 21675 37516 21684
rect 32496 21564 32548 21616
rect 33232 21564 33284 21616
rect 33692 21564 33744 21616
rect 30472 21539 30524 21548
rect 24584 21360 24636 21412
rect 14280 21292 14332 21344
rect 14740 21335 14792 21344
rect 14740 21301 14749 21335
rect 14749 21301 14783 21335
rect 14783 21301 14792 21335
rect 14740 21292 14792 21301
rect 15200 21335 15252 21344
rect 15200 21301 15209 21335
rect 15209 21301 15243 21335
rect 15243 21301 15252 21335
rect 15200 21292 15252 21301
rect 15384 21292 15436 21344
rect 15844 21292 15896 21344
rect 19340 21292 19392 21344
rect 25136 21292 25188 21344
rect 27436 21292 27488 21344
rect 27804 21292 27856 21344
rect 30472 21505 30481 21539
rect 30481 21505 30515 21539
rect 30515 21505 30524 21539
rect 30472 21496 30524 21505
rect 30748 21539 30800 21548
rect 30748 21505 30757 21539
rect 30757 21505 30791 21539
rect 30791 21505 30800 21539
rect 30748 21496 30800 21505
rect 31208 21539 31260 21548
rect 31208 21505 31217 21539
rect 31217 21505 31251 21539
rect 31251 21505 31260 21539
rect 31208 21496 31260 21505
rect 31484 21496 31536 21548
rect 32588 21496 32640 21548
rect 32956 21539 33008 21548
rect 32956 21505 32965 21539
rect 32965 21505 32999 21539
rect 32999 21505 33008 21539
rect 32956 21496 33008 21505
rect 34796 21496 34848 21548
rect 35256 21539 35308 21548
rect 30564 21428 30616 21480
rect 34428 21428 34480 21480
rect 34520 21428 34572 21480
rect 35256 21505 35265 21539
rect 35265 21505 35299 21539
rect 35299 21505 35308 21539
rect 35256 21496 35308 21505
rect 35532 21496 35584 21548
rect 37464 21641 37473 21675
rect 37473 21641 37507 21675
rect 37507 21641 37516 21675
rect 37464 21632 37516 21641
rect 37740 21564 37792 21616
rect 36360 21539 36412 21548
rect 36360 21505 36369 21539
rect 36369 21505 36403 21539
rect 36403 21505 36412 21539
rect 36636 21539 36688 21548
rect 36360 21496 36412 21505
rect 36636 21505 36645 21539
rect 36645 21505 36679 21539
rect 36679 21505 36688 21539
rect 36636 21496 36688 21505
rect 38292 21496 38344 21548
rect 38016 21471 38068 21480
rect 29092 21360 29144 21412
rect 31300 21360 31352 21412
rect 33140 21360 33192 21412
rect 38016 21437 38025 21471
rect 38025 21437 38059 21471
rect 38059 21437 38068 21471
rect 38016 21428 38068 21437
rect 35348 21360 35400 21412
rect 36544 21403 36596 21412
rect 36544 21369 36553 21403
rect 36553 21369 36587 21403
rect 36587 21369 36596 21403
rect 36544 21360 36596 21369
rect 29736 21292 29788 21344
rect 34428 21292 34480 21344
rect 35256 21292 35308 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 5908 21131 5960 21140
rect 5908 21097 5917 21131
rect 5917 21097 5951 21131
rect 5951 21097 5960 21131
rect 5908 21088 5960 21097
rect 9588 21088 9640 21140
rect 10692 21088 10744 21140
rect 10968 21131 11020 21140
rect 10968 21097 10977 21131
rect 10977 21097 11011 21131
rect 11011 21097 11020 21131
rect 10968 21088 11020 21097
rect 14556 21088 14608 21140
rect 15844 21088 15896 21140
rect 18512 21131 18564 21140
rect 18512 21097 18521 21131
rect 18521 21097 18555 21131
rect 18555 21097 18564 21131
rect 18512 21088 18564 21097
rect 21824 21131 21876 21140
rect 21824 21097 21833 21131
rect 21833 21097 21867 21131
rect 21867 21097 21876 21131
rect 21824 21088 21876 21097
rect 25044 21088 25096 21140
rect 25320 21088 25372 21140
rect 25688 21088 25740 21140
rect 26332 21088 26384 21140
rect 30472 21088 30524 21140
rect 31392 21088 31444 21140
rect 31944 21131 31996 21140
rect 31944 21097 31953 21131
rect 31953 21097 31987 21131
rect 31987 21097 31996 21131
rect 31944 21088 31996 21097
rect 13728 21020 13780 21072
rect 2780 20952 2832 21004
rect 3976 20952 4028 21004
rect 9220 20952 9272 21004
rect 15292 20952 15344 21004
rect 6000 20884 6052 20936
rect 7012 20884 7064 20936
rect 7196 20884 7248 20936
rect 9128 20884 9180 20936
rect 13544 20884 13596 20936
rect 16764 20952 16816 21004
rect 28908 21020 28960 21072
rect 30196 21020 30248 21072
rect 33600 21020 33652 21072
rect 24124 20952 24176 21004
rect 15568 20884 15620 20936
rect 17592 20927 17644 20936
rect 9956 20816 10008 20868
rect 13912 20816 13964 20868
rect 14464 20816 14516 20868
rect 17592 20893 17601 20927
rect 17601 20893 17635 20927
rect 17635 20893 17644 20927
rect 17592 20884 17644 20893
rect 20536 20927 20588 20936
rect 20536 20893 20545 20927
rect 20545 20893 20579 20927
rect 20579 20893 20588 20927
rect 20536 20884 20588 20893
rect 24492 20884 24544 20936
rect 24768 20952 24820 21004
rect 25320 20927 25372 20936
rect 15752 20859 15804 20868
rect 15752 20825 15761 20859
rect 15761 20825 15795 20859
rect 15795 20825 15804 20859
rect 15752 20816 15804 20825
rect 15936 20816 15988 20868
rect 17224 20859 17276 20868
rect 17224 20825 17233 20859
rect 17233 20825 17267 20859
rect 17267 20825 17276 20859
rect 17224 20816 17276 20825
rect 17868 20816 17920 20868
rect 17960 20859 18012 20868
rect 17960 20825 17969 20859
rect 17969 20825 18003 20859
rect 18003 20825 18012 20859
rect 17960 20816 18012 20825
rect 25320 20893 25329 20927
rect 25329 20893 25363 20927
rect 25363 20893 25372 20927
rect 25320 20884 25372 20893
rect 25412 20884 25464 20936
rect 26056 20884 26108 20936
rect 27252 20927 27304 20936
rect 27252 20893 27261 20927
rect 27261 20893 27295 20927
rect 27295 20893 27304 20927
rect 27252 20884 27304 20893
rect 27528 20927 27580 20936
rect 27528 20893 27537 20927
rect 27537 20893 27571 20927
rect 27571 20893 27580 20927
rect 27528 20884 27580 20893
rect 27620 20927 27672 20936
rect 27620 20893 27629 20927
rect 27629 20893 27663 20927
rect 27663 20893 27672 20927
rect 27620 20884 27672 20893
rect 27896 20884 27948 20936
rect 29920 20927 29972 20936
rect 29920 20893 29929 20927
rect 29929 20893 29963 20927
rect 29963 20893 29972 20927
rect 29920 20884 29972 20893
rect 26148 20859 26200 20868
rect 6552 20748 6604 20800
rect 7104 20748 7156 20800
rect 14280 20791 14332 20800
rect 14280 20757 14289 20791
rect 14289 20757 14323 20791
rect 14323 20757 14332 20791
rect 14280 20748 14332 20757
rect 14740 20791 14792 20800
rect 14740 20757 14749 20791
rect 14749 20757 14783 20791
rect 14783 20757 14792 20791
rect 14740 20748 14792 20757
rect 15200 20748 15252 20800
rect 15660 20748 15712 20800
rect 26148 20825 26157 20859
rect 26157 20825 26191 20859
rect 26191 20825 26200 20859
rect 26148 20816 26200 20825
rect 20076 20748 20128 20800
rect 20996 20748 21048 20800
rect 24768 20748 24820 20800
rect 25228 20748 25280 20800
rect 30656 20816 30708 20868
rect 30840 20952 30892 21004
rect 31760 20952 31812 21004
rect 31300 20927 31352 20936
rect 31300 20893 31309 20927
rect 31309 20893 31343 20927
rect 31343 20893 31352 20927
rect 31300 20884 31352 20893
rect 31576 20884 31628 20936
rect 34612 20952 34664 21004
rect 32956 20884 33008 20936
rect 36820 20884 36872 20936
rect 33140 20816 33192 20868
rect 37464 20816 37516 20868
rect 27068 20791 27120 20800
rect 27068 20757 27077 20791
rect 27077 20757 27111 20791
rect 27111 20757 27120 20791
rect 27068 20748 27120 20757
rect 29828 20791 29880 20800
rect 29828 20757 29837 20791
rect 29837 20757 29871 20791
rect 29871 20757 29880 20791
rect 29828 20748 29880 20757
rect 32772 20791 32824 20800
rect 32772 20757 32781 20791
rect 32781 20757 32815 20791
rect 32815 20757 32824 20791
rect 32772 20748 32824 20757
rect 35900 20748 35952 20800
rect 37648 20748 37700 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 4988 20544 5040 20596
rect 9956 20587 10008 20596
rect 9956 20553 9965 20587
rect 9965 20553 9999 20587
rect 9999 20553 10008 20587
rect 9956 20544 10008 20553
rect 13912 20544 13964 20596
rect 14740 20544 14792 20596
rect 9220 20476 9272 20528
rect 10968 20476 11020 20528
rect 14280 20476 14332 20528
rect 5356 20408 5408 20460
rect 7104 20408 7156 20460
rect 9404 20451 9456 20460
rect 9404 20417 9413 20451
rect 9413 20417 9447 20451
rect 9447 20417 9456 20451
rect 9404 20408 9456 20417
rect 9772 20451 9824 20460
rect 9772 20417 9781 20451
rect 9781 20417 9815 20451
rect 9815 20417 9824 20451
rect 9772 20408 9824 20417
rect 14464 20451 14516 20460
rect 14464 20417 14473 20451
rect 14473 20417 14507 20451
rect 14507 20417 14516 20451
rect 14464 20408 14516 20417
rect 4620 20340 4672 20392
rect 3976 20272 4028 20324
rect 11704 20340 11756 20392
rect 12164 20383 12216 20392
rect 12164 20349 12173 20383
rect 12173 20349 12207 20383
rect 12207 20349 12216 20383
rect 12164 20340 12216 20349
rect 14556 20383 14608 20392
rect 14556 20349 14565 20383
rect 14565 20349 14599 20383
rect 14599 20349 14608 20383
rect 14556 20340 14608 20349
rect 14740 20383 14792 20392
rect 14740 20349 14749 20383
rect 14749 20349 14783 20383
rect 14783 20349 14792 20383
rect 15292 20519 15344 20528
rect 15292 20485 15301 20519
rect 15301 20485 15335 20519
rect 15335 20485 15344 20519
rect 15292 20476 15344 20485
rect 15384 20476 15436 20528
rect 15752 20476 15804 20528
rect 17592 20476 17644 20528
rect 22652 20544 22704 20596
rect 22928 20544 22980 20596
rect 23388 20587 23440 20596
rect 23388 20553 23397 20587
rect 23397 20553 23431 20587
rect 23431 20553 23440 20587
rect 23388 20544 23440 20553
rect 25412 20544 25464 20596
rect 25872 20544 25924 20596
rect 27620 20544 27672 20596
rect 28080 20544 28132 20596
rect 32772 20544 32824 20596
rect 33140 20587 33192 20596
rect 33140 20553 33149 20587
rect 33149 20553 33183 20587
rect 33183 20553 33192 20587
rect 33140 20544 33192 20553
rect 33968 20587 34020 20596
rect 33968 20553 33977 20587
rect 33977 20553 34011 20587
rect 34011 20553 34020 20587
rect 33968 20544 34020 20553
rect 37464 20587 37516 20596
rect 37464 20553 37473 20587
rect 37473 20553 37507 20587
rect 37507 20553 37516 20587
rect 37464 20544 37516 20553
rect 14740 20340 14792 20349
rect 15384 20340 15436 20392
rect 16580 20408 16632 20460
rect 20444 20476 20496 20528
rect 18236 20408 18288 20460
rect 26700 20476 26752 20528
rect 27344 20476 27396 20528
rect 27528 20476 27580 20528
rect 29276 20519 29328 20528
rect 29276 20485 29285 20519
rect 29285 20485 29319 20519
rect 29319 20485 29328 20519
rect 29276 20476 29328 20485
rect 15660 20340 15712 20392
rect 11888 20272 11940 20324
rect 3884 20247 3936 20256
rect 3884 20213 3893 20247
rect 3893 20213 3927 20247
rect 3927 20213 3936 20247
rect 3884 20204 3936 20213
rect 6828 20204 6880 20256
rect 16488 20272 16540 20324
rect 18052 20272 18104 20324
rect 18512 20383 18564 20392
rect 18512 20349 18521 20383
rect 18521 20349 18555 20383
rect 18555 20349 18564 20383
rect 18512 20340 18564 20349
rect 19340 20340 19392 20392
rect 22100 20408 22152 20460
rect 24032 20451 24084 20460
rect 24032 20417 24041 20451
rect 24041 20417 24075 20451
rect 24075 20417 24084 20451
rect 24032 20408 24084 20417
rect 25044 20451 25096 20460
rect 25044 20417 25053 20451
rect 25053 20417 25087 20451
rect 25087 20417 25096 20451
rect 25044 20408 25096 20417
rect 25136 20408 25188 20460
rect 20904 20340 20956 20392
rect 23848 20340 23900 20392
rect 20996 20272 21048 20324
rect 24768 20272 24820 20324
rect 25780 20408 25832 20460
rect 26608 20408 26660 20460
rect 28816 20408 28868 20460
rect 29368 20408 29420 20460
rect 32220 20476 32272 20528
rect 33232 20476 33284 20528
rect 33600 20519 33652 20528
rect 33600 20485 33609 20519
rect 33609 20485 33643 20519
rect 33643 20485 33652 20519
rect 33600 20476 33652 20485
rect 29644 20451 29696 20460
rect 29644 20417 29653 20451
rect 29653 20417 29687 20451
rect 29687 20417 29696 20451
rect 29644 20408 29696 20417
rect 30104 20408 30156 20460
rect 26424 20340 26476 20392
rect 27804 20340 27856 20392
rect 27988 20383 28040 20392
rect 27988 20349 27997 20383
rect 27997 20349 28031 20383
rect 28031 20349 28040 20383
rect 27988 20340 28040 20349
rect 28264 20340 28316 20392
rect 28448 20340 28500 20392
rect 29184 20340 29236 20392
rect 29920 20340 29972 20392
rect 25412 20272 25464 20324
rect 32496 20451 32548 20460
rect 32496 20417 32505 20451
rect 32505 20417 32539 20451
rect 32539 20417 32548 20451
rect 32496 20408 32548 20417
rect 32680 20451 32732 20460
rect 32680 20417 32687 20451
rect 32687 20417 32732 20451
rect 32680 20408 32732 20417
rect 32772 20451 32824 20460
rect 32772 20417 32781 20451
rect 32781 20417 32815 20451
rect 32815 20417 32824 20451
rect 32772 20408 32824 20417
rect 33048 20408 33100 20460
rect 33140 20408 33192 20460
rect 30656 20340 30708 20392
rect 14004 20204 14056 20256
rect 14464 20204 14516 20256
rect 20536 20204 20588 20256
rect 22284 20204 22336 20256
rect 25228 20204 25280 20256
rect 26332 20204 26384 20256
rect 26884 20204 26936 20256
rect 28264 20204 28316 20256
rect 29460 20204 29512 20256
rect 30656 20247 30708 20256
rect 30656 20213 30665 20247
rect 30665 20213 30699 20247
rect 30699 20213 30708 20247
rect 30656 20204 30708 20213
rect 31484 20340 31536 20392
rect 31300 20272 31352 20324
rect 31944 20272 31996 20324
rect 32772 20272 32824 20324
rect 35532 20451 35584 20460
rect 35532 20417 35541 20451
rect 35541 20417 35575 20451
rect 35575 20417 35584 20451
rect 35532 20408 35584 20417
rect 35900 20451 35952 20460
rect 35900 20417 35909 20451
rect 35909 20417 35943 20451
rect 35943 20417 35952 20451
rect 35900 20408 35952 20417
rect 37648 20408 37700 20460
rect 38016 20383 38068 20392
rect 38016 20349 38025 20383
rect 38025 20349 38059 20383
rect 38059 20349 38068 20383
rect 38016 20340 38068 20349
rect 35992 20272 36044 20324
rect 36544 20272 36596 20324
rect 37832 20272 37884 20324
rect 34520 20204 34572 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 7104 20043 7156 20052
rect 7104 20009 7113 20043
rect 7113 20009 7147 20043
rect 7147 20009 7156 20043
rect 7104 20000 7156 20009
rect 5356 19975 5408 19984
rect 5356 19941 5365 19975
rect 5365 19941 5399 19975
rect 5399 19941 5408 19975
rect 5356 19932 5408 19941
rect 10416 19932 10468 19984
rect 3976 19907 4028 19916
rect 3976 19873 3985 19907
rect 3985 19873 4019 19907
rect 4019 19873 4028 19907
rect 3976 19864 4028 19873
rect 3884 19796 3936 19848
rect 6552 19839 6604 19848
rect 6552 19805 6561 19839
rect 6561 19805 6595 19839
rect 6595 19805 6604 19839
rect 6552 19796 6604 19805
rect 6828 19839 6880 19848
rect 6828 19805 6837 19839
rect 6837 19805 6871 19839
rect 6871 19805 6880 19839
rect 6828 19796 6880 19805
rect 6920 19839 6972 19848
rect 6920 19805 6929 19839
rect 6929 19805 6963 19839
rect 6963 19805 6972 19839
rect 6920 19796 6972 19805
rect 8208 19796 8260 19848
rect 9680 19864 9732 19916
rect 10232 19839 10284 19848
rect 6736 19771 6788 19780
rect 6736 19737 6745 19771
rect 6745 19737 6779 19771
rect 6779 19737 6788 19771
rect 6736 19728 6788 19737
rect 10232 19805 10241 19839
rect 10241 19805 10275 19839
rect 10275 19805 10284 19839
rect 10232 19796 10284 19805
rect 13820 20000 13872 20052
rect 14556 20000 14608 20052
rect 16488 20000 16540 20052
rect 19892 20000 19944 20052
rect 20260 20000 20312 20052
rect 18512 19932 18564 19984
rect 20536 19975 20588 19984
rect 16580 19864 16632 19916
rect 16672 19907 16724 19916
rect 16672 19873 16681 19907
rect 16681 19873 16715 19907
rect 16715 19873 16724 19907
rect 19432 19907 19484 19916
rect 16672 19864 16724 19873
rect 10600 19839 10652 19848
rect 10600 19805 10609 19839
rect 10609 19805 10643 19839
rect 10643 19805 10652 19839
rect 10600 19796 10652 19805
rect 15936 19796 15988 19848
rect 19432 19873 19441 19907
rect 19441 19873 19475 19907
rect 19475 19873 19484 19907
rect 19432 19864 19484 19873
rect 17408 19796 17460 19848
rect 18144 19796 18196 19848
rect 18420 19796 18472 19848
rect 20260 19864 20312 19916
rect 19892 19839 19944 19848
rect 19892 19805 19901 19839
rect 19901 19805 19935 19839
rect 19935 19805 19944 19839
rect 19892 19796 19944 19805
rect 20536 19941 20545 19975
rect 20545 19941 20579 19975
rect 20579 19941 20588 19975
rect 20536 19932 20588 19941
rect 20812 19864 20864 19916
rect 20904 19839 20956 19848
rect 20904 19805 20913 19839
rect 20913 19805 20947 19839
rect 20947 19805 20956 19839
rect 20904 19796 20956 19805
rect 21364 19796 21416 19848
rect 22284 20000 22336 20052
rect 22376 20000 22428 20052
rect 22100 19932 22152 19984
rect 22744 19932 22796 19984
rect 22376 19839 22428 19848
rect 22376 19805 22390 19839
rect 22390 19805 22424 19839
rect 22424 19805 22428 19839
rect 22376 19796 22428 19805
rect 23204 19796 23256 19848
rect 25320 20000 25372 20052
rect 29276 20000 29328 20052
rect 35900 20000 35952 20052
rect 23940 19932 23992 19984
rect 25964 19932 26016 19984
rect 26332 19932 26384 19984
rect 30748 19932 30800 19984
rect 32036 19932 32088 19984
rect 9772 19728 9824 19780
rect 10324 19728 10376 19780
rect 8392 19703 8444 19712
rect 8392 19669 8401 19703
rect 8401 19669 8435 19703
rect 8435 19669 8444 19703
rect 11704 19728 11756 19780
rect 15200 19728 15252 19780
rect 16304 19728 16356 19780
rect 16580 19771 16632 19780
rect 16580 19737 16589 19771
rect 16589 19737 16623 19771
rect 16623 19737 16632 19771
rect 16580 19728 16632 19737
rect 17776 19728 17828 19780
rect 21916 19728 21968 19780
rect 22192 19771 22244 19780
rect 22192 19737 22201 19771
rect 22201 19737 22235 19771
rect 22235 19737 22244 19771
rect 22192 19728 22244 19737
rect 8392 19660 8444 19669
rect 15292 19703 15344 19712
rect 15292 19669 15301 19703
rect 15301 19669 15335 19703
rect 15335 19669 15344 19703
rect 15292 19660 15344 19669
rect 18512 19660 18564 19712
rect 18788 19660 18840 19712
rect 28080 19864 28132 19916
rect 29828 19907 29880 19916
rect 29828 19873 29837 19907
rect 29837 19873 29871 19907
rect 29871 19873 29880 19907
rect 29828 19864 29880 19873
rect 30380 19864 30432 19916
rect 33600 19932 33652 19984
rect 24768 19839 24820 19848
rect 24768 19805 24777 19839
rect 24777 19805 24811 19839
rect 24811 19805 24820 19839
rect 24768 19796 24820 19805
rect 25136 19796 25188 19848
rect 26884 19796 26936 19848
rect 27988 19796 28040 19848
rect 29184 19796 29236 19848
rect 29460 19796 29512 19848
rect 29736 19839 29788 19848
rect 29736 19805 29745 19839
rect 29745 19805 29779 19839
rect 29779 19805 29788 19839
rect 29736 19796 29788 19805
rect 31116 19796 31168 19848
rect 31484 19839 31536 19848
rect 31484 19805 31493 19839
rect 31493 19805 31527 19839
rect 31527 19805 31536 19839
rect 31484 19796 31536 19805
rect 27068 19771 27120 19780
rect 27068 19737 27077 19771
rect 27077 19737 27111 19771
rect 27111 19737 27120 19771
rect 27068 19728 27120 19737
rect 24584 19660 24636 19712
rect 28632 19660 28684 19712
rect 29276 19728 29328 19780
rect 30288 19728 30340 19780
rect 38108 19907 38160 19916
rect 33140 19839 33192 19848
rect 33140 19805 33149 19839
rect 33149 19805 33183 19839
rect 33183 19805 33192 19839
rect 33140 19796 33192 19805
rect 33232 19728 33284 19780
rect 38108 19873 38117 19907
rect 38117 19873 38151 19907
rect 38151 19873 38160 19907
rect 38108 19864 38160 19873
rect 36820 19796 36872 19848
rect 37832 19839 37884 19848
rect 37832 19805 37841 19839
rect 37841 19805 37875 19839
rect 37875 19805 37884 19839
rect 37832 19796 37884 19805
rect 29552 19660 29604 19712
rect 31024 19660 31076 19712
rect 34980 19660 35032 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 5632 19388 5684 19440
rect 4620 19320 4672 19372
rect 6736 19320 6788 19372
rect 9496 19456 9548 19508
rect 15292 19499 15344 19508
rect 15292 19465 15301 19499
rect 15301 19465 15335 19499
rect 15335 19465 15344 19499
rect 15292 19456 15344 19465
rect 16580 19456 16632 19508
rect 19340 19499 19392 19508
rect 19340 19465 19349 19499
rect 19349 19465 19383 19499
rect 19383 19465 19392 19499
rect 19340 19456 19392 19465
rect 20536 19456 20588 19508
rect 7104 19252 7156 19304
rect 9312 19388 9364 19440
rect 7380 19184 7432 19236
rect 5080 19159 5132 19168
rect 5080 19125 5089 19159
rect 5089 19125 5123 19159
rect 5123 19125 5132 19159
rect 5080 19116 5132 19125
rect 8208 19184 8260 19236
rect 9128 19320 9180 19372
rect 9956 19320 10008 19372
rect 10600 19320 10652 19372
rect 12348 19388 12400 19440
rect 16672 19388 16724 19440
rect 20076 19388 20128 19440
rect 15660 19363 15712 19372
rect 15660 19329 15669 19363
rect 15669 19329 15703 19363
rect 15703 19329 15712 19363
rect 15660 19320 15712 19329
rect 15752 19363 15804 19372
rect 15752 19329 15761 19363
rect 15761 19329 15795 19363
rect 15795 19329 15804 19363
rect 17592 19363 17644 19372
rect 15752 19320 15804 19329
rect 17592 19329 17601 19363
rect 17601 19329 17635 19363
rect 17635 19329 17644 19363
rect 17592 19320 17644 19329
rect 17776 19363 17828 19372
rect 17776 19329 17785 19363
rect 17785 19329 17819 19363
rect 17819 19329 17828 19363
rect 17776 19320 17828 19329
rect 18512 19363 18564 19372
rect 18512 19329 18521 19363
rect 18521 19329 18555 19363
rect 18555 19329 18564 19363
rect 18512 19320 18564 19329
rect 18604 19363 18656 19372
rect 18604 19329 18613 19363
rect 18613 19329 18647 19363
rect 18647 19329 18656 19363
rect 18604 19320 18656 19329
rect 19984 19320 20036 19372
rect 20536 19363 20588 19372
rect 20536 19329 20545 19363
rect 20545 19329 20579 19363
rect 20579 19329 20588 19363
rect 20536 19320 20588 19329
rect 15936 19295 15988 19304
rect 15936 19261 15945 19295
rect 15945 19261 15979 19295
rect 15979 19261 15988 19295
rect 15936 19252 15988 19261
rect 10784 19227 10836 19236
rect 8576 19159 8628 19168
rect 8576 19125 8585 19159
rect 8585 19125 8619 19159
rect 8619 19125 8628 19159
rect 8576 19116 8628 19125
rect 10784 19193 10793 19227
rect 10793 19193 10827 19227
rect 10827 19193 10836 19227
rect 10784 19184 10836 19193
rect 14924 19184 14976 19236
rect 16764 19184 16816 19236
rect 17316 19184 17368 19236
rect 17960 19252 18012 19304
rect 20260 19252 20312 19304
rect 20812 19388 20864 19440
rect 22376 19320 22428 19372
rect 22560 19363 22612 19372
rect 22560 19329 22569 19363
rect 22569 19329 22603 19363
rect 22603 19329 22612 19363
rect 22560 19320 22612 19329
rect 22652 19363 22704 19372
rect 22652 19329 22661 19363
rect 22661 19329 22695 19363
rect 22695 19329 22704 19363
rect 22652 19320 22704 19329
rect 26884 19456 26936 19508
rect 27528 19456 27580 19508
rect 23480 19388 23532 19440
rect 25780 19388 25832 19440
rect 30012 19456 30064 19508
rect 32680 19456 32732 19508
rect 35532 19499 35584 19508
rect 23388 19363 23440 19372
rect 23388 19329 23397 19363
rect 23397 19329 23431 19363
rect 23431 19329 23440 19363
rect 23388 19320 23440 19329
rect 24308 19320 24360 19372
rect 24952 19320 25004 19372
rect 25044 19252 25096 19304
rect 22284 19184 22336 19236
rect 22836 19184 22888 19236
rect 23388 19184 23440 19236
rect 25412 19320 25464 19372
rect 26056 19363 26108 19372
rect 26056 19329 26065 19363
rect 26065 19329 26099 19363
rect 26099 19329 26108 19363
rect 26056 19320 26108 19329
rect 26332 19363 26384 19372
rect 26332 19329 26341 19363
rect 26341 19329 26375 19363
rect 26375 19329 26384 19363
rect 26332 19320 26384 19329
rect 26424 19363 26476 19372
rect 26424 19329 26433 19363
rect 26433 19329 26467 19363
rect 26467 19329 26476 19363
rect 26424 19320 26476 19329
rect 26884 19320 26936 19372
rect 27068 19252 27120 19304
rect 28816 19363 28868 19372
rect 28816 19329 28826 19363
rect 28826 19329 28860 19363
rect 28860 19329 28868 19363
rect 28816 19320 28868 19329
rect 28908 19252 28960 19304
rect 32312 19388 32364 19440
rect 33508 19388 33560 19440
rect 34428 19388 34480 19440
rect 35164 19431 35216 19440
rect 35164 19397 35173 19431
rect 35173 19397 35207 19431
rect 35207 19397 35216 19431
rect 35164 19388 35216 19397
rect 35532 19465 35541 19499
rect 35541 19465 35575 19499
rect 35575 19465 35584 19499
rect 35532 19456 35584 19465
rect 37648 19388 37700 19440
rect 29276 19320 29328 19372
rect 29828 19363 29880 19372
rect 29828 19329 29844 19363
rect 29844 19329 29878 19363
rect 29878 19329 29880 19363
rect 29828 19320 29880 19329
rect 30012 19320 30064 19372
rect 30288 19363 30340 19372
rect 30288 19329 30302 19363
rect 30302 19329 30336 19363
rect 30336 19329 30340 19363
rect 30288 19320 30340 19329
rect 30748 19320 30800 19372
rect 32680 19320 32732 19372
rect 33324 19320 33376 19372
rect 32956 19252 33008 19304
rect 34888 19363 34940 19372
rect 34888 19329 34897 19363
rect 34897 19329 34931 19363
rect 34931 19329 34940 19363
rect 35072 19363 35124 19372
rect 34888 19320 34940 19329
rect 35072 19329 35079 19363
rect 35079 19329 35124 19363
rect 35072 19320 35124 19329
rect 35532 19320 35584 19372
rect 37740 19320 37792 19372
rect 38108 19363 38160 19372
rect 38108 19329 38117 19363
rect 38117 19329 38151 19363
rect 38151 19329 38160 19363
rect 38108 19320 38160 19329
rect 31760 19184 31812 19236
rect 34980 19184 35032 19236
rect 35164 19252 35216 19304
rect 36360 19184 36412 19236
rect 9680 19116 9732 19168
rect 12256 19116 12308 19168
rect 18144 19116 18196 19168
rect 18696 19116 18748 19168
rect 20812 19116 20864 19168
rect 24492 19159 24544 19168
rect 24492 19125 24501 19159
rect 24501 19125 24535 19159
rect 24535 19125 24544 19159
rect 24492 19116 24544 19125
rect 26608 19159 26660 19168
rect 26608 19125 26617 19159
rect 26617 19125 26651 19159
rect 26651 19125 26660 19159
rect 26608 19116 26660 19125
rect 28540 19116 28592 19168
rect 29184 19116 29236 19168
rect 29736 19116 29788 19168
rect 30288 19116 30340 19168
rect 33324 19116 33376 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 9956 18955 10008 18964
rect 9956 18921 9965 18955
rect 9965 18921 9999 18955
rect 9999 18921 10008 18955
rect 9956 18912 10008 18921
rect 5632 18887 5684 18896
rect 5632 18853 5641 18887
rect 5641 18853 5675 18887
rect 5675 18853 5684 18887
rect 5632 18844 5684 18853
rect 3976 18776 4028 18828
rect 9128 18776 9180 18828
rect 9312 18844 9364 18896
rect 11428 18776 11480 18828
rect 5816 18708 5868 18760
rect 6460 18751 6512 18760
rect 6460 18717 6469 18751
rect 6469 18717 6503 18751
rect 6503 18717 6512 18751
rect 6460 18708 6512 18717
rect 7564 18708 7616 18760
rect 9496 18708 9548 18760
rect 9772 18751 9824 18760
rect 9772 18717 9781 18751
rect 9781 18717 9815 18751
rect 9815 18717 9824 18751
rect 9772 18708 9824 18717
rect 10416 18708 10468 18760
rect 13360 18708 13412 18760
rect 5080 18640 5132 18692
rect 6828 18683 6880 18692
rect 6828 18649 6837 18683
rect 6837 18649 6871 18683
rect 6871 18649 6880 18683
rect 6828 18640 6880 18649
rect 7196 18640 7248 18692
rect 7380 18683 7432 18692
rect 7380 18649 7389 18683
rect 7389 18649 7423 18683
rect 7423 18649 7432 18683
rect 7380 18640 7432 18649
rect 8392 18640 8444 18692
rect 10784 18640 10836 18692
rect 12440 18640 12492 18692
rect 13084 18640 13136 18692
rect 15660 18912 15712 18964
rect 17960 18955 18012 18964
rect 15476 18844 15528 18896
rect 15844 18844 15896 18896
rect 17960 18921 17969 18955
rect 17969 18921 18003 18955
rect 18003 18921 18012 18955
rect 17960 18912 18012 18921
rect 18144 18912 18196 18964
rect 19156 18912 19208 18964
rect 20628 18912 20680 18964
rect 24032 18912 24084 18964
rect 24492 18912 24544 18964
rect 24952 18955 25004 18964
rect 17040 18776 17092 18828
rect 14924 18708 14976 18760
rect 17132 18751 17184 18760
rect 17132 18717 17141 18751
rect 17141 18717 17175 18751
rect 17175 18717 17184 18751
rect 17132 18708 17184 18717
rect 18420 18819 18472 18828
rect 18420 18785 18429 18819
rect 18429 18785 18463 18819
rect 18463 18785 18472 18819
rect 18420 18776 18472 18785
rect 19984 18776 20036 18828
rect 21548 18776 21600 18828
rect 23480 18776 23532 18828
rect 21916 18708 21968 18760
rect 22468 18751 22520 18760
rect 22468 18717 22477 18751
rect 22477 18717 22511 18751
rect 22511 18717 22520 18751
rect 22468 18708 22520 18717
rect 23940 18819 23992 18828
rect 23940 18785 23949 18819
rect 23949 18785 23983 18819
rect 23983 18785 23992 18819
rect 24952 18921 24961 18955
rect 24961 18921 24995 18955
rect 24995 18921 25004 18955
rect 24952 18912 25004 18921
rect 29184 18912 29236 18964
rect 29736 18912 29788 18964
rect 33508 18912 33560 18964
rect 28908 18844 28960 18896
rect 29828 18844 29880 18896
rect 30472 18844 30524 18896
rect 31300 18844 31352 18896
rect 32312 18844 32364 18896
rect 32956 18844 33008 18896
rect 33048 18844 33100 18896
rect 33232 18844 33284 18896
rect 34888 18844 34940 18896
rect 36084 18844 36136 18896
rect 25872 18819 25924 18828
rect 23940 18776 23992 18785
rect 25872 18785 25881 18819
rect 25881 18785 25915 18819
rect 25915 18785 25924 18819
rect 25872 18776 25924 18785
rect 27896 18776 27948 18828
rect 30012 18776 30064 18828
rect 23848 18751 23900 18760
rect 6092 18572 6144 18624
rect 13452 18615 13504 18624
rect 13452 18581 13461 18615
rect 13461 18581 13495 18615
rect 13495 18581 13504 18615
rect 13452 18572 13504 18581
rect 14280 18572 14332 18624
rect 18512 18640 18564 18692
rect 21364 18640 21416 18692
rect 18604 18572 18656 18624
rect 19984 18572 20036 18624
rect 20168 18615 20220 18624
rect 20168 18581 20177 18615
rect 20177 18581 20211 18615
rect 20211 18581 20220 18615
rect 20168 18572 20220 18581
rect 20352 18572 20404 18624
rect 22560 18615 22612 18624
rect 22560 18581 22569 18615
rect 22569 18581 22603 18615
rect 22603 18581 22612 18615
rect 22560 18572 22612 18581
rect 23848 18717 23857 18751
rect 23857 18717 23891 18751
rect 23891 18717 23900 18751
rect 23848 18708 23900 18717
rect 29368 18708 29420 18760
rect 30840 18751 30892 18760
rect 30840 18717 30849 18751
rect 30849 18717 30883 18751
rect 30883 18717 30892 18751
rect 30840 18708 30892 18717
rect 28724 18640 28776 18692
rect 30012 18640 30064 18692
rect 31392 18708 31444 18760
rect 31576 18708 31628 18760
rect 31944 18708 31996 18760
rect 32496 18708 32548 18760
rect 33232 18751 33284 18760
rect 33232 18717 33246 18751
rect 33246 18717 33280 18751
rect 33280 18717 33284 18751
rect 33232 18708 33284 18717
rect 34796 18708 34848 18760
rect 35164 18751 35216 18760
rect 35164 18717 35174 18751
rect 35174 18717 35208 18751
rect 35208 18717 35216 18751
rect 35348 18751 35400 18760
rect 35164 18708 35216 18717
rect 35348 18717 35357 18751
rect 35357 18717 35391 18751
rect 35391 18717 35400 18751
rect 35348 18708 35400 18717
rect 33324 18640 33376 18692
rect 33600 18640 33652 18692
rect 33784 18640 33836 18692
rect 35532 18751 35584 18760
rect 35532 18717 35546 18751
rect 35546 18717 35580 18751
rect 35580 18717 35584 18751
rect 35532 18708 35584 18717
rect 36820 18708 36872 18760
rect 26792 18572 26844 18624
rect 30748 18572 30800 18624
rect 32864 18572 32916 18624
rect 32956 18572 33008 18624
rect 34888 18572 34940 18624
rect 35716 18615 35768 18624
rect 35716 18581 35725 18615
rect 35725 18581 35759 18615
rect 35759 18581 35768 18615
rect 35716 18572 35768 18581
rect 37464 18640 37516 18692
rect 37832 18572 37884 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 6460 18368 6512 18420
rect 8760 18368 8812 18420
rect 9312 18411 9364 18420
rect 9312 18377 9321 18411
rect 9321 18377 9355 18411
rect 9355 18377 9364 18411
rect 9312 18368 9364 18377
rect 10232 18368 10284 18420
rect 12256 18368 12308 18420
rect 14280 18411 14332 18420
rect 14280 18377 14289 18411
rect 14289 18377 14323 18411
rect 14323 18377 14332 18411
rect 14280 18368 14332 18377
rect 8576 18300 8628 18352
rect 7104 18232 7156 18284
rect 11428 18300 11480 18352
rect 10416 18275 10468 18284
rect 7932 18207 7984 18216
rect 7932 18173 7941 18207
rect 7941 18173 7975 18207
rect 7975 18173 7984 18207
rect 7932 18164 7984 18173
rect 9680 18164 9732 18216
rect 10416 18241 10425 18275
rect 10425 18241 10459 18275
rect 10459 18241 10468 18275
rect 10416 18232 10468 18241
rect 14740 18300 14792 18352
rect 15936 18300 15988 18352
rect 13452 18232 13504 18284
rect 15384 18232 15436 18284
rect 15844 18232 15896 18284
rect 13360 18096 13412 18148
rect 15200 18164 15252 18216
rect 17040 18232 17092 18284
rect 17316 18232 17368 18284
rect 17500 18232 17552 18284
rect 16672 18164 16724 18216
rect 17960 18368 18012 18420
rect 19984 18368 20036 18420
rect 20076 18300 20128 18352
rect 23388 18368 23440 18420
rect 25136 18368 25188 18420
rect 19340 18232 19392 18284
rect 19524 18232 19576 18284
rect 22008 18275 22060 18284
rect 22008 18241 22017 18275
rect 22017 18241 22051 18275
rect 22051 18241 22060 18275
rect 22008 18232 22060 18241
rect 18696 18207 18748 18216
rect 15752 18096 15804 18148
rect 18420 18096 18472 18148
rect 10600 18071 10652 18080
rect 10600 18037 10609 18071
rect 10609 18037 10643 18071
rect 10643 18037 10652 18071
rect 10600 18028 10652 18037
rect 12716 18071 12768 18080
rect 12716 18037 12725 18071
rect 12725 18037 12759 18071
rect 12759 18037 12768 18071
rect 12716 18028 12768 18037
rect 14004 18028 14056 18080
rect 16856 18071 16908 18080
rect 16856 18037 16865 18071
rect 16865 18037 16899 18071
rect 16899 18037 16908 18071
rect 16856 18028 16908 18037
rect 17316 18071 17368 18080
rect 17316 18037 17325 18071
rect 17325 18037 17359 18071
rect 17359 18037 17368 18071
rect 18144 18071 18196 18080
rect 17316 18028 17368 18037
rect 18144 18037 18153 18071
rect 18153 18037 18187 18071
rect 18187 18037 18196 18071
rect 18144 18028 18196 18037
rect 18696 18173 18705 18207
rect 18705 18173 18739 18207
rect 18739 18173 18748 18207
rect 18696 18164 18748 18173
rect 19432 18164 19484 18216
rect 18604 18096 18656 18148
rect 22560 18232 22612 18284
rect 23940 18300 23992 18352
rect 24676 18300 24728 18352
rect 33140 18368 33192 18420
rect 37464 18411 37516 18420
rect 37464 18377 37473 18411
rect 37473 18377 37507 18411
rect 37507 18377 37516 18411
rect 37464 18368 37516 18377
rect 37832 18411 37884 18420
rect 37832 18377 37841 18411
rect 37841 18377 37875 18411
rect 37875 18377 37884 18411
rect 37832 18368 37884 18377
rect 23480 18232 23532 18284
rect 24032 18275 24084 18284
rect 23572 18164 23624 18216
rect 24032 18241 24041 18275
rect 24041 18241 24075 18275
rect 24075 18241 24084 18275
rect 24032 18232 24084 18241
rect 26976 18232 27028 18284
rect 27712 18232 27764 18284
rect 30656 18300 30708 18352
rect 34428 18300 34480 18352
rect 37740 18300 37792 18352
rect 24124 18207 24176 18216
rect 24124 18173 24133 18207
rect 24133 18173 24167 18207
rect 24167 18173 24176 18207
rect 24124 18164 24176 18173
rect 25780 18164 25832 18216
rect 27160 18164 27212 18216
rect 30564 18275 30616 18284
rect 30564 18241 30573 18275
rect 30573 18241 30607 18275
rect 30607 18241 30616 18275
rect 30564 18232 30616 18241
rect 33416 18232 33468 18284
rect 33692 18232 33744 18284
rect 35716 18275 35768 18284
rect 35716 18241 35725 18275
rect 35725 18241 35759 18275
rect 35759 18241 35768 18275
rect 35716 18232 35768 18241
rect 35808 18275 35860 18284
rect 35808 18241 35817 18275
rect 35817 18241 35851 18275
rect 35851 18241 35860 18275
rect 35808 18232 35860 18241
rect 36360 18232 36412 18284
rect 28724 18207 28776 18216
rect 28724 18173 28733 18207
rect 28733 18173 28767 18207
rect 28767 18173 28776 18207
rect 28724 18164 28776 18173
rect 30656 18164 30708 18216
rect 31116 18207 31168 18216
rect 31116 18173 31125 18207
rect 31125 18173 31159 18207
rect 31159 18173 31168 18207
rect 31116 18164 31168 18173
rect 33600 18164 33652 18216
rect 36176 18164 36228 18216
rect 38016 18207 38068 18216
rect 38016 18173 38025 18207
rect 38025 18173 38059 18207
rect 38059 18173 38068 18207
rect 38016 18164 38068 18173
rect 19432 18028 19484 18080
rect 20168 18028 20220 18080
rect 23756 18096 23808 18148
rect 27896 18096 27948 18148
rect 29092 18096 29144 18148
rect 35440 18096 35492 18148
rect 35992 18139 36044 18148
rect 35992 18105 36001 18139
rect 36001 18105 36035 18139
rect 36035 18105 36044 18139
rect 35992 18096 36044 18105
rect 36636 18096 36688 18148
rect 22468 18071 22520 18080
rect 22468 18037 22477 18071
rect 22477 18037 22511 18071
rect 22511 18037 22520 18071
rect 22468 18028 22520 18037
rect 23204 18028 23256 18080
rect 23664 18028 23716 18080
rect 33508 18028 33560 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 11428 17867 11480 17876
rect 11428 17833 11437 17867
rect 11437 17833 11471 17867
rect 11471 17833 11480 17867
rect 11428 17824 11480 17833
rect 15108 17824 15160 17876
rect 21548 17824 21600 17876
rect 15200 17756 15252 17808
rect 17500 17756 17552 17808
rect 5816 17731 5868 17740
rect 5816 17697 5825 17731
rect 5825 17697 5859 17731
rect 5859 17697 5868 17731
rect 5816 17688 5868 17697
rect 9128 17688 9180 17740
rect 12716 17688 12768 17740
rect 14004 17688 14056 17740
rect 6092 17663 6144 17672
rect 6092 17629 6126 17663
rect 6126 17629 6144 17663
rect 6092 17620 6144 17629
rect 10600 17620 10652 17672
rect 13084 17620 13136 17672
rect 16856 17688 16908 17740
rect 13820 17552 13872 17604
rect 15108 17663 15160 17672
rect 15108 17629 15122 17663
rect 15122 17629 15156 17663
rect 15156 17629 15160 17663
rect 19524 17663 19576 17672
rect 15108 17620 15160 17629
rect 14924 17595 14976 17604
rect 14924 17561 14933 17595
rect 14933 17561 14967 17595
rect 14967 17561 14976 17595
rect 14924 17552 14976 17561
rect 19524 17629 19533 17663
rect 19533 17629 19567 17663
rect 19567 17629 19576 17663
rect 19524 17620 19576 17629
rect 20168 17756 20220 17808
rect 21272 17663 21324 17672
rect 21272 17629 21281 17663
rect 21281 17629 21315 17663
rect 21315 17629 21324 17663
rect 21272 17620 21324 17629
rect 22652 17688 22704 17740
rect 22100 17620 22152 17672
rect 24032 17824 24084 17876
rect 23112 17688 23164 17740
rect 24124 17688 24176 17740
rect 23204 17663 23256 17672
rect 23204 17629 23213 17663
rect 23213 17629 23247 17663
rect 23247 17629 23256 17663
rect 23204 17620 23256 17629
rect 23572 17620 23624 17672
rect 23940 17620 23992 17672
rect 7196 17527 7248 17536
rect 7196 17493 7205 17527
rect 7205 17493 7239 17527
rect 7239 17493 7248 17527
rect 7196 17484 7248 17493
rect 12348 17527 12400 17536
rect 12348 17493 12357 17527
rect 12357 17493 12391 17527
rect 12391 17493 12400 17527
rect 12348 17484 12400 17493
rect 13084 17484 13136 17536
rect 15476 17552 15528 17604
rect 18052 17552 18104 17604
rect 21456 17595 21508 17604
rect 21456 17561 21465 17595
rect 21465 17561 21499 17595
rect 21499 17561 21508 17595
rect 21456 17552 21508 17561
rect 22192 17552 22244 17604
rect 23756 17552 23808 17604
rect 25596 17824 25648 17876
rect 24676 17731 24728 17740
rect 24676 17697 24685 17731
rect 24685 17697 24719 17731
rect 24719 17697 24728 17731
rect 24676 17688 24728 17697
rect 24768 17663 24820 17672
rect 24768 17629 24777 17663
rect 24777 17629 24811 17663
rect 24811 17629 24820 17663
rect 24768 17620 24820 17629
rect 25320 17663 25372 17672
rect 25320 17629 25329 17663
rect 25329 17629 25363 17663
rect 25363 17629 25372 17663
rect 25320 17620 25372 17629
rect 26332 17620 26384 17672
rect 29092 17824 29144 17876
rect 30288 17867 30340 17876
rect 30288 17833 30297 17867
rect 30297 17833 30331 17867
rect 30331 17833 30340 17867
rect 30288 17824 30340 17833
rect 31116 17824 31168 17876
rect 33508 17867 33560 17876
rect 33508 17833 33517 17867
rect 33517 17833 33551 17867
rect 33551 17833 33560 17867
rect 33508 17824 33560 17833
rect 28724 17756 28776 17808
rect 27344 17688 27396 17740
rect 30564 17688 30616 17740
rect 26608 17620 26660 17672
rect 27160 17663 27212 17672
rect 27160 17629 27170 17663
rect 27170 17629 27204 17663
rect 27204 17629 27212 17663
rect 27160 17620 27212 17629
rect 28080 17620 28132 17672
rect 29828 17663 29880 17672
rect 29828 17629 29870 17663
rect 29870 17629 29880 17663
rect 30380 17663 30432 17672
rect 29828 17620 29880 17629
rect 30380 17629 30389 17663
rect 30389 17629 30423 17663
rect 30423 17629 30432 17663
rect 30380 17620 30432 17629
rect 30932 17620 30984 17672
rect 26700 17552 26752 17604
rect 27436 17595 27488 17604
rect 27436 17561 27445 17595
rect 27445 17561 27479 17595
rect 27479 17561 27488 17595
rect 31024 17595 31076 17604
rect 27436 17552 27488 17561
rect 31024 17561 31033 17595
rect 31033 17561 31067 17595
rect 31067 17561 31076 17595
rect 31024 17552 31076 17561
rect 31300 17552 31352 17604
rect 15660 17484 15712 17536
rect 16120 17527 16172 17536
rect 16120 17493 16129 17527
rect 16129 17493 16163 17527
rect 16163 17493 16172 17527
rect 16120 17484 16172 17493
rect 17960 17484 18012 17536
rect 20076 17484 20128 17536
rect 23112 17527 23164 17536
rect 23112 17493 23121 17527
rect 23121 17493 23155 17527
rect 23155 17493 23164 17527
rect 23112 17484 23164 17493
rect 24124 17484 24176 17536
rect 24584 17484 24636 17536
rect 25688 17484 25740 17536
rect 27988 17484 28040 17536
rect 29736 17527 29788 17536
rect 29736 17493 29745 17527
rect 29745 17493 29779 17527
rect 29779 17493 29788 17527
rect 29736 17484 29788 17493
rect 29920 17527 29972 17536
rect 29920 17493 29929 17527
rect 29929 17493 29963 17527
rect 29963 17493 29972 17527
rect 29920 17484 29972 17493
rect 36728 17756 36780 17808
rect 33048 17688 33100 17740
rect 38108 17731 38160 17740
rect 38108 17697 38117 17731
rect 38117 17697 38151 17731
rect 38151 17697 38160 17731
rect 38108 17688 38160 17697
rect 33140 17663 33192 17672
rect 31944 17552 31996 17604
rect 32128 17595 32180 17604
rect 32128 17561 32137 17595
rect 32137 17561 32171 17595
rect 32171 17561 32180 17595
rect 32128 17552 32180 17561
rect 33140 17629 33149 17663
rect 33149 17629 33183 17663
rect 33183 17629 33192 17663
rect 33140 17620 33192 17629
rect 33324 17620 33376 17672
rect 37832 17663 37884 17672
rect 37832 17629 37841 17663
rect 37841 17629 37875 17663
rect 37875 17629 37884 17663
rect 37832 17620 37884 17629
rect 33232 17484 33284 17536
rect 33692 17484 33744 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 7196 17280 7248 17332
rect 7656 17212 7708 17264
rect 10508 17212 10560 17264
rect 12348 17212 12400 17264
rect 14924 17280 14976 17332
rect 15476 17323 15528 17332
rect 15476 17289 15485 17323
rect 15485 17289 15519 17323
rect 15519 17289 15528 17323
rect 15476 17280 15528 17289
rect 19340 17280 19392 17332
rect 23112 17280 23164 17332
rect 23848 17280 23900 17332
rect 25320 17280 25372 17332
rect 30380 17280 30432 17332
rect 8024 17144 8076 17196
rect 8208 17144 8260 17196
rect 17316 17212 17368 17264
rect 18144 17212 18196 17264
rect 15200 17144 15252 17196
rect 15660 17187 15712 17196
rect 15660 17153 15669 17187
rect 15669 17153 15703 17187
rect 15703 17153 15712 17187
rect 15660 17144 15712 17153
rect 15844 17187 15896 17196
rect 15844 17153 15853 17187
rect 15853 17153 15887 17187
rect 15887 17153 15896 17187
rect 15844 17144 15896 17153
rect 18052 17144 18104 17196
rect 18236 17187 18288 17196
rect 18236 17153 18245 17187
rect 18245 17153 18279 17187
rect 18279 17153 18288 17187
rect 18236 17144 18288 17153
rect 22928 17212 22980 17264
rect 23204 17212 23256 17264
rect 23020 17144 23072 17196
rect 27344 17255 27396 17264
rect 27344 17221 27353 17255
rect 27353 17221 27387 17255
rect 27387 17221 27396 17255
rect 27344 17212 27396 17221
rect 27712 17212 27764 17264
rect 7840 17076 7892 17128
rect 11704 17119 11756 17128
rect 11704 17085 11713 17119
rect 11713 17085 11747 17119
rect 11747 17085 11756 17119
rect 11704 17076 11756 17085
rect 15568 17076 15620 17128
rect 17132 17076 17184 17128
rect 22836 17076 22888 17128
rect 24584 17187 24636 17196
rect 24584 17153 24593 17187
rect 24593 17153 24627 17187
rect 24627 17153 24636 17187
rect 26056 17187 26108 17196
rect 24584 17144 24636 17153
rect 26056 17153 26065 17187
rect 26065 17153 26099 17187
rect 26099 17153 26108 17187
rect 26056 17144 26108 17153
rect 26332 17187 26384 17196
rect 26332 17153 26341 17187
rect 26341 17153 26375 17187
rect 26375 17153 26384 17187
rect 26332 17144 26384 17153
rect 26424 17187 26476 17196
rect 26424 17153 26433 17187
rect 26433 17153 26467 17187
rect 26467 17153 26476 17187
rect 26424 17144 26476 17153
rect 27436 17187 27488 17196
rect 24032 17076 24084 17128
rect 24768 17119 24820 17128
rect 24768 17085 24777 17119
rect 24777 17085 24811 17119
rect 24811 17085 24820 17119
rect 24768 17076 24820 17085
rect 25780 17076 25832 17128
rect 13084 17051 13136 17060
rect 13084 17017 13093 17051
rect 13093 17017 13127 17051
rect 13127 17017 13136 17051
rect 13084 17008 13136 17017
rect 13544 17008 13596 17060
rect 15384 17008 15436 17060
rect 8668 16983 8720 16992
rect 8668 16949 8677 16983
rect 8677 16949 8711 16983
rect 8711 16949 8720 16983
rect 8668 16940 8720 16949
rect 14740 16940 14792 16992
rect 15108 16940 15160 16992
rect 22468 17008 22520 17060
rect 23940 17008 23992 17060
rect 27436 17153 27445 17187
rect 27445 17153 27479 17187
rect 27479 17153 27488 17187
rect 27436 17144 27488 17153
rect 28724 17212 28776 17264
rect 29184 17212 29236 17264
rect 30656 17212 30708 17264
rect 31300 17212 31352 17264
rect 32588 17212 32640 17264
rect 37740 17280 37792 17332
rect 37832 17280 37884 17332
rect 27344 17076 27396 17128
rect 28080 17076 28132 17128
rect 28724 17076 28776 17128
rect 30012 17187 30064 17196
rect 30012 17153 30021 17187
rect 30021 17153 30055 17187
rect 30055 17153 30064 17187
rect 30012 17144 30064 17153
rect 30840 17144 30892 17196
rect 33232 17144 33284 17196
rect 31944 17076 31996 17128
rect 32404 17076 32456 17128
rect 32864 17119 32916 17128
rect 32864 17085 32873 17119
rect 32873 17085 32907 17119
rect 32907 17085 32916 17119
rect 32864 17076 32916 17085
rect 34244 17144 34296 17196
rect 34796 17144 34848 17196
rect 35164 17187 35216 17196
rect 35164 17153 35174 17187
rect 35174 17153 35208 17187
rect 35208 17153 35216 17187
rect 35348 17187 35400 17196
rect 35164 17144 35216 17153
rect 35348 17153 35357 17187
rect 35357 17153 35391 17187
rect 35391 17153 35400 17187
rect 35348 17144 35400 17153
rect 35532 17187 35584 17196
rect 35532 17153 35546 17187
rect 35546 17153 35580 17187
rect 35580 17153 35584 17187
rect 35532 17144 35584 17153
rect 23112 16940 23164 16992
rect 31024 17008 31076 17060
rect 33324 17008 33376 17060
rect 36728 17187 36780 17196
rect 27712 16983 27764 16992
rect 27712 16949 27721 16983
rect 27721 16949 27755 16983
rect 27755 16949 27764 16983
rect 27712 16940 27764 16949
rect 29276 16940 29328 16992
rect 32956 16940 33008 16992
rect 35348 16940 35400 16992
rect 36728 17153 36737 17187
rect 36737 17153 36771 17187
rect 36771 17153 36780 17187
rect 36728 17144 36780 17153
rect 37740 17144 37792 17196
rect 36636 17119 36688 17128
rect 36636 17085 36645 17119
rect 36645 17085 36679 17119
rect 36679 17085 36688 17119
rect 36636 17076 36688 17085
rect 38016 17119 38068 17128
rect 38016 17085 38025 17119
rect 38025 17085 38059 17119
rect 38059 17085 38068 17119
rect 38016 17076 38068 17085
rect 37096 16940 37148 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 8024 16779 8076 16788
rect 8024 16745 8033 16779
rect 8033 16745 8067 16779
rect 8067 16745 8076 16779
rect 8024 16736 8076 16745
rect 8208 16736 8260 16788
rect 10508 16779 10560 16788
rect 7932 16668 7984 16720
rect 10508 16745 10517 16779
rect 10517 16745 10551 16779
rect 10551 16745 10560 16779
rect 10508 16736 10560 16745
rect 7840 16600 7892 16652
rect 10876 16668 10928 16720
rect 6920 16532 6972 16584
rect 8208 16575 8260 16584
rect 8208 16541 8217 16575
rect 8217 16541 8251 16575
rect 8251 16541 8260 16575
rect 8208 16532 8260 16541
rect 8668 16532 8720 16584
rect 13084 16668 13136 16720
rect 15476 16668 15528 16720
rect 11704 16600 11756 16652
rect 14188 16600 14240 16652
rect 18236 16736 18288 16788
rect 17960 16668 18012 16720
rect 22008 16736 22060 16788
rect 22836 16779 22888 16788
rect 22836 16745 22845 16779
rect 22845 16745 22879 16779
rect 22879 16745 22888 16779
rect 22836 16736 22888 16745
rect 23940 16736 23992 16788
rect 22652 16668 22704 16720
rect 26332 16668 26384 16720
rect 27712 16736 27764 16788
rect 27896 16668 27948 16720
rect 26424 16600 26476 16652
rect 11888 16575 11940 16584
rect 11888 16541 11897 16575
rect 11897 16541 11931 16575
rect 11931 16541 11940 16575
rect 11888 16532 11940 16541
rect 12440 16532 12492 16584
rect 13636 16532 13688 16584
rect 15384 16575 15436 16584
rect 15384 16541 15393 16575
rect 15393 16541 15427 16575
rect 15427 16541 15436 16575
rect 15384 16532 15436 16541
rect 15568 16532 15620 16584
rect 16120 16532 16172 16584
rect 20076 16532 20128 16584
rect 21824 16532 21876 16584
rect 22100 16532 22152 16584
rect 22468 16575 22520 16584
rect 22468 16541 22477 16575
rect 22477 16541 22511 16575
rect 22511 16541 22520 16575
rect 22468 16532 22520 16541
rect 22928 16575 22980 16584
rect 22928 16541 22937 16575
rect 22937 16541 22971 16575
rect 22971 16541 22980 16575
rect 22928 16532 22980 16541
rect 23112 16532 23164 16584
rect 26240 16532 26292 16584
rect 26516 16575 26568 16584
rect 26516 16541 26525 16575
rect 26525 16541 26559 16575
rect 26559 16541 26568 16575
rect 26516 16532 26568 16541
rect 26700 16575 26752 16584
rect 26700 16541 26709 16575
rect 26709 16541 26743 16575
rect 26743 16541 26752 16575
rect 26700 16532 26752 16541
rect 27344 16600 27396 16652
rect 28908 16736 28960 16788
rect 32220 16736 32272 16788
rect 33140 16736 33192 16788
rect 37740 16736 37792 16788
rect 29092 16643 29144 16652
rect 29092 16609 29101 16643
rect 29101 16609 29135 16643
rect 29135 16609 29144 16643
rect 29092 16600 29144 16609
rect 28908 16575 28960 16584
rect 28908 16541 28917 16575
rect 28917 16541 28951 16575
rect 28951 16541 28960 16575
rect 29184 16575 29236 16584
rect 28908 16532 28960 16541
rect 29184 16541 29193 16575
rect 29193 16541 29227 16575
rect 29227 16541 29236 16575
rect 29460 16600 29512 16652
rect 31576 16600 31628 16652
rect 33416 16600 33468 16652
rect 34704 16600 34756 16652
rect 29184 16532 29236 16541
rect 31300 16575 31352 16584
rect 6552 16464 6604 16516
rect 10692 16464 10744 16516
rect 13544 16464 13596 16516
rect 17960 16464 18012 16516
rect 26056 16464 26108 16516
rect 26792 16507 26844 16516
rect 26792 16473 26801 16507
rect 26801 16473 26835 16507
rect 26835 16473 26844 16507
rect 26792 16464 26844 16473
rect 30932 16464 30984 16516
rect 31300 16541 31309 16575
rect 31309 16541 31343 16575
rect 31343 16541 31352 16575
rect 31300 16532 31352 16541
rect 31392 16575 31444 16584
rect 31392 16541 31401 16575
rect 31401 16541 31435 16575
rect 31435 16541 31444 16575
rect 31852 16575 31904 16584
rect 31392 16532 31444 16541
rect 31852 16541 31861 16575
rect 31861 16541 31895 16575
rect 31895 16541 31904 16575
rect 31852 16532 31904 16541
rect 31668 16464 31720 16516
rect 7012 16439 7064 16448
rect 7012 16405 7021 16439
rect 7021 16405 7055 16439
rect 7055 16405 7064 16439
rect 7012 16396 7064 16405
rect 12072 16439 12124 16448
rect 12072 16405 12081 16439
rect 12081 16405 12115 16439
rect 12115 16405 12124 16439
rect 12072 16396 12124 16405
rect 22928 16396 22980 16448
rect 27620 16396 27672 16448
rect 27804 16396 27856 16448
rect 28908 16396 28960 16448
rect 30656 16396 30708 16448
rect 30840 16439 30892 16448
rect 30840 16405 30849 16439
rect 30849 16405 30883 16439
rect 30883 16405 30892 16439
rect 30840 16396 30892 16405
rect 32220 16575 32272 16584
rect 32220 16541 32229 16575
rect 32229 16541 32263 16575
rect 32263 16541 32272 16575
rect 32220 16532 32272 16541
rect 32404 16532 32456 16584
rect 33692 16575 33744 16584
rect 33692 16541 33701 16575
rect 33701 16541 33735 16575
rect 33735 16541 33744 16575
rect 33692 16532 33744 16541
rect 34796 16532 34848 16584
rect 35072 16575 35124 16584
rect 35072 16541 35081 16575
rect 35081 16541 35115 16575
rect 35115 16541 35124 16575
rect 35072 16532 35124 16541
rect 35164 16575 35216 16584
rect 35164 16541 35174 16575
rect 35174 16541 35208 16575
rect 35208 16541 35216 16575
rect 35440 16600 35492 16652
rect 36820 16643 36872 16652
rect 36820 16609 36829 16643
rect 36829 16609 36863 16643
rect 36863 16609 36872 16643
rect 36820 16600 36872 16609
rect 35164 16532 35216 16541
rect 35532 16575 35584 16584
rect 35532 16541 35546 16575
rect 35546 16541 35580 16575
rect 35580 16541 35584 16575
rect 37096 16575 37148 16584
rect 35532 16532 35584 16541
rect 37096 16541 37130 16575
rect 37130 16541 37148 16575
rect 37096 16532 37148 16541
rect 32864 16464 32916 16516
rect 37832 16464 37884 16516
rect 35716 16439 35768 16448
rect 35716 16405 35725 16439
rect 35725 16405 35759 16439
rect 35759 16405 35768 16439
rect 35716 16396 35768 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 6552 16235 6604 16244
rect 6552 16201 6561 16235
rect 6561 16201 6595 16235
rect 6595 16201 6604 16235
rect 6552 16192 6604 16201
rect 8392 16192 8444 16244
rect 13544 16235 13596 16244
rect 7012 16124 7064 16176
rect 12072 16124 12124 16176
rect 13544 16201 13553 16235
rect 13553 16201 13587 16235
rect 13587 16201 13596 16235
rect 13544 16192 13596 16201
rect 17224 16192 17276 16244
rect 25320 16235 25372 16244
rect 15752 16124 15804 16176
rect 25320 16201 25329 16235
rect 25329 16201 25363 16235
rect 25363 16201 25372 16235
rect 25320 16192 25372 16201
rect 8116 16056 8168 16108
rect 14188 16099 14240 16108
rect 14188 16065 14197 16099
rect 14197 16065 14231 16099
rect 14231 16065 14240 16099
rect 14188 16056 14240 16065
rect 17592 16099 17644 16108
rect 17592 16065 17601 16099
rect 17601 16065 17635 16099
rect 17635 16065 17644 16099
rect 17592 16056 17644 16065
rect 17776 16099 17828 16108
rect 17776 16065 17785 16099
rect 17785 16065 17819 16099
rect 17819 16065 17828 16099
rect 17776 16056 17828 16065
rect 17868 16099 17920 16108
rect 17868 16065 17877 16099
rect 17877 16065 17911 16099
rect 17911 16065 17920 16099
rect 21640 16124 21692 16176
rect 22468 16124 22520 16176
rect 23020 16124 23072 16176
rect 17868 16056 17920 16065
rect 7104 15988 7156 16040
rect 8392 16031 8444 16040
rect 8392 15997 8401 16031
rect 8401 15997 8435 16031
rect 8435 15997 8444 16031
rect 8392 15988 8444 15997
rect 12164 16031 12216 16040
rect 12164 15997 12173 16031
rect 12173 15997 12207 16031
rect 12207 15997 12216 16031
rect 12164 15988 12216 15997
rect 14464 16031 14516 16040
rect 14464 15997 14473 16031
rect 14473 15997 14507 16031
rect 14507 15997 14516 16031
rect 14464 15988 14516 15997
rect 20536 16056 20588 16108
rect 22560 16056 22612 16108
rect 26516 16056 26568 16108
rect 27160 16056 27212 16108
rect 27620 16099 27672 16108
rect 27620 16065 27629 16099
rect 27629 16065 27663 16099
rect 27663 16065 27672 16099
rect 27620 16056 27672 16065
rect 27896 16056 27948 16108
rect 29828 16124 29880 16176
rect 29276 16099 29328 16108
rect 29276 16065 29285 16099
rect 29285 16065 29319 16099
rect 29319 16065 29328 16099
rect 29460 16099 29512 16108
rect 29276 16056 29328 16065
rect 29460 16065 29469 16099
rect 29469 16065 29503 16099
rect 29503 16065 29512 16099
rect 29460 16056 29512 16065
rect 25780 15988 25832 16040
rect 26056 15988 26108 16040
rect 27528 16031 27580 16040
rect 27528 15997 27541 16031
rect 27541 15997 27575 16031
rect 27575 15997 27580 16031
rect 27528 15988 27580 15997
rect 29000 15988 29052 16040
rect 31392 16192 31444 16244
rect 32220 16192 32272 16244
rect 35532 16192 35584 16244
rect 37832 16235 37884 16244
rect 30564 16124 30616 16176
rect 31484 16124 31536 16176
rect 31944 16124 31996 16176
rect 32588 16167 32640 16176
rect 30472 16056 30524 16108
rect 31208 16056 31260 16108
rect 32588 16133 32597 16167
rect 32597 16133 32631 16167
rect 32631 16133 32640 16167
rect 32588 16124 32640 16133
rect 32956 16124 33008 16176
rect 32680 16099 32732 16108
rect 32680 16065 32689 16099
rect 32689 16065 32723 16099
rect 32723 16065 32732 16099
rect 32680 16056 32732 16065
rect 35716 16099 35768 16108
rect 35716 16065 35725 16099
rect 35725 16065 35759 16099
rect 35759 16065 35768 16099
rect 35716 16056 35768 16065
rect 37832 16201 37841 16235
rect 37841 16201 37875 16235
rect 37875 16201 37884 16235
rect 37832 16192 37884 16201
rect 38016 16031 38068 16040
rect 38016 15997 38025 16031
rect 38025 15997 38059 16031
rect 38059 15997 38068 16031
rect 38016 15988 38068 15997
rect 24952 15920 25004 15972
rect 26976 15920 27028 15972
rect 30472 15920 30524 15972
rect 31300 15920 31352 15972
rect 36636 15920 36688 15972
rect 37832 15920 37884 15972
rect 7748 15895 7800 15904
rect 7748 15861 7757 15895
rect 7757 15861 7791 15895
rect 7791 15861 7800 15895
rect 7748 15852 7800 15861
rect 8300 15895 8352 15904
rect 8300 15861 8309 15895
rect 8309 15861 8343 15895
rect 8343 15861 8352 15895
rect 8300 15852 8352 15861
rect 17500 15852 17552 15904
rect 22928 15895 22980 15904
rect 22928 15861 22937 15895
rect 22937 15861 22971 15895
rect 22971 15861 22980 15895
rect 22928 15852 22980 15861
rect 25228 15852 25280 15904
rect 27344 15852 27396 15904
rect 29276 15852 29328 15904
rect 30012 15852 30064 15904
rect 32680 15852 32732 15904
rect 37188 15852 37240 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 6920 15648 6972 15700
rect 8392 15648 8444 15700
rect 17776 15648 17828 15700
rect 24952 15691 25004 15700
rect 24952 15657 24961 15691
rect 24961 15657 24995 15691
rect 24995 15657 25004 15691
rect 24952 15648 25004 15657
rect 11152 15623 11204 15632
rect 11152 15589 11161 15623
rect 11161 15589 11195 15623
rect 11195 15589 11204 15623
rect 11152 15580 11204 15589
rect 7748 15444 7800 15496
rect 12164 15444 12216 15496
rect 17868 15580 17920 15632
rect 20168 15623 20220 15632
rect 17776 15512 17828 15564
rect 20168 15589 20177 15623
rect 20177 15589 20211 15623
rect 20211 15589 20220 15623
rect 20168 15580 20220 15589
rect 26792 15648 26844 15700
rect 27896 15648 27948 15700
rect 29460 15648 29512 15700
rect 25872 15623 25924 15632
rect 16028 15487 16080 15496
rect 10048 15419 10100 15428
rect 10048 15385 10082 15419
rect 10082 15385 10100 15419
rect 16028 15453 16037 15487
rect 16037 15453 16071 15487
rect 16071 15453 16080 15487
rect 16028 15444 16080 15453
rect 17592 15487 17644 15496
rect 17592 15453 17601 15487
rect 17601 15453 17635 15487
rect 17635 15453 17644 15487
rect 17592 15444 17644 15453
rect 20260 15512 20312 15564
rect 10048 15376 10100 15385
rect 17776 15376 17828 15428
rect 21456 15444 21508 15496
rect 25872 15589 25881 15623
rect 25881 15589 25915 15623
rect 25915 15589 25924 15623
rect 25872 15580 25924 15589
rect 26056 15580 26108 15632
rect 31116 15648 31168 15700
rect 34520 15648 34572 15700
rect 36360 15691 36412 15700
rect 36360 15657 36369 15691
rect 36369 15657 36403 15691
rect 36403 15657 36412 15691
rect 36360 15648 36412 15657
rect 22836 15512 22888 15564
rect 22192 15487 22244 15496
rect 22192 15453 22201 15487
rect 22201 15453 22235 15487
rect 22235 15453 22244 15487
rect 22192 15444 22244 15453
rect 22468 15444 22520 15496
rect 23020 15444 23072 15496
rect 24216 15512 24268 15564
rect 24400 15444 24452 15496
rect 25504 15444 25556 15496
rect 25320 15376 25372 15428
rect 15936 15308 15988 15360
rect 17684 15351 17736 15360
rect 17684 15317 17693 15351
rect 17693 15317 17727 15351
rect 17727 15317 17736 15351
rect 17684 15308 17736 15317
rect 20168 15308 20220 15360
rect 25136 15351 25188 15360
rect 25136 15317 25145 15351
rect 25145 15317 25179 15351
rect 25179 15317 25188 15351
rect 25136 15308 25188 15317
rect 26516 15512 26568 15564
rect 33140 15580 33192 15632
rect 30840 15512 30892 15564
rect 31576 15555 31628 15564
rect 31576 15521 31585 15555
rect 31585 15521 31619 15555
rect 31619 15521 31628 15555
rect 31576 15512 31628 15521
rect 33508 15580 33560 15632
rect 38108 15555 38160 15564
rect 26976 15487 27028 15496
rect 26976 15453 26985 15487
rect 26985 15453 27019 15487
rect 27019 15453 27028 15487
rect 26976 15444 27028 15453
rect 27160 15487 27212 15496
rect 27160 15453 27169 15487
rect 27169 15453 27203 15487
rect 27203 15453 27212 15487
rect 27160 15444 27212 15453
rect 28080 15487 28132 15496
rect 28080 15453 28089 15487
rect 28089 15453 28123 15487
rect 28123 15453 28132 15487
rect 28080 15444 28132 15453
rect 28172 15444 28224 15496
rect 28632 15444 28684 15496
rect 29736 15487 29788 15496
rect 29736 15453 29745 15487
rect 29745 15453 29779 15487
rect 29779 15453 29788 15487
rect 29736 15444 29788 15453
rect 29828 15444 29880 15496
rect 38108 15521 38117 15555
rect 38117 15521 38151 15555
rect 38151 15521 38160 15555
rect 38108 15512 38160 15521
rect 33508 15444 33560 15496
rect 34796 15444 34848 15496
rect 37832 15487 37884 15496
rect 37832 15453 37841 15487
rect 37841 15453 37875 15487
rect 37875 15453 37884 15487
rect 37832 15444 37884 15453
rect 28724 15308 28776 15360
rect 31116 15351 31168 15360
rect 31116 15317 31125 15351
rect 31125 15317 31159 15351
rect 31159 15317 31168 15351
rect 31116 15308 31168 15317
rect 31668 15308 31720 15360
rect 33416 15351 33468 15360
rect 33416 15317 33425 15351
rect 33425 15317 33459 15351
rect 33459 15317 33468 15351
rect 33416 15308 33468 15317
rect 33508 15308 33560 15360
rect 34704 15376 34756 15428
rect 38016 15308 38068 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 8852 15147 8904 15156
rect 8852 15113 8861 15147
rect 8861 15113 8895 15147
rect 8895 15113 8904 15147
rect 8852 15104 8904 15113
rect 10048 15147 10100 15156
rect 10048 15113 10057 15147
rect 10057 15113 10091 15147
rect 10091 15113 10100 15147
rect 10048 15104 10100 15113
rect 14464 15104 14516 15156
rect 16028 15104 16080 15156
rect 16764 15104 16816 15156
rect 20352 15104 20404 15156
rect 9312 14968 9364 15020
rect 10140 14968 10192 15020
rect 11152 14968 11204 15020
rect 16580 15036 16632 15088
rect 11888 14968 11940 15020
rect 13360 15011 13412 15020
rect 13360 14977 13369 15011
rect 13369 14977 13403 15011
rect 13403 14977 13412 15011
rect 13360 14968 13412 14977
rect 15200 15011 15252 15020
rect 8300 14900 8352 14952
rect 10600 14900 10652 14952
rect 13452 14943 13504 14952
rect 13452 14909 13461 14943
rect 13461 14909 13495 14943
rect 13495 14909 13504 14943
rect 13452 14900 13504 14909
rect 15200 14977 15209 15011
rect 15209 14977 15243 15011
rect 15243 14977 15252 15011
rect 15200 14968 15252 14977
rect 15936 15011 15988 15020
rect 15936 14977 15945 15011
rect 15945 14977 15979 15011
rect 15979 14977 15988 15011
rect 15936 14968 15988 14977
rect 16856 14968 16908 15020
rect 17040 14968 17092 15020
rect 17868 15036 17920 15088
rect 18052 15036 18104 15088
rect 21088 15079 21140 15088
rect 17592 14968 17644 15020
rect 17776 14968 17828 15020
rect 18880 14968 18932 15020
rect 19340 15011 19392 15020
rect 19340 14977 19349 15011
rect 19349 14977 19383 15011
rect 19383 14977 19392 15011
rect 19340 14968 19392 14977
rect 19432 15011 19484 15020
rect 19432 14977 19441 15011
rect 19441 14977 19475 15011
rect 19475 14977 19484 15011
rect 21088 15045 21097 15079
rect 21097 15045 21131 15079
rect 21131 15045 21140 15079
rect 21088 15036 21140 15045
rect 19432 14968 19484 14977
rect 20720 14968 20772 15020
rect 12532 14832 12584 14884
rect 13544 14832 13596 14884
rect 15384 14875 15436 14884
rect 15384 14841 15393 14875
rect 15393 14841 15427 14875
rect 15427 14841 15436 14875
rect 15384 14832 15436 14841
rect 8392 14807 8444 14816
rect 8392 14773 8401 14807
rect 8401 14773 8435 14807
rect 8435 14773 8444 14807
rect 8392 14764 8444 14773
rect 11152 14764 11204 14816
rect 15292 14764 15344 14816
rect 16672 14764 16724 14816
rect 17868 14900 17920 14952
rect 17960 14943 18012 14952
rect 17960 14909 17969 14943
rect 17969 14909 18003 14943
rect 18003 14909 18012 14943
rect 17960 14900 18012 14909
rect 19708 14900 19760 14952
rect 18328 14875 18380 14884
rect 18328 14841 18337 14875
rect 18337 14841 18371 14875
rect 18371 14841 18380 14875
rect 18328 14832 18380 14841
rect 20352 14832 20404 14884
rect 21916 14968 21968 15020
rect 25136 15036 25188 15088
rect 31576 15104 31628 15156
rect 26240 15036 26292 15088
rect 31484 15079 31536 15088
rect 31484 15045 31493 15079
rect 31493 15045 31527 15079
rect 31527 15045 31536 15079
rect 31484 15036 31536 15045
rect 33416 15036 33468 15088
rect 22468 15011 22520 15020
rect 22468 14977 22471 15011
rect 22471 14977 22520 15011
rect 21456 14900 21508 14952
rect 21640 14900 21692 14952
rect 22468 14968 22520 14977
rect 22560 15011 22612 15020
rect 22560 14977 22586 15011
rect 22586 14977 22612 15011
rect 22560 14968 22612 14977
rect 23664 14968 23716 15020
rect 24216 15011 24268 15020
rect 24216 14977 24225 15011
rect 24225 14977 24259 15011
rect 24259 14977 24268 15011
rect 24216 14968 24268 14977
rect 24584 14968 24636 15020
rect 24952 14968 25004 15020
rect 25412 15011 25464 15020
rect 25412 14977 25421 15011
rect 25421 14977 25455 15011
rect 25455 14977 25464 15011
rect 25412 14968 25464 14977
rect 25780 15011 25832 15020
rect 25780 14977 25794 15011
rect 25794 14977 25828 15011
rect 25828 14977 25832 15011
rect 27804 15011 27856 15020
rect 25780 14968 25832 14977
rect 27804 14977 27813 15011
rect 27813 14977 27847 15011
rect 27847 14977 27856 15011
rect 27804 14968 27856 14977
rect 28080 14968 28132 15020
rect 32312 14968 32364 15020
rect 33508 15011 33560 15020
rect 33508 14977 33517 15011
rect 33517 14977 33551 15011
rect 33551 14977 33560 15011
rect 33508 14968 33560 14977
rect 38108 15079 38160 15088
rect 38108 15045 38117 15079
rect 38117 15045 38151 15079
rect 38151 15045 38160 15079
rect 38108 15036 38160 15045
rect 27436 14900 27488 14952
rect 29092 14900 29144 14952
rect 30656 14900 30708 14952
rect 23940 14832 23992 14884
rect 25044 14832 25096 14884
rect 29000 14832 29052 14884
rect 32128 14832 32180 14884
rect 35440 14832 35492 14884
rect 17776 14764 17828 14816
rect 20720 14764 20772 14816
rect 24124 14764 24176 14816
rect 24400 14807 24452 14816
rect 24400 14773 24409 14807
rect 24409 14773 24443 14807
rect 24443 14773 24452 14807
rect 24400 14764 24452 14773
rect 27896 14764 27948 14816
rect 33968 14764 34020 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 13452 14603 13504 14612
rect 13452 14569 13461 14603
rect 13461 14569 13495 14603
rect 13495 14569 13504 14603
rect 13452 14560 13504 14569
rect 16580 14560 16632 14612
rect 19340 14560 19392 14612
rect 19708 14560 19760 14612
rect 25044 14560 25096 14612
rect 25412 14603 25464 14612
rect 25412 14569 25421 14603
rect 25421 14569 25455 14603
rect 25455 14569 25464 14603
rect 25412 14560 25464 14569
rect 27804 14603 27856 14612
rect 27804 14569 27813 14603
rect 27813 14569 27847 14603
rect 27847 14569 27856 14603
rect 27804 14560 27856 14569
rect 28816 14560 28868 14612
rect 15936 14492 15988 14544
rect 6920 14424 6972 14476
rect 7932 14424 7984 14476
rect 7380 14356 7432 14408
rect 12440 14424 12492 14476
rect 11888 14399 11940 14408
rect 11888 14365 11897 14399
rect 11897 14365 11931 14399
rect 11931 14365 11940 14399
rect 11888 14356 11940 14365
rect 12072 14399 12124 14408
rect 12072 14365 12081 14399
rect 12081 14365 12115 14399
rect 12115 14365 12124 14399
rect 12072 14356 12124 14365
rect 13176 14356 13228 14408
rect 12992 14288 13044 14340
rect 14648 14356 14700 14408
rect 16396 14424 16448 14476
rect 17776 14467 17828 14476
rect 16856 14356 16908 14408
rect 17224 14356 17276 14408
rect 17776 14433 17785 14467
rect 17785 14433 17819 14467
rect 17819 14433 17828 14467
rect 17776 14424 17828 14433
rect 18052 14356 18104 14408
rect 20904 14492 20956 14544
rect 24400 14492 24452 14544
rect 20168 14467 20220 14476
rect 20168 14433 20177 14467
rect 20177 14433 20211 14467
rect 20211 14433 20220 14467
rect 20168 14424 20220 14433
rect 22744 14424 22796 14476
rect 15292 14288 15344 14340
rect 17684 14288 17736 14340
rect 18972 14356 19024 14408
rect 19156 14356 19208 14408
rect 21456 14399 21508 14408
rect 21456 14365 21465 14399
rect 21465 14365 21499 14399
rect 21499 14365 21508 14399
rect 21456 14356 21508 14365
rect 21640 14399 21692 14408
rect 21640 14365 21649 14399
rect 21649 14365 21683 14399
rect 21683 14365 21692 14399
rect 21640 14356 21692 14365
rect 21916 14399 21968 14408
rect 21916 14365 21919 14399
rect 21919 14365 21968 14399
rect 21916 14356 21968 14365
rect 22192 14356 22244 14408
rect 23572 14399 23624 14408
rect 23572 14365 23595 14399
rect 23595 14365 23624 14399
rect 23572 14356 23624 14365
rect 23940 14424 23992 14476
rect 24124 14424 24176 14476
rect 35348 14560 35400 14612
rect 37924 14560 37976 14612
rect 35624 14492 35676 14544
rect 24584 14399 24636 14408
rect 24584 14365 24593 14399
rect 24593 14365 24627 14399
rect 24627 14365 24636 14399
rect 24584 14356 24636 14365
rect 25044 14356 25096 14408
rect 33324 14467 33376 14476
rect 33324 14433 33333 14467
rect 33333 14433 33367 14467
rect 33367 14433 33376 14467
rect 33324 14424 33376 14433
rect 34520 14424 34572 14476
rect 35440 14467 35492 14476
rect 35440 14433 35449 14467
rect 35449 14433 35483 14467
rect 35483 14433 35492 14467
rect 35440 14424 35492 14433
rect 23112 14288 23164 14340
rect 23204 14288 23256 14340
rect 25780 14356 25832 14408
rect 27804 14356 27856 14408
rect 28356 14356 28408 14408
rect 29920 14399 29972 14408
rect 27252 14288 27304 14340
rect 29920 14365 29929 14399
rect 29929 14365 29963 14399
rect 29963 14365 29972 14399
rect 29920 14356 29972 14365
rect 33416 14356 33468 14408
rect 35164 14399 35216 14408
rect 35164 14365 35174 14399
rect 35174 14365 35208 14399
rect 35208 14365 35216 14399
rect 35164 14356 35216 14365
rect 35716 14356 35768 14408
rect 37188 14399 37240 14408
rect 37188 14365 37222 14399
rect 37222 14365 37240 14399
rect 37188 14356 37240 14365
rect 32680 14288 32732 14340
rect 33508 14288 33560 14340
rect 17040 14220 17092 14272
rect 18880 14220 18932 14272
rect 19340 14220 19392 14272
rect 19984 14263 20036 14272
rect 19984 14229 19993 14263
rect 19993 14229 20027 14263
rect 20027 14229 20036 14263
rect 19984 14220 20036 14229
rect 20352 14220 20404 14272
rect 22560 14220 22612 14272
rect 23848 14220 23900 14272
rect 24216 14220 24268 14272
rect 25044 14220 25096 14272
rect 29000 14220 29052 14272
rect 30840 14220 30892 14272
rect 34704 14220 34756 14272
rect 36452 14288 36504 14340
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 9312 14059 9364 14068
rect 9312 14025 9321 14059
rect 9321 14025 9355 14059
rect 9355 14025 9364 14059
rect 9312 14016 9364 14025
rect 17868 14016 17920 14068
rect 19432 14016 19484 14068
rect 22744 14059 22796 14068
rect 22744 14025 22753 14059
rect 22753 14025 22787 14059
rect 22787 14025 22796 14059
rect 22744 14016 22796 14025
rect 29920 14016 29972 14068
rect 31668 14016 31720 14068
rect 32772 14059 32824 14068
rect 32772 14025 32781 14059
rect 32781 14025 32815 14059
rect 32815 14025 32824 14059
rect 32772 14016 32824 14025
rect 8392 13948 8444 14000
rect 7932 13923 7984 13932
rect 7932 13889 7941 13923
rect 7941 13889 7975 13923
rect 7975 13889 7984 13923
rect 7932 13880 7984 13889
rect 10600 13923 10652 13932
rect 10600 13889 10609 13923
rect 10609 13889 10643 13923
rect 10643 13889 10652 13923
rect 10600 13880 10652 13889
rect 12072 13948 12124 14000
rect 11888 13923 11940 13932
rect 11888 13889 11897 13923
rect 11897 13889 11931 13923
rect 11931 13889 11940 13923
rect 11888 13880 11940 13889
rect 13636 13948 13688 14000
rect 12992 13923 13044 13932
rect 12992 13889 13001 13923
rect 13001 13889 13035 13923
rect 13035 13889 13044 13923
rect 12992 13880 13044 13889
rect 13268 13880 13320 13932
rect 13544 13880 13596 13932
rect 10692 13855 10744 13864
rect 10692 13821 10701 13855
rect 10701 13821 10735 13855
rect 10735 13821 10744 13855
rect 10692 13812 10744 13821
rect 12716 13812 12768 13864
rect 13176 13812 13228 13864
rect 17960 13948 18012 14000
rect 18696 13948 18748 14000
rect 20260 13948 20312 14000
rect 15016 13880 15068 13932
rect 15384 13923 15436 13932
rect 15384 13889 15393 13923
rect 15393 13889 15427 13923
rect 15427 13889 15436 13923
rect 15384 13880 15436 13889
rect 17224 13923 17276 13932
rect 17224 13889 17233 13923
rect 17233 13889 17267 13923
rect 17267 13889 17276 13923
rect 17224 13880 17276 13889
rect 19340 13880 19392 13932
rect 20076 13880 20128 13932
rect 20352 13880 20404 13932
rect 23940 13948 23992 14000
rect 27160 13991 27212 14000
rect 27160 13957 27169 13991
rect 27169 13957 27203 13991
rect 27203 13957 27212 13991
rect 27160 13948 27212 13957
rect 27252 13948 27304 14000
rect 23204 13923 23256 13932
rect 23204 13889 23213 13923
rect 23213 13889 23247 13923
rect 23247 13889 23256 13923
rect 23204 13880 23256 13889
rect 24216 13923 24268 13932
rect 24216 13889 24225 13923
rect 24225 13889 24259 13923
rect 24259 13889 24268 13923
rect 24216 13880 24268 13889
rect 24584 13880 24636 13932
rect 25044 13923 25096 13932
rect 25044 13889 25053 13923
rect 25053 13889 25087 13923
rect 25087 13889 25096 13923
rect 25044 13880 25096 13889
rect 25872 13880 25924 13932
rect 26332 13923 26384 13932
rect 26332 13889 26341 13923
rect 26341 13889 26375 13923
rect 26375 13889 26384 13923
rect 26332 13880 26384 13889
rect 26976 13880 27028 13932
rect 27988 13923 28040 13932
rect 15200 13855 15252 13864
rect 13728 13744 13780 13796
rect 15200 13821 15209 13855
rect 15209 13821 15243 13855
rect 15243 13821 15252 13855
rect 15200 13812 15252 13821
rect 17408 13812 17460 13864
rect 18328 13812 18380 13864
rect 22744 13812 22796 13864
rect 23480 13812 23532 13864
rect 24124 13855 24176 13864
rect 24124 13821 24133 13855
rect 24133 13821 24167 13855
rect 24167 13821 24176 13855
rect 24124 13812 24176 13821
rect 27988 13889 27997 13923
rect 27997 13889 28031 13923
rect 28031 13889 28040 13923
rect 27988 13880 28040 13889
rect 28816 13923 28868 13932
rect 28816 13889 28825 13923
rect 28825 13889 28859 13923
rect 28859 13889 28868 13923
rect 28816 13880 28868 13889
rect 33508 13948 33560 14000
rect 31116 13880 31168 13932
rect 31208 13880 31260 13932
rect 33048 13923 33100 13932
rect 33048 13889 33057 13923
rect 33057 13889 33091 13923
rect 33091 13889 33100 13923
rect 33048 13880 33100 13889
rect 15108 13744 15160 13796
rect 21364 13744 21416 13796
rect 27620 13812 27672 13864
rect 28632 13812 28684 13864
rect 30380 13855 30432 13864
rect 30380 13821 30389 13855
rect 30389 13821 30423 13855
rect 30423 13821 30432 13855
rect 30380 13812 30432 13821
rect 32864 13812 32916 13864
rect 33324 13855 33376 13864
rect 33324 13821 33333 13855
rect 33333 13821 33367 13855
rect 33367 13821 33376 13855
rect 33324 13812 33376 13821
rect 35532 14016 35584 14068
rect 34796 13948 34848 14000
rect 35716 13948 35768 14000
rect 36452 13991 36504 14000
rect 36452 13957 36461 13991
rect 36461 13957 36495 13991
rect 36495 13957 36504 13991
rect 36452 13948 36504 13957
rect 33968 13880 34020 13932
rect 35164 13880 35216 13932
rect 36176 13880 36228 13932
rect 35348 13812 35400 13864
rect 35624 13812 35676 13864
rect 38292 13855 38344 13864
rect 38292 13821 38301 13855
rect 38301 13821 38335 13855
rect 38335 13821 38344 13855
rect 38292 13812 38344 13821
rect 16028 13676 16080 13728
rect 18144 13676 18196 13728
rect 27804 13744 27856 13796
rect 35808 13787 35860 13796
rect 35808 13753 35817 13787
rect 35817 13753 35851 13787
rect 35851 13753 35860 13787
rect 35808 13744 35860 13753
rect 22836 13676 22888 13728
rect 23388 13676 23440 13728
rect 25044 13676 25096 13728
rect 26976 13676 27028 13728
rect 28172 13719 28224 13728
rect 28172 13685 28181 13719
rect 28181 13685 28215 13719
rect 28215 13685 28224 13719
rect 28172 13676 28224 13685
rect 29184 13676 29236 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 10692 13515 10744 13524
rect 10692 13481 10701 13515
rect 10701 13481 10735 13515
rect 10735 13481 10744 13515
rect 10692 13472 10744 13481
rect 10784 13472 10836 13524
rect 15108 13472 15160 13524
rect 15200 13472 15252 13524
rect 23572 13515 23624 13524
rect 23572 13481 23581 13515
rect 23581 13481 23615 13515
rect 23615 13481 23624 13515
rect 23572 13472 23624 13481
rect 11152 13336 11204 13388
rect 10784 13268 10836 13320
rect 12440 13268 12492 13320
rect 15384 13336 15436 13388
rect 15016 13268 15068 13320
rect 15752 13268 15804 13320
rect 18144 13404 18196 13456
rect 23296 13404 23348 13456
rect 30196 13472 30248 13524
rect 36728 13472 36780 13524
rect 25596 13404 25648 13456
rect 28816 13404 28868 13456
rect 30932 13404 30984 13456
rect 33784 13404 33836 13456
rect 17592 13336 17644 13388
rect 16488 13311 16540 13320
rect 16488 13277 16497 13311
rect 16497 13277 16531 13311
rect 16531 13277 16540 13311
rect 16488 13268 16540 13277
rect 16856 13311 16908 13320
rect 12900 13243 12952 13252
rect 12900 13209 12909 13243
rect 12909 13209 12943 13243
rect 12943 13209 12952 13243
rect 12900 13200 12952 13209
rect 13268 13132 13320 13184
rect 14556 13132 14608 13184
rect 16856 13277 16865 13311
rect 16865 13277 16899 13311
rect 16899 13277 16908 13311
rect 16856 13268 16908 13277
rect 19984 13336 20036 13388
rect 18144 13311 18196 13320
rect 18144 13277 18153 13311
rect 18153 13277 18187 13311
rect 18187 13277 18196 13311
rect 18144 13268 18196 13277
rect 20904 13311 20956 13320
rect 17776 13200 17828 13252
rect 20904 13277 20913 13311
rect 20913 13277 20947 13311
rect 20947 13277 20956 13311
rect 20904 13268 20956 13277
rect 21732 13336 21784 13388
rect 26976 13379 27028 13388
rect 26976 13345 26985 13379
rect 26985 13345 27019 13379
rect 27019 13345 27028 13379
rect 26976 13336 27028 13345
rect 21548 13311 21600 13320
rect 21548 13277 21557 13311
rect 21557 13277 21591 13311
rect 21591 13277 21600 13311
rect 21548 13268 21600 13277
rect 21640 13311 21692 13320
rect 21640 13277 21649 13311
rect 21649 13277 21683 13311
rect 21683 13277 21692 13311
rect 21640 13268 21692 13277
rect 23480 13268 23532 13320
rect 23940 13268 23992 13320
rect 25872 13311 25924 13320
rect 25872 13277 25881 13311
rect 25881 13277 25915 13311
rect 25915 13277 25924 13311
rect 25872 13268 25924 13277
rect 27620 13336 27672 13388
rect 29000 13336 29052 13388
rect 30840 13379 30892 13388
rect 30840 13345 30849 13379
rect 30849 13345 30883 13379
rect 30883 13345 30892 13379
rect 30840 13336 30892 13345
rect 35716 13379 35768 13388
rect 35716 13345 35725 13379
rect 35725 13345 35759 13379
rect 35759 13345 35768 13379
rect 35716 13336 35768 13345
rect 27804 13268 27856 13320
rect 28356 13311 28408 13320
rect 28356 13277 28365 13311
rect 28365 13277 28399 13311
rect 28399 13277 28408 13311
rect 28356 13268 28408 13277
rect 21916 13200 21968 13252
rect 22744 13200 22796 13252
rect 24216 13200 24268 13252
rect 25044 13200 25096 13252
rect 27620 13200 27672 13252
rect 28264 13200 28316 13252
rect 30932 13311 30984 13320
rect 28632 13200 28684 13252
rect 30932 13277 30941 13311
rect 30941 13277 30975 13311
rect 30975 13277 30984 13311
rect 30932 13268 30984 13277
rect 31024 13268 31076 13320
rect 34704 13268 34756 13320
rect 31668 13200 31720 13252
rect 19340 13132 19392 13184
rect 21088 13175 21140 13184
rect 21088 13141 21097 13175
rect 21097 13141 21131 13175
rect 21131 13141 21140 13175
rect 21088 13132 21140 13141
rect 22192 13132 22244 13184
rect 22468 13132 22520 13184
rect 30012 13132 30064 13184
rect 34520 13132 34572 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 7932 12928 7984 12980
rect 11152 12903 11204 12912
rect 11152 12869 11161 12903
rect 11161 12869 11195 12903
rect 11195 12869 11204 12903
rect 11152 12860 11204 12869
rect 12164 12860 12216 12912
rect 12900 12860 12952 12912
rect 12716 12835 12768 12844
rect 9772 12767 9824 12776
rect 9772 12733 9781 12767
rect 9781 12733 9815 12767
rect 9815 12733 9824 12767
rect 9772 12724 9824 12733
rect 12716 12801 12725 12835
rect 12725 12801 12759 12835
rect 12759 12801 12768 12835
rect 12716 12792 12768 12801
rect 13360 12928 13412 12980
rect 14648 12928 14700 12980
rect 16856 12928 16908 12980
rect 17776 12971 17828 12980
rect 17776 12937 17785 12971
rect 17785 12937 17819 12971
rect 17819 12937 17828 12971
rect 17776 12928 17828 12937
rect 21088 12928 21140 12980
rect 13268 12903 13320 12912
rect 13268 12869 13277 12903
rect 13277 12869 13311 12903
rect 13311 12869 13320 12903
rect 13268 12860 13320 12869
rect 13452 12860 13504 12912
rect 14004 12792 14056 12844
rect 14556 12792 14608 12844
rect 15568 12792 15620 12844
rect 16488 12860 16540 12912
rect 15752 12835 15804 12844
rect 15752 12801 15761 12835
rect 15761 12801 15795 12835
rect 15795 12801 15804 12835
rect 15752 12792 15804 12801
rect 17224 12792 17276 12844
rect 17500 12792 17552 12844
rect 19340 12792 19392 12844
rect 19708 12835 19760 12844
rect 14832 12767 14884 12776
rect 12716 12656 12768 12708
rect 13452 12656 13504 12708
rect 13636 12699 13688 12708
rect 13636 12665 13645 12699
rect 13645 12665 13679 12699
rect 13679 12665 13688 12699
rect 13636 12656 13688 12665
rect 14832 12733 14841 12767
rect 14841 12733 14875 12767
rect 14875 12733 14884 12767
rect 14832 12724 14884 12733
rect 19708 12801 19717 12835
rect 19717 12801 19751 12835
rect 19751 12801 19760 12835
rect 19708 12792 19760 12801
rect 19984 12792 20036 12844
rect 21180 12835 21232 12844
rect 21180 12801 21189 12835
rect 21189 12801 21223 12835
rect 21223 12801 21232 12835
rect 21180 12792 21232 12801
rect 21364 12792 21416 12844
rect 22192 12835 22244 12844
rect 22192 12801 22201 12835
rect 22201 12801 22235 12835
rect 22235 12801 22244 12835
rect 22192 12792 22244 12801
rect 25136 12860 25188 12912
rect 29736 12928 29788 12980
rect 32036 12928 32088 12980
rect 25412 12835 25464 12844
rect 25412 12801 25421 12835
rect 25421 12801 25455 12835
rect 25455 12801 25464 12835
rect 25412 12792 25464 12801
rect 25596 12835 25648 12844
rect 25596 12801 25605 12835
rect 25605 12801 25639 12835
rect 25639 12801 25648 12835
rect 25596 12792 25648 12801
rect 27804 12792 27856 12844
rect 29092 12860 29144 12912
rect 20076 12724 20128 12776
rect 21548 12724 21600 12776
rect 22468 12767 22520 12776
rect 22468 12733 22477 12767
rect 22477 12733 22511 12767
rect 22511 12733 22520 12767
rect 22468 12724 22520 12733
rect 27988 12767 28040 12776
rect 27988 12733 27997 12767
rect 27997 12733 28031 12767
rect 28031 12733 28040 12767
rect 27988 12724 28040 12733
rect 28816 12724 28868 12776
rect 29184 12792 29236 12844
rect 33876 12792 33928 12844
rect 16764 12656 16816 12708
rect 17776 12656 17828 12708
rect 32864 12724 32916 12776
rect 33048 12724 33100 12776
rect 9220 12588 9272 12640
rect 12532 12631 12584 12640
rect 12532 12597 12541 12631
rect 12541 12597 12575 12631
rect 12575 12597 12584 12631
rect 12532 12588 12584 12597
rect 14188 12631 14240 12640
rect 14188 12597 14197 12631
rect 14197 12597 14231 12631
rect 14231 12597 14240 12631
rect 14188 12588 14240 12597
rect 15660 12588 15712 12640
rect 19708 12588 19760 12640
rect 20628 12588 20680 12640
rect 21456 12588 21508 12640
rect 27804 12631 27856 12640
rect 27804 12597 27813 12631
rect 27813 12597 27847 12631
rect 27847 12597 27856 12631
rect 27804 12588 27856 12597
rect 32588 12631 32640 12640
rect 32588 12597 32597 12631
rect 32597 12597 32631 12631
rect 32631 12597 32640 12631
rect 32588 12588 32640 12597
rect 35532 12588 35584 12640
rect 38292 12631 38344 12640
rect 38292 12597 38301 12631
rect 38301 12597 38335 12631
rect 38335 12597 38344 12631
rect 38292 12588 38344 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 10600 12384 10652 12436
rect 13176 12427 13228 12436
rect 13176 12393 13185 12427
rect 13185 12393 13219 12427
rect 13219 12393 13228 12427
rect 13176 12384 13228 12393
rect 15016 12427 15068 12436
rect 15016 12393 15025 12427
rect 15025 12393 15059 12427
rect 15059 12393 15068 12427
rect 15016 12384 15068 12393
rect 15660 12384 15712 12436
rect 17040 12384 17092 12436
rect 17592 12384 17644 12436
rect 18788 12384 18840 12436
rect 20168 12384 20220 12436
rect 20720 12384 20772 12436
rect 21180 12384 21232 12436
rect 11796 12316 11848 12368
rect 15384 12316 15436 12368
rect 9220 12291 9272 12300
rect 9220 12257 9229 12291
rect 9229 12257 9263 12291
rect 9263 12257 9272 12291
rect 9220 12248 9272 12257
rect 12624 12248 12676 12300
rect 14188 12248 14240 12300
rect 15568 12291 15620 12300
rect 15568 12257 15577 12291
rect 15577 12257 15611 12291
rect 15611 12257 15620 12291
rect 15568 12248 15620 12257
rect 16396 12248 16448 12300
rect 16948 12248 17000 12300
rect 17224 12291 17276 12300
rect 17224 12257 17233 12291
rect 17233 12257 17267 12291
rect 17267 12257 17276 12291
rect 17224 12248 17276 12257
rect 9312 12223 9364 12232
rect 9312 12189 9321 12223
rect 9321 12189 9355 12223
rect 9355 12189 9364 12223
rect 9312 12180 9364 12189
rect 12348 12180 12400 12232
rect 13268 12180 13320 12232
rect 13452 12180 13504 12232
rect 12440 12112 12492 12164
rect 15660 12112 15712 12164
rect 15476 12087 15528 12096
rect 15476 12053 15485 12087
rect 15485 12053 15519 12087
rect 15519 12053 15528 12087
rect 15476 12044 15528 12053
rect 17040 12180 17092 12232
rect 18788 12223 18840 12232
rect 18788 12189 18797 12223
rect 18797 12189 18831 12223
rect 18831 12189 18840 12223
rect 18788 12180 18840 12189
rect 19064 12180 19116 12232
rect 21548 12316 21600 12368
rect 19708 12223 19760 12232
rect 19708 12189 19717 12223
rect 19717 12189 19751 12223
rect 19751 12189 19760 12223
rect 19708 12180 19760 12189
rect 19340 12112 19392 12164
rect 17684 12044 17736 12096
rect 18880 12044 18932 12096
rect 20076 12180 20128 12232
rect 21640 12248 21692 12300
rect 26332 12384 26384 12436
rect 27988 12384 28040 12436
rect 29000 12427 29052 12436
rect 29000 12393 29009 12427
rect 29009 12393 29043 12427
rect 29043 12393 29052 12427
rect 29000 12384 29052 12393
rect 21916 12223 21968 12232
rect 21916 12189 21925 12223
rect 21925 12189 21959 12223
rect 21959 12189 21968 12223
rect 21916 12180 21968 12189
rect 20444 12112 20496 12164
rect 22284 12180 22336 12232
rect 24860 12223 24912 12232
rect 24860 12189 24869 12223
rect 24869 12189 24903 12223
rect 24903 12189 24912 12223
rect 24860 12180 24912 12189
rect 25964 12291 26016 12300
rect 25964 12257 25973 12291
rect 25973 12257 26007 12291
rect 26007 12257 26016 12291
rect 25964 12248 26016 12257
rect 28448 12248 28500 12300
rect 27620 12180 27672 12232
rect 28264 12223 28316 12232
rect 28264 12189 28273 12223
rect 28273 12189 28307 12223
rect 28307 12189 28316 12223
rect 28264 12180 28316 12189
rect 28632 12180 28684 12232
rect 28816 12248 28868 12300
rect 28908 12180 28960 12232
rect 25780 12112 25832 12164
rect 33232 12384 33284 12436
rect 33876 12427 33928 12436
rect 33876 12393 33885 12427
rect 33885 12393 33919 12427
rect 33919 12393 33928 12427
rect 33876 12384 33928 12393
rect 30840 12248 30892 12300
rect 34428 12248 34480 12300
rect 35716 12248 35768 12300
rect 30380 12180 30432 12232
rect 32496 12223 32548 12232
rect 32496 12189 32505 12223
rect 32505 12189 32539 12223
rect 32539 12189 32548 12223
rect 32496 12180 32548 12189
rect 32588 12180 32640 12232
rect 33048 12180 33100 12232
rect 38200 12180 38252 12232
rect 20812 12044 20864 12096
rect 21364 12044 21416 12096
rect 24768 12087 24820 12096
rect 24768 12053 24777 12087
rect 24777 12053 24811 12087
rect 24811 12053 24820 12087
rect 24768 12044 24820 12053
rect 25872 12087 25924 12096
rect 25872 12053 25881 12087
rect 25881 12053 25915 12087
rect 25915 12053 25924 12087
rect 25872 12044 25924 12053
rect 27804 12044 27856 12096
rect 28264 12044 28316 12096
rect 32036 12112 32088 12164
rect 34336 12112 34388 12164
rect 31116 12087 31168 12096
rect 31116 12053 31125 12087
rect 31125 12053 31159 12087
rect 31159 12053 31168 12087
rect 31116 12044 31168 12053
rect 31484 12087 31536 12096
rect 31484 12053 31493 12087
rect 31493 12053 31527 12087
rect 31527 12053 31536 12087
rect 31484 12044 31536 12053
rect 34796 12044 34848 12096
rect 35808 12112 35860 12164
rect 37464 12112 37516 12164
rect 35716 12044 35768 12096
rect 37832 12044 37884 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 9312 11883 9364 11892
rect 9312 11849 9321 11883
rect 9321 11849 9355 11883
rect 9355 11849 9364 11883
rect 9312 11840 9364 11849
rect 9772 11840 9824 11892
rect 15476 11840 15528 11892
rect 16764 11840 16816 11892
rect 19064 11883 19116 11892
rect 19064 11849 19073 11883
rect 19073 11849 19107 11883
rect 19107 11849 19116 11883
rect 19064 11840 19116 11849
rect 19340 11840 19392 11892
rect 19708 11840 19760 11892
rect 20260 11840 20312 11892
rect 25228 11883 25280 11892
rect 11060 11772 11112 11824
rect 12348 11815 12400 11824
rect 12348 11781 12357 11815
rect 12357 11781 12391 11815
rect 12391 11781 12400 11815
rect 12348 11772 12400 11781
rect 12624 11772 12676 11824
rect 17500 11815 17552 11824
rect 17500 11781 17509 11815
rect 17509 11781 17543 11815
rect 17543 11781 17552 11815
rect 17500 11772 17552 11781
rect 7932 11679 7984 11688
rect 7932 11645 7941 11679
rect 7941 11645 7975 11679
rect 7975 11645 7984 11679
rect 7932 11636 7984 11645
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 10508 11636 10560 11688
rect 15660 11704 15712 11756
rect 17776 11704 17828 11756
rect 21640 11772 21692 11824
rect 19984 11747 20036 11756
rect 15384 11679 15436 11688
rect 15384 11645 15393 11679
rect 15393 11645 15427 11679
rect 15427 11645 15436 11679
rect 15384 11636 15436 11645
rect 19340 11636 19392 11688
rect 19708 11636 19760 11688
rect 19984 11713 19993 11747
rect 19993 11713 20027 11747
rect 20027 11713 20036 11747
rect 19984 11704 20036 11713
rect 20260 11704 20312 11756
rect 22008 11704 22060 11756
rect 23480 11772 23532 11824
rect 25228 11849 25237 11883
rect 25237 11849 25271 11883
rect 25271 11849 25280 11883
rect 25228 11840 25280 11849
rect 25780 11840 25832 11892
rect 34612 11840 34664 11892
rect 37464 11883 37516 11892
rect 37464 11849 37473 11883
rect 37473 11849 37507 11883
rect 37507 11849 37516 11883
rect 37464 11840 37516 11849
rect 37832 11883 37884 11892
rect 37832 11849 37841 11883
rect 37841 11849 37875 11883
rect 37875 11849 37884 11883
rect 37832 11840 37884 11849
rect 25964 11815 26016 11824
rect 25964 11781 25973 11815
rect 25973 11781 26007 11815
rect 26007 11781 26016 11815
rect 25964 11772 26016 11781
rect 26056 11772 26108 11824
rect 31116 11772 31168 11824
rect 11704 11568 11756 11620
rect 17684 11568 17736 11620
rect 21732 11568 21784 11620
rect 24768 11568 24820 11620
rect 30104 11704 30156 11756
rect 30380 11747 30432 11756
rect 30380 11713 30389 11747
rect 30389 11713 30423 11747
rect 30423 11713 30432 11747
rect 30380 11704 30432 11713
rect 30472 11704 30524 11756
rect 33048 11772 33100 11824
rect 32312 11747 32364 11756
rect 32312 11713 32321 11747
rect 32321 11713 32355 11747
rect 32355 11713 32364 11747
rect 32312 11704 32364 11713
rect 32864 11747 32916 11756
rect 32864 11713 32873 11747
rect 32873 11713 32907 11747
rect 32907 11713 32916 11747
rect 32864 11704 32916 11713
rect 33140 11747 33192 11756
rect 33140 11713 33149 11747
rect 33149 11713 33183 11747
rect 33183 11713 33192 11747
rect 33140 11704 33192 11713
rect 33876 11704 33928 11756
rect 34704 11704 34756 11756
rect 35900 11747 35952 11756
rect 35900 11713 35909 11747
rect 35909 11713 35943 11747
rect 35943 11713 35952 11747
rect 35900 11704 35952 11713
rect 25780 11636 25832 11688
rect 26148 11636 26200 11688
rect 26240 11636 26292 11688
rect 31484 11636 31536 11688
rect 35808 11679 35860 11688
rect 35808 11645 35817 11679
rect 35817 11645 35851 11679
rect 35851 11645 35860 11679
rect 35808 11636 35860 11645
rect 10324 11500 10376 11552
rect 11244 11500 11296 11552
rect 11980 11500 12032 11552
rect 26148 11543 26200 11552
rect 26148 11509 26157 11543
rect 26157 11509 26191 11543
rect 26191 11509 26200 11543
rect 26148 11500 26200 11509
rect 29000 11500 29052 11552
rect 31852 11500 31904 11552
rect 36176 11568 36228 11620
rect 35716 11500 35768 11552
rect 38200 11636 38252 11688
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 10784 11296 10836 11348
rect 11060 11296 11112 11348
rect 14832 11296 14884 11348
rect 19984 11296 20036 11348
rect 21456 11296 21508 11348
rect 15752 11228 15804 11280
rect 10324 11135 10376 11144
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 11060 11092 11112 11144
rect 11244 11135 11296 11144
rect 11244 11101 11253 11135
rect 11253 11101 11287 11135
rect 11287 11101 11296 11135
rect 11244 11092 11296 11101
rect 12348 11092 12400 11144
rect 12624 11092 12676 11144
rect 14004 11092 14056 11144
rect 15384 11092 15436 11144
rect 10508 10999 10560 11008
rect 10508 10965 10517 10999
rect 10517 10965 10551 10999
rect 10551 10965 10560 10999
rect 10508 10956 10560 10965
rect 12440 10999 12492 11008
rect 12440 10965 12449 10999
rect 12449 10965 12483 10999
rect 12483 10965 12492 10999
rect 12440 10956 12492 10965
rect 13360 10956 13412 11008
rect 17776 11228 17828 11280
rect 18052 11271 18104 11280
rect 18052 11237 18061 11271
rect 18061 11237 18095 11271
rect 18095 11237 18104 11271
rect 18052 11228 18104 11237
rect 18604 11228 18656 11280
rect 19340 11160 19392 11212
rect 16856 11024 16908 11076
rect 17592 11092 17644 11144
rect 20168 11160 20220 11212
rect 18512 11024 18564 11076
rect 18972 11024 19024 11076
rect 20444 11092 20496 11144
rect 22468 11160 22520 11212
rect 22928 11160 22980 11212
rect 25228 11160 25280 11212
rect 21640 11092 21692 11144
rect 26700 11135 26752 11144
rect 26700 11101 26709 11135
rect 26709 11101 26743 11135
rect 26743 11101 26752 11135
rect 26700 11092 26752 11101
rect 27252 11092 27304 11144
rect 30840 11296 30892 11348
rect 34428 11296 34480 11348
rect 35808 11296 35860 11348
rect 28908 11228 28960 11280
rect 25964 11024 26016 11076
rect 27160 11024 27212 11076
rect 15292 10956 15344 11008
rect 16948 10956 17000 11008
rect 17224 10999 17276 11008
rect 17224 10965 17233 10999
rect 17233 10965 17267 10999
rect 17267 10965 17276 10999
rect 17224 10956 17276 10965
rect 18236 10999 18288 11008
rect 18236 10965 18245 10999
rect 18245 10965 18279 10999
rect 18279 10965 18288 10999
rect 18236 10956 18288 10965
rect 22008 10956 22060 11008
rect 24860 10956 24912 11008
rect 28080 10999 28132 11008
rect 28080 10965 28089 10999
rect 28089 10965 28123 10999
rect 28123 10965 28132 10999
rect 29184 11092 29236 11144
rect 30288 11092 30340 11144
rect 33140 11228 33192 11280
rect 33600 11228 33652 11280
rect 32496 11160 32548 11212
rect 32956 11160 33008 11212
rect 31392 11135 31444 11144
rect 30104 11024 30156 11076
rect 31392 11101 31401 11135
rect 31401 11101 31435 11135
rect 31435 11101 31444 11135
rect 31392 11092 31444 11101
rect 33232 11024 33284 11076
rect 34796 11024 34848 11076
rect 37464 11024 37516 11076
rect 28080 10956 28132 10965
rect 37832 10956 37884 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 17224 10752 17276 10804
rect 18512 10795 18564 10804
rect 18512 10761 18521 10795
rect 18521 10761 18555 10795
rect 18555 10761 18564 10795
rect 18512 10752 18564 10761
rect 24952 10752 25004 10804
rect 25964 10795 26016 10804
rect 25964 10761 25973 10795
rect 25973 10761 26007 10795
rect 26007 10761 26016 10795
rect 25964 10752 26016 10761
rect 27160 10795 27212 10804
rect 27160 10761 27169 10795
rect 27169 10761 27203 10795
rect 27203 10761 27212 10795
rect 27160 10752 27212 10761
rect 28080 10752 28132 10804
rect 30104 10795 30156 10804
rect 30104 10761 30113 10795
rect 30113 10761 30147 10795
rect 30147 10761 30156 10795
rect 30104 10752 30156 10761
rect 37464 10795 37516 10804
rect 37464 10761 37473 10795
rect 37473 10761 37507 10795
rect 37507 10761 37516 10795
rect 37464 10752 37516 10761
rect 17684 10727 17736 10736
rect 17684 10693 17693 10727
rect 17693 10693 17727 10727
rect 17727 10693 17736 10727
rect 17684 10684 17736 10693
rect 21456 10684 21508 10736
rect 11796 10659 11848 10668
rect 11796 10625 11805 10659
rect 11805 10625 11839 10659
rect 11839 10625 11848 10659
rect 11796 10616 11848 10625
rect 11980 10659 12032 10668
rect 11980 10625 11989 10659
rect 11989 10625 12023 10659
rect 12023 10625 12032 10659
rect 11980 10616 12032 10625
rect 13176 10659 13228 10668
rect 13176 10625 13185 10659
rect 13185 10625 13219 10659
rect 13219 10625 13228 10659
rect 13176 10616 13228 10625
rect 13360 10659 13412 10668
rect 13360 10625 13369 10659
rect 13369 10625 13403 10659
rect 13403 10625 13412 10659
rect 13360 10616 13412 10625
rect 15476 10616 15528 10668
rect 15660 10616 15712 10668
rect 18052 10616 18104 10668
rect 20812 10616 20864 10668
rect 22008 10659 22060 10668
rect 18236 10548 18288 10600
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 22192 10659 22244 10668
rect 22192 10625 22201 10659
rect 22201 10625 22235 10659
rect 22235 10625 22244 10659
rect 22192 10616 22244 10625
rect 22376 10659 22428 10668
rect 22376 10625 22385 10659
rect 22385 10625 22419 10659
rect 22419 10625 22428 10659
rect 22376 10616 22428 10625
rect 17776 10480 17828 10532
rect 11244 10412 11296 10464
rect 13544 10455 13596 10464
rect 13544 10421 13553 10455
rect 13553 10421 13587 10455
rect 13587 10421 13596 10455
rect 13544 10412 13596 10421
rect 15384 10455 15436 10464
rect 15384 10421 15393 10455
rect 15393 10421 15427 10455
rect 15427 10421 15436 10455
rect 15384 10412 15436 10421
rect 17408 10412 17460 10464
rect 17500 10412 17552 10464
rect 20720 10455 20772 10464
rect 20720 10421 20729 10455
rect 20729 10421 20763 10455
rect 20763 10421 20772 10455
rect 20720 10412 20772 10421
rect 23480 10548 23532 10600
rect 26700 10684 26752 10736
rect 29000 10727 29052 10736
rect 24860 10659 24912 10668
rect 24860 10625 24894 10659
rect 24894 10625 24912 10659
rect 24860 10616 24912 10625
rect 26240 10616 26292 10668
rect 27528 10616 27580 10668
rect 29000 10693 29034 10727
rect 29034 10693 29052 10727
rect 29000 10684 29052 10693
rect 34244 10659 34296 10668
rect 34244 10625 34253 10659
rect 34253 10625 34287 10659
rect 34287 10625 34296 10659
rect 34244 10616 34296 10625
rect 27252 10548 27304 10600
rect 22652 10412 22704 10464
rect 25688 10412 25740 10464
rect 33324 10548 33376 10600
rect 38016 10684 38068 10736
rect 37372 10616 37424 10668
rect 37832 10659 37884 10668
rect 37832 10625 37841 10659
rect 37841 10625 37875 10659
rect 37875 10625 37884 10659
rect 37832 10616 37884 10625
rect 34428 10591 34480 10600
rect 34428 10557 34437 10591
rect 34437 10557 34471 10591
rect 34471 10557 34480 10591
rect 34428 10548 34480 10557
rect 38200 10548 38252 10600
rect 33508 10412 33560 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 10692 10251 10744 10260
rect 10692 10217 10701 10251
rect 10701 10217 10735 10251
rect 10735 10217 10744 10251
rect 10692 10208 10744 10217
rect 12532 10208 12584 10260
rect 12900 10208 12952 10260
rect 13360 10208 13412 10260
rect 20536 10208 20588 10260
rect 22192 10208 22244 10260
rect 24860 10251 24912 10260
rect 24860 10217 24869 10251
rect 24869 10217 24903 10251
rect 24903 10217 24912 10251
rect 24860 10208 24912 10217
rect 25872 10208 25924 10260
rect 32312 10208 32364 10260
rect 14832 10140 14884 10192
rect 21732 10140 21784 10192
rect 22376 10140 22428 10192
rect 34244 10140 34296 10192
rect 7932 10072 7984 10124
rect 13268 10115 13320 10124
rect 13268 10081 13277 10115
rect 13277 10081 13311 10115
rect 13311 10081 13320 10115
rect 13268 10072 13320 10081
rect 14464 10072 14516 10124
rect 10876 10004 10928 10056
rect 11244 10047 11296 10056
rect 11244 10013 11253 10047
rect 11253 10013 11287 10047
rect 11287 10013 11296 10047
rect 11244 10004 11296 10013
rect 13176 10047 13228 10056
rect 11428 9979 11480 9988
rect 11428 9945 11437 9979
rect 11437 9945 11471 9979
rect 11471 9945 11480 9979
rect 11428 9936 11480 9945
rect 13176 10013 13185 10047
rect 13185 10013 13219 10047
rect 13219 10013 13228 10047
rect 13176 10004 13228 10013
rect 20352 10072 20404 10124
rect 26332 10072 26384 10124
rect 26700 10072 26752 10124
rect 32956 10115 33008 10124
rect 32956 10081 32965 10115
rect 32965 10081 32999 10115
rect 32999 10081 33008 10115
rect 32956 10072 33008 10081
rect 34520 10140 34572 10192
rect 36176 10115 36228 10124
rect 36176 10081 36185 10115
rect 36185 10081 36219 10115
rect 36219 10081 36228 10115
rect 36176 10072 36228 10081
rect 15384 10047 15436 10056
rect 15384 10013 15393 10047
rect 15393 10013 15427 10047
rect 15427 10013 15436 10047
rect 15384 10004 15436 10013
rect 16764 10047 16816 10056
rect 16764 10013 16773 10047
rect 16773 10013 16807 10047
rect 16807 10013 16816 10047
rect 16764 10004 16816 10013
rect 17408 10047 17460 10056
rect 17408 10013 17417 10047
rect 17417 10013 17451 10047
rect 17451 10013 17460 10047
rect 17408 10004 17460 10013
rect 18696 10047 18748 10056
rect 18696 10013 18705 10047
rect 18705 10013 18739 10047
rect 18739 10013 18748 10047
rect 18696 10004 18748 10013
rect 11336 9911 11388 9920
rect 11336 9877 11345 9911
rect 11345 9877 11379 9911
rect 11379 9877 11388 9911
rect 11336 9868 11388 9877
rect 12440 9868 12492 9920
rect 16948 9936 17000 9988
rect 15660 9868 15712 9920
rect 17500 9911 17552 9920
rect 17500 9877 17509 9911
rect 17509 9877 17543 9911
rect 17543 9877 17552 9911
rect 17500 9868 17552 9877
rect 20812 10004 20864 10056
rect 21456 10004 21508 10056
rect 22468 10047 22520 10056
rect 22468 10013 22477 10047
rect 22477 10013 22511 10047
rect 22511 10013 22520 10047
rect 22468 10004 22520 10013
rect 22652 10047 22704 10056
rect 22652 10013 22661 10047
rect 22661 10013 22695 10047
rect 22695 10013 22704 10047
rect 22652 10004 22704 10013
rect 24768 10047 24820 10056
rect 24768 10013 24777 10047
rect 24777 10013 24811 10047
rect 24811 10013 24820 10047
rect 24768 10004 24820 10013
rect 32128 10047 32180 10056
rect 32128 10013 32137 10047
rect 32137 10013 32171 10047
rect 32171 10013 32180 10047
rect 32128 10004 32180 10013
rect 22100 9936 22152 9988
rect 26240 9936 26292 9988
rect 31944 9936 31996 9988
rect 33508 10004 33560 10056
rect 34520 10004 34572 10056
rect 35900 10047 35952 10056
rect 35900 10013 35909 10047
rect 35909 10013 35943 10047
rect 35943 10013 35952 10047
rect 35900 10004 35952 10013
rect 37372 10072 37424 10124
rect 38108 10115 38160 10124
rect 38108 10081 38117 10115
rect 38117 10081 38151 10115
rect 38151 10081 38160 10115
rect 38108 10072 38160 10081
rect 37832 10047 37884 10056
rect 37832 10013 37841 10047
rect 37841 10013 37875 10047
rect 37875 10013 37884 10047
rect 37832 10004 37884 10013
rect 33416 9936 33468 9988
rect 33600 9936 33652 9988
rect 32772 9868 32824 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 12440 9664 12492 9716
rect 15384 9664 15436 9716
rect 14740 9596 14792 9648
rect 14924 9596 14976 9648
rect 11428 9528 11480 9580
rect 11796 9528 11848 9580
rect 11244 9460 11296 9512
rect 11336 9460 11388 9512
rect 11060 9392 11112 9444
rect 11704 9435 11756 9444
rect 11704 9401 11713 9435
rect 11713 9401 11747 9435
rect 11747 9401 11756 9435
rect 11704 9392 11756 9401
rect 12164 9571 12216 9580
rect 12164 9537 12173 9571
rect 12173 9537 12207 9571
rect 12207 9537 12216 9571
rect 12164 9528 12216 9537
rect 15660 9528 15712 9580
rect 12440 9503 12492 9512
rect 12440 9469 12449 9503
rect 12449 9469 12483 9503
rect 12483 9469 12492 9503
rect 12992 9503 13044 9512
rect 12440 9460 12492 9469
rect 12992 9469 13001 9503
rect 13001 9469 13035 9503
rect 13035 9469 13044 9503
rect 12992 9460 13044 9469
rect 18052 9460 18104 9512
rect 18420 9528 18472 9580
rect 19156 9571 19208 9580
rect 19156 9537 19165 9571
rect 19165 9537 19199 9571
rect 19199 9537 19208 9571
rect 19156 9528 19208 9537
rect 21088 9571 21140 9580
rect 21088 9537 21097 9571
rect 21097 9537 21131 9571
rect 21131 9537 21140 9571
rect 21088 9528 21140 9537
rect 21272 9528 21324 9580
rect 22284 9528 22336 9580
rect 19892 9460 19944 9512
rect 22468 9460 22520 9512
rect 11980 9324 12032 9376
rect 14648 9324 14700 9376
rect 15568 9324 15620 9376
rect 18328 9324 18380 9376
rect 18420 9324 18472 9376
rect 22560 9392 22612 9444
rect 20536 9324 20588 9376
rect 23480 9596 23532 9648
rect 24860 9664 24912 9716
rect 24768 9596 24820 9648
rect 25228 9596 25280 9648
rect 26240 9664 26292 9716
rect 33232 9664 33284 9716
rect 33600 9707 33652 9716
rect 33600 9673 33609 9707
rect 33609 9673 33643 9707
rect 33643 9673 33652 9707
rect 33600 9664 33652 9673
rect 26424 9596 26476 9648
rect 29184 9639 29236 9648
rect 29184 9605 29193 9639
rect 29193 9605 29227 9639
rect 29227 9605 29236 9639
rect 29184 9596 29236 9605
rect 30196 9596 30248 9648
rect 30840 9639 30892 9648
rect 25320 9460 25372 9512
rect 26700 9528 26752 9580
rect 27988 9528 28040 9580
rect 28356 9392 28408 9444
rect 29644 9571 29696 9580
rect 29644 9537 29653 9571
rect 29653 9537 29687 9571
rect 29687 9537 29696 9571
rect 29828 9571 29880 9580
rect 29644 9528 29696 9537
rect 29828 9537 29837 9571
rect 29837 9537 29871 9571
rect 29871 9537 29880 9571
rect 29828 9528 29880 9537
rect 30288 9571 30340 9580
rect 30288 9537 30297 9571
rect 30297 9537 30331 9571
rect 30331 9537 30340 9571
rect 30288 9528 30340 9537
rect 30840 9605 30849 9639
rect 30849 9605 30883 9639
rect 30883 9605 30892 9639
rect 30840 9596 30892 9605
rect 32128 9596 32180 9648
rect 32588 9596 32640 9648
rect 32772 9596 32824 9648
rect 38108 9639 38160 9648
rect 32036 9528 32088 9580
rect 34152 9571 34204 9580
rect 34152 9537 34161 9571
rect 34161 9537 34195 9571
rect 34195 9537 34204 9571
rect 34152 9528 34204 9537
rect 38108 9605 38117 9639
rect 38117 9605 38151 9639
rect 38151 9605 38160 9639
rect 38108 9596 38160 9605
rect 35532 9528 35584 9580
rect 37832 9571 37884 9580
rect 37832 9537 37841 9571
rect 37841 9537 37875 9571
rect 37875 9537 37884 9571
rect 37832 9528 37884 9537
rect 30748 9460 30800 9512
rect 32772 9503 32824 9512
rect 29920 9392 29972 9444
rect 32772 9469 32781 9503
rect 32781 9469 32815 9503
rect 32815 9469 32824 9503
rect 32772 9460 32824 9469
rect 31760 9324 31812 9376
rect 34152 9324 34204 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 10876 9163 10928 9172
rect 10876 9129 10885 9163
rect 10885 9129 10919 9163
rect 10919 9129 10928 9163
rect 10876 9120 10928 9129
rect 17132 9120 17184 9172
rect 16764 9052 16816 9104
rect 11060 8984 11112 9036
rect 12164 8984 12216 9036
rect 12532 8984 12584 9036
rect 12900 8984 12952 9036
rect 13544 8984 13596 9036
rect 17316 8984 17368 9036
rect 11336 8916 11388 8968
rect 14464 8959 14516 8968
rect 14464 8925 14473 8959
rect 14473 8925 14507 8959
rect 14507 8925 14516 8959
rect 14464 8916 14516 8925
rect 14648 8959 14700 8968
rect 14648 8925 14657 8959
rect 14657 8925 14691 8959
rect 14691 8925 14700 8959
rect 14648 8916 14700 8925
rect 15660 8959 15712 8968
rect 15660 8925 15669 8959
rect 15669 8925 15703 8959
rect 15703 8925 15712 8959
rect 15660 8916 15712 8925
rect 16764 8959 16816 8968
rect 16764 8925 16773 8959
rect 16773 8925 16807 8959
rect 16807 8925 16816 8959
rect 16764 8916 16816 8925
rect 18420 9052 18472 9104
rect 20812 9095 20864 9104
rect 18788 8984 18840 9036
rect 17868 8916 17920 8968
rect 18512 8959 18564 8968
rect 18512 8925 18521 8959
rect 18521 8925 18555 8959
rect 18555 8925 18564 8959
rect 20812 9061 20821 9095
rect 20821 9061 20855 9095
rect 20855 9061 20864 9095
rect 20812 9052 20864 9061
rect 26332 9120 26384 9172
rect 27988 9163 28040 9172
rect 27988 9129 27997 9163
rect 27997 9129 28031 9163
rect 28031 9129 28040 9163
rect 27988 9120 28040 9129
rect 29552 9120 29604 9172
rect 31484 9120 31536 9172
rect 32588 9163 32640 9172
rect 32588 9129 32597 9163
rect 32597 9129 32631 9163
rect 32631 9129 32640 9163
rect 32588 9120 32640 9129
rect 33416 9163 33468 9172
rect 33416 9129 33425 9163
rect 33425 9129 33459 9163
rect 33459 9129 33468 9163
rect 33416 9120 33468 9129
rect 29644 9052 29696 9104
rect 35348 9052 35400 9104
rect 36176 9052 36228 9104
rect 20168 8984 20220 9036
rect 21916 8984 21968 9036
rect 25228 8984 25280 9036
rect 25688 9027 25740 9036
rect 25688 8993 25697 9027
rect 25697 8993 25731 9027
rect 25731 8993 25740 9027
rect 25688 8984 25740 8993
rect 26056 8984 26108 9036
rect 18512 8916 18564 8925
rect 14924 8848 14976 8900
rect 18880 8891 18932 8900
rect 18880 8857 18889 8891
rect 18889 8857 18923 8891
rect 18923 8857 18932 8891
rect 18880 8848 18932 8857
rect 19248 8848 19300 8900
rect 24216 8916 24268 8968
rect 25872 8916 25924 8968
rect 27528 8984 27580 9036
rect 36084 9027 36136 9036
rect 28356 8959 28408 8968
rect 28356 8925 28365 8959
rect 28365 8925 28399 8959
rect 28399 8925 28408 8959
rect 28356 8916 28408 8925
rect 36084 8993 36093 9027
rect 36093 8993 36127 9027
rect 36127 8993 36136 9027
rect 36084 8984 36136 8993
rect 21088 8891 21140 8900
rect 12716 8780 12768 8832
rect 16304 8823 16356 8832
rect 16304 8789 16313 8823
rect 16313 8789 16347 8823
rect 16347 8789 16356 8823
rect 16304 8780 16356 8789
rect 17868 8780 17920 8832
rect 21088 8857 21097 8891
rect 21097 8857 21131 8891
rect 21131 8857 21140 8891
rect 21088 8848 21140 8857
rect 21272 8891 21324 8900
rect 21272 8857 21281 8891
rect 21281 8857 21315 8891
rect 21315 8857 21324 8891
rect 21272 8848 21324 8857
rect 26148 8848 26200 8900
rect 19892 8823 19944 8832
rect 19892 8789 19901 8823
rect 19901 8789 19935 8823
rect 19935 8789 19944 8823
rect 25044 8823 25096 8832
rect 19892 8780 19944 8789
rect 25044 8789 25053 8823
rect 25053 8789 25087 8823
rect 25087 8789 25096 8823
rect 25044 8780 25096 8789
rect 25320 8780 25372 8832
rect 28448 8780 28500 8832
rect 30196 8916 30248 8968
rect 31208 8959 31260 8968
rect 31208 8925 31217 8959
rect 31217 8925 31251 8959
rect 31251 8925 31260 8959
rect 31208 8916 31260 8925
rect 31760 8916 31812 8968
rect 32864 8916 32916 8968
rect 35440 8959 35492 8968
rect 35440 8925 35449 8959
rect 35449 8925 35483 8959
rect 35483 8925 35492 8959
rect 35440 8916 35492 8925
rect 35900 8916 35952 8968
rect 30472 8848 30524 8900
rect 30932 8848 30984 8900
rect 33876 8848 33928 8900
rect 37740 8848 37792 8900
rect 31392 8780 31444 8832
rect 31484 8780 31536 8832
rect 38108 8891 38160 8900
rect 38108 8857 38117 8891
rect 38117 8857 38151 8891
rect 38151 8857 38160 8891
rect 38108 8848 38160 8857
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 12440 8576 12492 8628
rect 14464 8576 14516 8628
rect 11796 8483 11848 8492
rect 11796 8449 11805 8483
rect 11805 8449 11839 8483
rect 11839 8449 11848 8483
rect 11796 8440 11848 8449
rect 12808 8440 12860 8492
rect 14924 8508 14976 8560
rect 25872 8619 25924 8628
rect 18512 8551 18564 8560
rect 14832 8483 14884 8492
rect 14832 8449 14841 8483
rect 14841 8449 14875 8483
rect 14875 8449 14884 8483
rect 14832 8440 14884 8449
rect 14464 8372 14516 8424
rect 18512 8517 18521 8551
rect 18521 8517 18555 8551
rect 18555 8517 18564 8551
rect 18512 8508 18564 8517
rect 25872 8585 25881 8619
rect 25881 8585 25915 8619
rect 25915 8585 25924 8619
rect 25872 8576 25924 8585
rect 27528 8576 27580 8628
rect 29184 8576 29236 8628
rect 31392 8619 31444 8628
rect 25044 8508 25096 8560
rect 28448 8508 28500 8560
rect 30748 8508 30800 8560
rect 31392 8585 31401 8619
rect 31401 8585 31435 8619
rect 31435 8585 31444 8619
rect 31392 8576 31444 8585
rect 32772 8576 32824 8628
rect 36084 8576 36136 8628
rect 37740 8576 37792 8628
rect 15568 8304 15620 8356
rect 16764 8440 16816 8492
rect 16488 8372 16540 8424
rect 18880 8440 18932 8492
rect 20720 8440 20772 8492
rect 18788 8372 18840 8424
rect 20536 8415 20588 8424
rect 20536 8381 20545 8415
rect 20545 8381 20579 8415
rect 20579 8381 20588 8415
rect 20536 8372 20588 8381
rect 20904 8372 20956 8424
rect 19984 8304 20036 8356
rect 23480 8440 23532 8492
rect 27896 8440 27948 8492
rect 29184 8440 29236 8492
rect 29644 8440 29696 8492
rect 30196 8440 30248 8492
rect 30932 8483 30984 8492
rect 30932 8449 30941 8483
rect 30941 8449 30975 8483
rect 30975 8449 30984 8483
rect 30932 8440 30984 8449
rect 33876 8508 33928 8560
rect 32680 8440 32732 8492
rect 32864 8483 32916 8492
rect 32864 8449 32873 8483
rect 32873 8449 32907 8483
rect 32907 8449 32916 8483
rect 32864 8440 32916 8449
rect 33968 8483 34020 8492
rect 33968 8449 33977 8483
rect 33977 8449 34011 8483
rect 34011 8449 34020 8483
rect 33968 8440 34020 8449
rect 35348 8440 35400 8492
rect 25688 8372 25740 8424
rect 26516 8372 26568 8424
rect 14188 8279 14240 8288
rect 14188 8245 14197 8279
rect 14197 8245 14231 8279
rect 14231 8245 14240 8279
rect 14188 8236 14240 8245
rect 18696 8236 18748 8288
rect 28356 8372 28408 8424
rect 31392 8372 31444 8424
rect 31852 8372 31904 8424
rect 34796 8415 34848 8424
rect 29552 8304 29604 8356
rect 34796 8381 34805 8415
rect 34805 8381 34839 8415
rect 34839 8381 34848 8415
rect 34796 8372 34848 8381
rect 37924 8415 37976 8424
rect 37924 8381 37933 8415
rect 37933 8381 37967 8415
rect 37967 8381 37976 8415
rect 37924 8372 37976 8381
rect 38200 8372 38252 8424
rect 34612 8304 34664 8356
rect 37188 8304 37240 8356
rect 27160 8279 27212 8288
rect 27160 8245 27169 8279
rect 27169 8245 27203 8279
rect 27203 8245 27212 8279
rect 27160 8236 27212 8245
rect 32496 8279 32548 8288
rect 32496 8245 32505 8279
rect 32505 8245 32539 8279
rect 32539 8245 32548 8279
rect 32496 8236 32548 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 11796 8075 11848 8084
rect 11796 8041 11805 8075
rect 11805 8041 11839 8075
rect 11839 8041 11848 8075
rect 11796 8032 11848 8041
rect 12808 8075 12860 8084
rect 12808 8041 12817 8075
rect 12817 8041 12851 8075
rect 12851 8041 12860 8075
rect 12808 8032 12860 8041
rect 15568 8075 15620 8084
rect 15568 8041 15577 8075
rect 15577 8041 15611 8075
rect 15611 8041 15620 8075
rect 15568 8032 15620 8041
rect 16672 8032 16724 8084
rect 18788 8032 18840 8084
rect 20904 8032 20956 8084
rect 23020 8075 23072 8084
rect 23020 8041 23029 8075
rect 23029 8041 23063 8075
rect 23063 8041 23072 8075
rect 23020 8032 23072 8041
rect 27896 8075 27948 8084
rect 27896 8041 27905 8075
rect 27905 8041 27939 8075
rect 27939 8041 27948 8075
rect 27896 8032 27948 8041
rect 29828 8032 29880 8084
rect 32864 8032 32916 8084
rect 35348 8032 35400 8084
rect 37832 8032 37884 8084
rect 31668 7964 31720 8016
rect 34428 7964 34480 8016
rect 12256 7871 12308 7880
rect 12256 7837 12265 7871
rect 12265 7837 12299 7871
rect 12299 7837 12308 7871
rect 12256 7828 12308 7837
rect 12716 7871 12768 7880
rect 12716 7837 12725 7871
rect 12725 7837 12759 7871
rect 12759 7837 12768 7871
rect 12716 7828 12768 7837
rect 12900 7803 12952 7812
rect 12900 7769 12909 7803
rect 12909 7769 12943 7803
rect 12943 7769 12952 7803
rect 12900 7760 12952 7769
rect 14188 7828 14240 7880
rect 14832 7896 14884 7948
rect 14924 7871 14976 7880
rect 14924 7837 14933 7871
rect 14933 7837 14967 7871
rect 14967 7837 14976 7871
rect 14924 7828 14976 7837
rect 16304 7828 16356 7880
rect 16488 7871 16540 7880
rect 16488 7837 16497 7871
rect 16497 7837 16531 7871
rect 16531 7837 16540 7871
rect 16672 7871 16724 7880
rect 16488 7828 16540 7837
rect 16672 7837 16681 7871
rect 16681 7837 16715 7871
rect 16715 7837 16724 7871
rect 16672 7828 16724 7837
rect 16856 7828 16908 7880
rect 18604 7896 18656 7948
rect 20628 7896 20680 7948
rect 18420 7871 18472 7880
rect 14740 7803 14792 7812
rect 14740 7769 14749 7803
rect 14749 7769 14783 7803
rect 14783 7769 14792 7803
rect 14740 7760 14792 7769
rect 18420 7837 18429 7871
rect 18429 7837 18463 7871
rect 18463 7837 18472 7871
rect 18420 7828 18472 7837
rect 18696 7871 18748 7880
rect 18696 7837 18705 7871
rect 18705 7837 18739 7871
rect 18739 7837 18748 7871
rect 18696 7828 18748 7837
rect 20536 7871 20588 7880
rect 20536 7837 20545 7871
rect 20545 7837 20579 7871
rect 20579 7837 20588 7871
rect 35256 7896 35308 7948
rect 35348 7896 35400 7948
rect 35532 7896 35584 7948
rect 20536 7828 20588 7837
rect 22468 7828 22520 7880
rect 26608 7828 26660 7880
rect 27160 7828 27212 7880
rect 27896 7828 27948 7880
rect 31208 7828 31260 7880
rect 31668 7828 31720 7880
rect 33232 7871 33284 7880
rect 20812 7760 20864 7812
rect 16212 7735 16264 7744
rect 16212 7701 16221 7735
rect 16221 7701 16255 7735
rect 16255 7701 16264 7735
rect 16212 7692 16264 7701
rect 16580 7692 16632 7744
rect 20260 7692 20312 7744
rect 21732 7760 21784 7812
rect 28356 7803 28408 7812
rect 28356 7769 28365 7803
rect 28365 7769 28399 7803
rect 28399 7769 28408 7803
rect 28356 7760 28408 7769
rect 32496 7760 32548 7812
rect 33232 7837 33241 7871
rect 33241 7837 33275 7871
rect 33275 7837 33284 7871
rect 33232 7828 33284 7837
rect 34796 7760 34848 7812
rect 36728 7828 36780 7880
rect 37188 7871 37240 7880
rect 37188 7837 37222 7871
rect 37222 7837 37240 7871
rect 37188 7828 37240 7837
rect 36084 7760 36136 7812
rect 34612 7692 34664 7744
rect 35164 7692 35216 7744
rect 35256 7692 35308 7744
rect 35900 7692 35952 7744
rect 37924 7692 37976 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 20536 7488 20588 7540
rect 22560 7488 22612 7540
rect 26056 7488 26108 7540
rect 33968 7488 34020 7540
rect 34520 7531 34572 7540
rect 34520 7497 34529 7531
rect 34529 7497 34563 7531
rect 34563 7497 34572 7531
rect 34520 7488 34572 7497
rect 37832 7531 37884 7540
rect 13360 7463 13412 7472
rect 13360 7429 13369 7463
rect 13369 7429 13403 7463
rect 13403 7429 13412 7463
rect 13360 7420 13412 7429
rect 12992 7352 13044 7404
rect 15936 7420 15988 7472
rect 14372 7395 14424 7404
rect 14372 7361 14381 7395
rect 14381 7361 14415 7395
rect 14415 7361 14424 7395
rect 14372 7352 14424 7361
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14740 7395 14792 7404
rect 14464 7352 14516 7361
rect 14740 7361 14749 7395
rect 14749 7361 14783 7395
rect 14783 7361 14792 7395
rect 14740 7352 14792 7361
rect 18696 7420 18748 7472
rect 11980 7327 12032 7336
rect 11980 7293 11989 7327
rect 11989 7293 12023 7327
rect 12023 7293 12032 7327
rect 11980 7284 12032 7293
rect 14188 7284 14240 7336
rect 18604 7352 18656 7404
rect 20812 7420 20864 7472
rect 24032 7463 24084 7472
rect 24032 7429 24041 7463
rect 24041 7429 24075 7463
rect 24075 7429 24084 7463
rect 24032 7420 24084 7429
rect 29184 7420 29236 7472
rect 20260 7395 20312 7404
rect 20260 7361 20269 7395
rect 20269 7361 20303 7395
rect 20303 7361 20312 7395
rect 20260 7352 20312 7361
rect 20628 7395 20680 7404
rect 18144 7327 18196 7336
rect 18144 7293 18153 7327
rect 18153 7293 18187 7327
rect 18187 7293 18196 7327
rect 18144 7284 18196 7293
rect 18788 7327 18840 7336
rect 18788 7293 18797 7327
rect 18797 7293 18831 7327
rect 18831 7293 18840 7327
rect 18788 7284 18840 7293
rect 12900 7216 12952 7268
rect 17960 7216 18012 7268
rect 20628 7361 20637 7395
rect 20637 7361 20671 7395
rect 20671 7361 20680 7395
rect 20628 7352 20680 7361
rect 20904 7352 20956 7404
rect 29644 7395 29696 7404
rect 29644 7361 29653 7395
rect 29653 7361 29687 7395
rect 29687 7361 29696 7395
rect 29644 7352 29696 7361
rect 31668 7352 31720 7404
rect 32956 7352 33008 7404
rect 37832 7497 37841 7531
rect 37841 7497 37875 7531
rect 37875 7497 37884 7531
rect 37832 7488 37884 7497
rect 38016 7488 38068 7540
rect 18236 7148 18288 7200
rect 20076 7191 20128 7200
rect 20076 7157 20085 7191
rect 20085 7157 20119 7191
rect 20119 7157 20128 7191
rect 20076 7148 20128 7157
rect 24216 7191 24268 7200
rect 24216 7157 24225 7191
rect 24225 7157 24259 7191
rect 24259 7157 24268 7191
rect 24216 7148 24268 7157
rect 24400 7191 24452 7200
rect 24400 7157 24409 7191
rect 24409 7157 24443 7191
rect 24443 7157 24452 7191
rect 24400 7148 24452 7157
rect 29092 7148 29144 7200
rect 29552 7148 29604 7200
rect 31024 7148 31076 7200
rect 31944 7148 31996 7200
rect 34796 7148 34848 7200
rect 35072 7352 35124 7404
rect 35164 7395 35216 7404
rect 35164 7361 35173 7395
rect 35173 7361 35207 7395
rect 35207 7361 35216 7395
rect 35164 7352 35216 7361
rect 38016 7327 38068 7336
rect 38016 7293 38025 7327
rect 38025 7293 38059 7327
rect 38059 7293 38068 7327
rect 38016 7284 38068 7293
rect 37004 7148 37056 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 14464 6944 14516 6996
rect 11980 6808 12032 6860
rect 12256 6783 12308 6792
rect 12256 6749 12265 6783
rect 12265 6749 12299 6783
rect 12299 6749 12308 6783
rect 12256 6740 12308 6749
rect 14740 6876 14792 6928
rect 14740 6783 14792 6792
rect 14188 6672 14240 6724
rect 14740 6749 14749 6783
rect 14749 6749 14783 6783
rect 14783 6749 14792 6783
rect 14740 6740 14792 6749
rect 21732 6944 21784 6996
rect 24032 6944 24084 6996
rect 25136 6987 25188 6996
rect 25136 6953 25145 6987
rect 25145 6953 25179 6987
rect 25179 6953 25188 6987
rect 25136 6944 25188 6953
rect 32956 6987 33008 6996
rect 32956 6953 32965 6987
rect 32965 6953 32999 6987
rect 32999 6953 33008 6987
rect 32956 6944 33008 6953
rect 35440 6944 35492 6996
rect 37832 6944 37884 6996
rect 26056 6876 26108 6928
rect 16212 6808 16264 6860
rect 17960 6851 18012 6860
rect 17960 6817 17969 6851
rect 17969 6817 18003 6851
rect 18003 6817 18012 6851
rect 17960 6808 18012 6817
rect 16028 6783 16080 6792
rect 16028 6749 16037 6783
rect 16037 6749 16071 6783
rect 16071 6749 16080 6783
rect 16028 6740 16080 6749
rect 17408 6783 17460 6792
rect 17408 6749 17417 6783
rect 17417 6749 17451 6783
rect 17451 6749 17460 6783
rect 17408 6740 17460 6749
rect 18420 6808 18472 6860
rect 20444 6808 20496 6860
rect 18328 6740 18380 6792
rect 19984 6783 20036 6792
rect 19984 6749 19993 6783
rect 19993 6749 20027 6783
rect 20027 6749 20036 6783
rect 19984 6740 20036 6749
rect 20076 6740 20128 6792
rect 20536 6783 20588 6792
rect 20536 6749 20545 6783
rect 20545 6749 20579 6783
rect 20579 6749 20588 6783
rect 20536 6740 20588 6749
rect 25780 6808 25832 6860
rect 26148 6808 26200 6860
rect 22468 6783 22520 6792
rect 16580 6672 16632 6724
rect 18052 6672 18104 6724
rect 22468 6749 22477 6783
rect 22477 6749 22511 6783
rect 22511 6749 22520 6783
rect 22468 6740 22520 6749
rect 23204 6740 23256 6792
rect 23296 6672 23348 6724
rect 25412 6715 25464 6724
rect 25412 6681 25421 6715
rect 25421 6681 25455 6715
rect 25455 6681 25464 6715
rect 25412 6672 25464 6681
rect 26240 6783 26292 6792
rect 26240 6749 26249 6783
rect 26249 6749 26283 6783
rect 26283 6749 26292 6783
rect 26240 6740 26292 6749
rect 34152 6876 34204 6928
rect 28356 6808 28408 6860
rect 29736 6808 29788 6860
rect 29276 6740 29328 6792
rect 30104 6783 30156 6792
rect 30104 6749 30113 6783
rect 30113 6749 30147 6783
rect 30147 6749 30156 6783
rect 30656 6808 30708 6860
rect 33048 6808 33100 6860
rect 30104 6740 30156 6749
rect 18696 6604 18748 6656
rect 21364 6604 21416 6656
rect 25964 6604 26016 6656
rect 27436 6672 27488 6724
rect 33968 6740 34020 6792
rect 35072 6740 35124 6792
rect 36728 6851 36780 6860
rect 36728 6817 36737 6851
rect 36737 6817 36771 6851
rect 36771 6817 36780 6851
rect 36728 6808 36780 6817
rect 35532 6783 35584 6792
rect 35532 6749 35541 6783
rect 35541 6749 35575 6783
rect 35575 6749 35584 6783
rect 35532 6740 35584 6749
rect 37004 6783 37056 6792
rect 37004 6749 37038 6783
rect 37038 6749 37056 6783
rect 37004 6740 37056 6749
rect 29184 6604 29236 6656
rect 33324 6604 33376 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 20444 6400 20496 6452
rect 23296 6443 23348 6452
rect 16580 6332 16632 6384
rect 18420 6332 18472 6384
rect 18972 6332 19024 6384
rect 19984 6332 20036 6384
rect 16212 6264 16264 6316
rect 18144 6307 18196 6316
rect 18144 6273 18153 6307
rect 18153 6273 18187 6307
rect 18187 6273 18196 6307
rect 18144 6264 18196 6273
rect 18604 6307 18656 6316
rect 18604 6273 18613 6307
rect 18613 6273 18647 6307
rect 18647 6273 18656 6307
rect 18604 6264 18656 6273
rect 23296 6409 23305 6443
rect 23305 6409 23339 6443
rect 23339 6409 23348 6443
rect 23296 6400 23348 6409
rect 24032 6400 24084 6452
rect 25412 6400 25464 6452
rect 26148 6400 26200 6452
rect 29276 6443 29328 6452
rect 23848 6332 23900 6384
rect 24400 6332 24452 6384
rect 21364 6307 21416 6316
rect 21364 6273 21373 6307
rect 21373 6273 21407 6307
rect 21407 6273 21416 6307
rect 21364 6264 21416 6273
rect 24676 6307 24728 6316
rect 24676 6273 24685 6307
rect 24685 6273 24719 6307
rect 24719 6273 24728 6307
rect 24676 6264 24728 6273
rect 26424 6332 26476 6384
rect 26148 6264 26200 6316
rect 28080 6264 28132 6316
rect 28448 6332 28500 6384
rect 29276 6409 29285 6443
rect 29285 6409 29319 6443
rect 29319 6409 29328 6443
rect 29276 6400 29328 6409
rect 30104 6400 30156 6452
rect 35532 6400 35584 6452
rect 33876 6332 33928 6384
rect 34704 6332 34756 6384
rect 34888 6332 34940 6384
rect 29092 6264 29144 6316
rect 30840 6307 30892 6316
rect 30840 6273 30849 6307
rect 30849 6273 30883 6307
rect 30883 6273 30892 6307
rect 30840 6264 30892 6273
rect 33784 6307 33836 6316
rect 33784 6273 33793 6307
rect 33793 6273 33827 6307
rect 33827 6273 33836 6307
rect 33784 6264 33836 6273
rect 35348 6332 35400 6384
rect 38108 6375 38160 6384
rect 38108 6341 38117 6375
rect 38117 6341 38151 6375
rect 38151 6341 38160 6375
rect 38108 6332 38160 6341
rect 35440 6307 35492 6316
rect 27436 6239 27488 6248
rect 27436 6205 27445 6239
rect 27445 6205 27479 6239
rect 27479 6205 27488 6239
rect 27436 6196 27488 6205
rect 15476 6060 15528 6112
rect 20536 6103 20588 6112
rect 20536 6069 20545 6103
rect 20545 6069 20579 6103
rect 20579 6069 20588 6103
rect 20536 6060 20588 6069
rect 21180 6103 21232 6112
rect 21180 6069 21189 6103
rect 21189 6069 21223 6103
rect 21223 6069 21232 6103
rect 21180 6060 21232 6069
rect 26056 6060 26108 6112
rect 26240 6128 26292 6180
rect 29736 6239 29788 6248
rect 29736 6205 29745 6239
rect 29745 6205 29779 6239
rect 29779 6205 29788 6239
rect 29736 6196 29788 6205
rect 29920 6239 29972 6248
rect 29920 6205 29929 6239
rect 29929 6205 29963 6239
rect 29963 6205 29972 6239
rect 29920 6196 29972 6205
rect 30932 6239 30984 6248
rect 30932 6205 30941 6239
rect 30941 6205 30975 6239
rect 30975 6205 30984 6239
rect 30932 6196 30984 6205
rect 31024 6239 31076 6248
rect 31024 6205 31033 6239
rect 31033 6205 31067 6239
rect 31067 6205 31076 6239
rect 35440 6273 35449 6307
rect 35449 6273 35483 6307
rect 35483 6273 35492 6307
rect 35440 6264 35492 6273
rect 35624 6264 35676 6316
rect 31024 6196 31076 6205
rect 38292 6196 38344 6248
rect 27252 6060 27304 6112
rect 35072 6060 35124 6112
rect 36636 6060 36688 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 17408 5856 17460 5908
rect 25964 5899 26016 5908
rect 25964 5865 25973 5899
rect 25973 5865 26007 5899
rect 26007 5865 26016 5899
rect 25964 5856 26016 5865
rect 28080 5899 28132 5908
rect 28080 5865 28089 5899
rect 28089 5865 28123 5899
rect 28123 5865 28132 5899
rect 28080 5856 28132 5865
rect 35440 5856 35492 5908
rect 38292 5899 38344 5908
rect 38292 5865 38301 5899
rect 38301 5865 38335 5899
rect 38335 5865 38344 5899
rect 38292 5856 38344 5865
rect 22100 5720 22152 5772
rect 23848 5720 23900 5772
rect 24768 5720 24820 5772
rect 25320 5720 25372 5772
rect 26424 5788 26476 5840
rect 27252 5788 27304 5840
rect 26056 5763 26108 5772
rect 15476 5695 15528 5704
rect 15476 5661 15485 5695
rect 15485 5661 15519 5695
rect 15519 5661 15528 5695
rect 15476 5652 15528 5661
rect 16028 5695 16080 5704
rect 16028 5661 16037 5695
rect 16037 5661 16071 5695
rect 16071 5661 16080 5695
rect 16028 5652 16080 5661
rect 18236 5695 18288 5704
rect 18236 5661 18245 5695
rect 18245 5661 18279 5695
rect 18279 5661 18288 5695
rect 18236 5652 18288 5661
rect 18788 5652 18840 5704
rect 21180 5695 21232 5704
rect 21180 5661 21189 5695
rect 21189 5661 21223 5695
rect 21223 5661 21232 5695
rect 21180 5652 21232 5661
rect 26056 5729 26065 5763
rect 26065 5729 26099 5763
rect 26099 5729 26108 5763
rect 26056 5720 26108 5729
rect 27988 5720 28040 5772
rect 28356 5720 28408 5772
rect 33048 5720 33100 5772
rect 36728 5720 36780 5772
rect 28264 5652 28316 5704
rect 28448 5695 28500 5704
rect 28448 5661 28457 5695
rect 28457 5661 28491 5695
rect 28491 5661 28500 5695
rect 28448 5652 28500 5661
rect 31668 5652 31720 5704
rect 30564 5584 30616 5636
rect 33876 5584 33928 5636
rect 35348 5584 35400 5636
rect 37464 5584 37516 5636
rect 18328 5559 18380 5568
rect 18328 5525 18337 5559
rect 18337 5525 18371 5559
rect 18371 5525 18380 5559
rect 18328 5516 18380 5525
rect 24584 5559 24636 5568
rect 24584 5525 24593 5559
rect 24593 5525 24627 5559
rect 24627 5525 24636 5559
rect 24584 5516 24636 5525
rect 24952 5559 25004 5568
rect 24952 5525 24961 5559
rect 24961 5525 24995 5559
rect 24995 5525 25004 5559
rect 24952 5516 25004 5525
rect 30840 5516 30892 5568
rect 33692 5516 33744 5568
rect 35716 5516 35768 5568
rect 37924 5516 37976 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 22836 5312 22888 5364
rect 23480 5312 23532 5364
rect 24676 5312 24728 5364
rect 24952 5312 25004 5364
rect 30564 5312 30616 5364
rect 30840 5355 30892 5364
rect 30840 5321 30849 5355
rect 30849 5321 30883 5355
rect 30883 5321 30892 5355
rect 30840 5312 30892 5321
rect 33784 5312 33836 5364
rect 36636 5355 36688 5364
rect 36636 5321 36645 5355
rect 36645 5321 36679 5355
rect 36679 5321 36688 5355
rect 36636 5312 36688 5321
rect 37464 5355 37516 5364
rect 37464 5321 37473 5355
rect 37473 5321 37507 5355
rect 37507 5321 37516 5355
rect 37464 5312 37516 5321
rect 38292 5312 38344 5364
rect 18328 5244 18380 5296
rect 22100 5176 22152 5228
rect 23204 5244 23256 5296
rect 24584 5244 24636 5296
rect 24768 5244 24820 5296
rect 28356 5244 28408 5296
rect 37924 5287 37976 5296
rect 23020 5176 23072 5228
rect 26240 5219 26292 5228
rect 26240 5185 26249 5219
rect 26249 5185 26283 5219
rect 26283 5185 26292 5219
rect 26240 5176 26292 5185
rect 26976 5176 27028 5228
rect 31760 5176 31812 5228
rect 32588 5219 32640 5228
rect 32588 5185 32622 5219
rect 32622 5185 32640 5219
rect 32588 5176 32640 5185
rect 37924 5253 37933 5287
rect 37933 5253 37967 5287
rect 37967 5253 37976 5287
rect 37924 5244 37976 5253
rect 35532 5219 35584 5228
rect 35532 5185 35566 5219
rect 35566 5185 35584 5219
rect 35532 5176 35584 5185
rect 18972 5108 19024 5160
rect 23204 5108 23256 5160
rect 24032 5151 24084 5160
rect 24032 5117 24041 5151
rect 24041 5117 24075 5151
rect 24075 5117 24084 5151
rect 24032 5108 24084 5117
rect 26516 5151 26568 5160
rect 26516 5117 26525 5151
rect 26525 5117 26559 5151
rect 26559 5117 26568 5151
rect 26516 5108 26568 5117
rect 30748 5108 30800 5160
rect 32220 5108 32272 5160
rect 33600 5108 33652 5160
rect 38016 5151 38068 5160
rect 38016 5117 38025 5151
rect 38025 5117 38059 5151
rect 38059 5117 38068 5151
rect 38016 5108 38068 5117
rect 17960 5040 18012 5092
rect 18512 5015 18564 5024
rect 18512 4981 18521 5015
rect 18521 4981 18555 5015
rect 18555 4981 18564 5015
rect 18512 4972 18564 4981
rect 25872 5015 25924 5024
rect 25872 4981 25881 5015
rect 25881 4981 25915 5015
rect 25915 4981 25924 5015
rect 25872 4972 25924 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 23020 4811 23072 4820
rect 23020 4777 23029 4811
rect 23029 4777 23063 4811
rect 23063 4777 23072 4811
rect 23020 4768 23072 4777
rect 26976 4811 27028 4820
rect 26976 4777 26985 4811
rect 26985 4777 27019 4811
rect 27019 4777 27028 4811
rect 26976 4768 27028 4777
rect 29000 4768 29052 4820
rect 29736 4768 29788 4820
rect 30932 4768 30984 4820
rect 32588 4811 32640 4820
rect 32588 4777 32597 4811
rect 32597 4777 32631 4811
rect 32631 4777 32640 4811
rect 32588 4768 32640 4777
rect 35532 4768 35584 4820
rect 23664 4700 23716 4752
rect 32220 4700 32272 4752
rect 17408 4632 17460 4684
rect 23572 4675 23624 4684
rect 23572 4641 23581 4675
rect 23581 4641 23615 4675
rect 23615 4641 23624 4675
rect 23572 4632 23624 4641
rect 15936 4607 15988 4616
rect 15936 4573 15945 4607
rect 15945 4573 15979 4607
rect 15979 4573 15988 4607
rect 15936 4564 15988 4573
rect 23480 4564 23532 4616
rect 24032 4564 24084 4616
rect 27436 4607 27488 4616
rect 27436 4573 27445 4607
rect 27445 4573 27479 4607
rect 27479 4573 27488 4607
rect 27436 4564 27488 4573
rect 30288 4564 30340 4616
rect 33048 4632 33100 4684
rect 35900 4632 35952 4684
rect 38016 4700 38068 4752
rect 38108 4675 38160 4684
rect 38108 4641 38117 4675
rect 38117 4641 38151 4675
rect 38151 4641 38160 4675
rect 38108 4632 38160 4641
rect 33784 4564 33836 4616
rect 36636 4564 36688 4616
rect 25872 4539 25924 4548
rect 25872 4505 25906 4539
rect 25906 4505 25924 4539
rect 25872 4496 25924 4505
rect 27896 4496 27948 4548
rect 30012 4539 30064 4548
rect 30012 4505 30046 4539
rect 30046 4505 30064 4539
rect 30012 4496 30064 4505
rect 23848 4428 23900 4480
rect 28172 4428 28224 4480
rect 35900 4428 35952 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 27896 4267 27948 4276
rect 27896 4233 27905 4267
rect 27905 4233 27939 4267
rect 27939 4233 27948 4267
rect 27896 4224 27948 4233
rect 29000 4224 29052 4276
rect 30012 4224 30064 4276
rect 30932 4224 30984 4276
rect 30472 4156 30524 4208
rect 15936 4088 15988 4140
rect 18512 4088 18564 4140
rect 28356 4131 28408 4140
rect 28356 4097 28365 4131
rect 28365 4097 28399 4131
rect 28399 4097 28408 4131
rect 28356 4088 28408 4097
rect 33600 4131 33652 4140
rect 19432 4020 19484 4072
rect 23572 4020 23624 4072
rect 33600 4097 33609 4131
rect 33609 4097 33643 4131
rect 33643 4097 33652 4131
rect 33600 4088 33652 4097
rect 33692 4088 33744 4140
rect 38108 4131 38160 4140
rect 29552 4020 29604 4072
rect 30288 4020 30340 4072
rect 38108 4097 38117 4131
rect 38117 4097 38151 4131
rect 38151 4097 38160 4131
rect 38108 4088 38160 4097
rect 29368 3884 29420 3936
rect 35348 3884 35400 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 27712 3000 27764 3052
rect 38108 2975 38160 2984
rect 38108 2941 38117 2975
rect 38117 2941 38151 2975
rect 38151 2941 38160 2975
rect 38108 2932 38160 2941
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 27344 2388 27396 2440
rect 38108 2363 38160 2372
rect 38108 2329 38117 2363
rect 38117 2329 38151 2363
rect 38151 2329 38160 2363
rect 38108 2320 38160 2329
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 1766 39200 1822 40000
rect 5078 39200 5134 40000
rect 8390 39200 8446 40000
rect 11702 39200 11758 40000
rect 15014 39200 15070 40000
rect 18326 39200 18382 40000
rect 21638 39200 21694 40000
rect 21744 39222 22048 39250
rect 1780 37262 1808 39200
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 5092 37262 5120 39200
rect 8404 37262 8432 39200
rect 9404 37324 9456 37330
rect 9404 37266 9456 37272
rect 1768 37256 1820 37262
rect 1768 37198 1820 37204
rect 5080 37256 5132 37262
rect 5080 37198 5132 37204
rect 8392 37256 8444 37262
rect 8392 37198 8444 37204
rect 5540 37188 5592 37194
rect 5540 37130 5592 37136
rect 5724 37188 5776 37194
rect 5724 37130 5776 37136
rect 9312 37188 9364 37194
rect 9312 37130 9364 37136
rect 5552 36786 5580 37130
rect 4528 36780 4580 36786
rect 5540 36780 5592 36786
rect 4580 36740 4660 36768
rect 4528 36722 4580 36728
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4632 36174 4660 36740
rect 5540 36722 5592 36728
rect 4620 36168 4672 36174
rect 4620 36110 4672 36116
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4632 34746 4660 36110
rect 5552 36106 5580 36722
rect 5632 36644 5684 36650
rect 5632 36586 5684 36592
rect 5644 36242 5672 36586
rect 5632 36236 5684 36242
rect 5632 36178 5684 36184
rect 5540 36100 5592 36106
rect 5540 36042 5592 36048
rect 5264 36032 5316 36038
rect 5264 35974 5316 35980
rect 5080 34944 5132 34950
rect 5080 34886 5132 34892
rect 4620 34740 4672 34746
rect 4620 34682 4672 34688
rect 5092 34610 5120 34886
rect 5080 34604 5132 34610
rect 5080 34546 5132 34552
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 5172 33516 5224 33522
rect 5172 33458 5224 33464
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4620 32972 4672 32978
rect 4620 32914 4672 32920
rect 4528 32904 4580 32910
rect 4528 32846 4580 32852
rect 4540 32366 4568 32846
rect 4632 32434 4660 32914
rect 5184 32910 5212 33458
rect 5276 32910 5304 35974
rect 5736 35018 5764 37130
rect 9128 37120 9180 37126
rect 9128 37062 9180 37068
rect 9140 36854 9168 37062
rect 9128 36848 9180 36854
rect 9128 36790 9180 36796
rect 7656 36712 7708 36718
rect 7656 36654 7708 36660
rect 7932 36712 7984 36718
rect 7932 36654 7984 36660
rect 5908 36236 5960 36242
rect 5908 36178 5960 36184
rect 5724 35012 5776 35018
rect 5724 34954 5776 34960
rect 5540 34944 5592 34950
rect 5540 34886 5592 34892
rect 5552 34746 5580 34886
rect 5540 34740 5592 34746
rect 5540 34682 5592 34688
rect 5552 34066 5580 34682
rect 5540 34060 5592 34066
rect 5540 34002 5592 34008
rect 5736 33998 5764 34954
rect 5920 34474 5948 36178
rect 7104 36100 7156 36106
rect 7104 36042 7156 36048
rect 7116 35834 7144 36042
rect 7104 35828 7156 35834
rect 7104 35770 7156 35776
rect 7668 35630 7696 36654
rect 7944 36174 7972 36654
rect 9324 36310 9352 37130
rect 8576 36304 8628 36310
rect 8576 36246 8628 36252
rect 9312 36304 9364 36310
rect 9312 36246 9364 36252
rect 7932 36168 7984 36174
rect 7932 36110 7984 36116
rect 7840 36100 7892 36106
rect 7840 36042 7892 36048
rect 7748 36032 7800 36038
rect 7748 35974 7800 35980
rect 7760 35834 7788 35974
rect 7748 35828 7800 35834
rect 7748 35770 7800 35776
rect 7656 35624 7708 35630
rect 7656 35566 7708 35572
rect 7668 35154 7696 35566
rect 7656 35148 7708 35154
rect 7656 35090 7708 35096
rect 7012 34740 7064 34746
rect 7012 34682 7064 34688
rect 5908 34468 5960 34474
rect 5908 34410 5960 34416
rect 5920 34066 5948 34410
rect 5908 34060 5960 34066
rect 5908 34002 5960 34008
rect 5724 33992 5776 33998
rect 5722 33960 5724 33969
rect 5776 33960 5778 33969
rect 5722 33895 5778 33904
rect 5356 33856 5408 33862
rect 5356 33798 5408 33804
rect 5368 32978 5396 33798
rect 7024 33522 7052 34682
rect 7760 34610 7788 35770
rect 7852 34610 7880 36042
rect 8300 35760 8352 35766
rect 8300 35702 8352 35708
rect 8312 34678 8340 35702
rect 8300 34672 8352 34678
rect 8300 34614 8352 34620
rect 7748 34604 7800 34610
rect 7748 34546 7800 34552
rect 7840 34604 7892 34610
rect 7840 34546 7892 34552
rect 7748 34468 7800 34474
rect 7748 34410 7800 34416
rect 7760 33998 7788 34410
rect 8208 34060 8260 34066
rect 8208 34002 8260 34008
rect 7748 33992 7800 33998
rect 7748 33934 7800 33940
rect 7380 33584 7432 33590
rect 7380 33526 7432 33532
rect 6552 33516 6604 33522
rect 6552 33458 6604 33464
rect 7012 33516 7064 33522
rect 7064 33476 7144 33504
rect 7012 33458 7064 33464
rect 5356 32972 5408 32978
rect 5356 32914 5408 32920
rect 5816 32972 5868 32978
rect 5816 32914 5868 32920
rect 5172 32904 5224 32910
rect 5172 32846 5224 32852
rect 5264 32904 5316 32910
rect 5264 32846 5316 32852
rect 4712 32836 4764 32842
rect 4712 32778 4764 32784
rect 5724 32836 5776 32842
rect 5724 32778 5776 32784
rect 4724 32502 4752 32778
rect 4712 32496 4764 32502
rect 4712 32438 4764 32444
rect 4620 32428 4672 32434
rect 4620 32370 4672 32376
rect 4528 32360 4580 32366
rect 4528 32302 4580 32308
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4724 31890 4752 32438
rect 5736 32434 5764 32778
rect 5724 32428 5776 32434
rect 5724 32370 5776 32376
rect 5448 32292 5500 32298
rect 5448 32234 5500 32240
rect 4896 31952 4948 31958
rect 4896 31894 4948 31900
rect 4712 31884 4764 31890
rect 4712 31826 4764 31832
rect 4908 31754 4936 31894
rect 5170 31784 5226 31793
rect 4908 31726 5028 31754
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4896 30660 4948 30666
rect 4896 30602 4948 30608
rect 4908 30394 4936 30602
rect 4896 30388 4948 30394
rect 4896 30330 4948 30336
rect 2780 30252 2832 30258
rect 2780 30194 2832 30200
rect 3976 30252 4028 30258
rect 3976 30194 4028 30200
rect 2792 26994 2820 30194
rect 3988 29850 4016 30194
rect 4620 30048 4672 30054
rect 4620 29990 4672 29996
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 3976 29844 4028 29850
rect 3976 29786 4028 29792
rect 4160 29708 4212 29714
rect 4160 29650 4212 29656
rect 3332 29504 3384 29510
rect 3332 29446 3384 29452
rect 3344 29238 3372 29446
rect 3332 29232 3384 29238
rect 3332 29174 3384 29180
rect 4068 29164 4120 29170
rect 4068 29106 4120 29112
rect 3976 28960 4028 28966
rect 3976 28902 4028 28908
rect 3988 27674 4016 28902
rect 4080 28529 4108 29106
rect 4172 28966 4200 29650
rect 4632 29646 4660 29990
rect 4620 29640 4672 29646
rect 4620 29582 4672 29588
rect 4804 29232 4856 29238
rect 4804 29174 4856 29180
rect 4620 29028 4672 29034
rect 4620 28970 4672 28976
rect 4160 28960 4212 28966
rect 4160 28902 4212 28908
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4066 28520 4122 28529
rect 4066 28455 4122 28464
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3976 27668 4028 27674
rect 3976 27610 4028 27616
rect 4436 27668 4488 27674
rect 4488 27628 4568 27656
rect 4436 27610 4488 27616
rect 4436 27464 4488 27470
rect 4540 27452 4568 27628
rect 4632 27606 4660 28970
rect 4712 28960 4764 28966
rect 4712 28902 4764 28908
rect 4724 28558 4752 28902
rect 4816 28762 4844 29174
rect 4896 29164 4948 29170
rect 4896 29106 4948 29112
rect 4908 29034 4936 29106
rect 4896 29028 4948 29034
rect 4896 28970 4948 28976
rect 4804 28756 4856 28762
rect 4804 28698 4856 28704
rect 4712 28552 4764 28558
rect 4712 28494 4764 28500
rect 4620 27600 4672 27606
rect 4620 27542 4672 27548
rect 4724 27538 4752 28494
rect 4804 28076 4856 28082
rect 4804 28018 4856 28024
rect 4816 27674 4844 28018
rect 4804 27668 4856 27674
rect 4804 27610 4856 27616
rect 4712 27532 4764 27538
rect 4712 27474 4764 27480
rect 4620 27464 4672 27470
rect 4540 27424 4620 27452
rect 4436 27406 4488 27412
rect 4816 27418 4844 27610
rect 4620 27406 4672 27412
rect 3976 27328 4028 27334
rect 3976 27270 4028 27276
rect 3988 27062 4016 27270
rect 4448 27130 4476 27406
rect 4528 27328 4580 27334
rect 4528 27270 4580 27276
rect 4436 27124 4488 27130
rect 4436 27066 4488 27072
rect 4540 27062 4568 27270
rect 3976 27056 4028 27062
rect 3976 26998 4028 27004
rect 4528 27056 4580 27062
rect 4528 26998 4580 27004
rect 2780 26988 2832 26994
rect 2780 26930 2832 26936
rect 2792 24818 2820 26930
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4528 26580 4580 26586
rect 4528 26522 4580 26528
rect 4436 26512 4488 26518
rect 4436 26454 4488 26460
rect 4448 25770 4476 26454
rect 4540 25786 4568 26522
rect 4632 25888 4660 27406
rect 4724 27390 4844 27418
rect 4724 26246 4752 27390
rect 4802 27160 4858 27169
rect 4802 27095 4858 27104
rect 4816 26586 4844 27095
rect 4804 26580 4856 26586
rect 4804 26522 4856 26528
rect 4804 26444 4856 26450
rect 4804 26386 4856 26392
rect 4712 26240 4764 26246
rect 4712 26182 4764 26188
rect 4632 25860 4752 25888
rect 4436 25764 4488 25770
rect 4540 25758 4660 25786
rect 4436 25706 4488 25712
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4160 25288 4212 25294
rect 4160 25230 4212 25236
rect 4436 25288 4488 25294
rect 4436 25230 4488 25236
rect 3976 25152 4028 25158
rect 3976 25094 4028 25100
rect 3988 24886 4016 25094
rect 4172 24954 4200 25230
rect 4160 24948 4212 24954
rect 4160 24890 4212 24896
rect 3976 24880 4028 24886
rect 3976 24822 4028 24828
rect 2780 24812 2832 24818
rect 2780 24754 2832 24760
rect 4448 24614 4476 25230
rect 4436 24608 4488 24614
rect 4436 24550 4488 24556
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4160 24132 4212 24138
rect 4160 24074 4212 24080
rect 4172 23866 4200 24074
rect 4160 23860 4212 23866
rect 4160 23802 4212 23808
rect 2780 23724 2832 23730
rect 2780 23666 2832 23672
rect 3976 23724 4028 23730
rect 3976 23666 4028 23672
rect 2792 21554 2820 23666
rect 3988 23322 4016 23666
rect 4172 23508 4200 23802
rect 4632 23798 4660 25758
rect 4724 25362 4752 25860
rect 4712 25356 4764 25362
rect 4712 25298 4764 25304
rect 4724 24052 4752 25298
rect 4816 24818 4844 26386
rect 4908 25838 4936 28970
rect 5000 27962 5028 31726
rect 5170 31719 5226 31728
rect 5184 29866 5212 31719
rect 5460 31346 5488 32234
rect 5736 32212 5764 32370
rect 5552 32184 5764 32212
rect 5552 31890 5580 32184
rect 5540 31884 5592 31890
rect 5540 31826 5592 31832
rect 5552 31346 5580 31826
rect 5828 31822 5856 32914
rect 6460 32360 6512 32366
rect 6460 32302 6512 32308
rect 6472 32026 6500 32302
rect 6564 32026 6592 33458
rect 6828 33312 6880 33318
rect 6828 33254 6880 33260
rect 6736 32292 6788 32298
rect 6736 32234 6788 32240
rect 6644 32224 6696 32230
rect 6644 32166 6696 32172
rect 6460 32020 6512 32026
rect 6460 31962 6512 31968
rect 6552 32020 6604 32026
rect 6552 31962 6604 31968
rect 5632 31816 5684 31822
rect 5632 31758 5684 31764
rect 5816 31816 5868 31822
rect 5816 31758 5868 31764
rect 5448 31340 5500 31346
rect 5448 31282 5500 31288
rect 5540 31340 5592 31346
rect 5540 31282 5592 31288
rect 5264 30660 5316 30666
rect 5264 30602 5316 30608
rect 5092 29838 5212 29866
rect 5092 29714 5120 29838
rect 5276 29782 5304 30602
rect 5460 30122 5488 31282
rect 5540 31136 5592 31142
rect 5540 31078 5592 31084
rect 5552 30258 5580 31078
rect 5540 30252 5592 30258
rect 5540 30194 5592 30200
rect 5448 30116 5500 30122
rect 5448 30058 5500 30064
rect 5264 29776 5316 29782
rect 5184 29724 5264 29730
rect 5184 29718 5316 29724
rect 5080 29708 5132 29714
rect 5080 29650 5132 29656
rect 5184 29702 5304 29718
rect 5184 29306 5212 29702
rect 5356 29640 5408 29646
rect 5356 29582 5408 29588
rect 5448 29640 5500 29646
rect 5448 29582 5500 29588
rect 5264 29572 5316 29578
rect 5264 29514 5316 29520
rect 5172 29300 5224 29306
rect 5172 29242 5224 29248
rect 5276 29170 5304 29514
rect 5264 29164 5316 29170
rect 5264 29106 5316 29112
rect 5276 28014 5304 29106
rect 5368 29102 5396 29582
rect 5460 29238 5488 29582
rect 5448 29232 5500 29238
rect 5448 29174 5500 29180
rect 5356 29096 5408 29102
rect 5356 29038 5408 29044
rect 5368 28558 5396 29038
rect 5552 28694 5580 30194
rect 5644 29714 5672 31758
rect 6656 31686 6684 32166
rect 6748 31822 6776 32234
rect 6840 31958 6868 33254
rect 6920 32428 6972 32434
rect 6920 32370 6972 32376
rect 6828 31952 6880 31958
rect 6828 31894 6880 31900
rect 6736 31816 6788 31822
rect 6736 31758 6788 31764
rect 6644 31680 6696 31686
rect 6472 31640 6644 31668
rect 6092 31136 6144 31142
rect 6092 31078 6144 31084
rect 6104 30666 6132 31078
rect 6092 30660 6144 30666
rect 6092 30602 6144 30608
rect 5632 29708 5684 29714
rect 5632 29650 5684 29656
rect 6000 29708 6052 29714
rect 6000 29650 6052 29656
rect 5540 28688 5592 28694
rect 5540 28630 5592 28636
rect 5356 28552 5408 28558
rect 5356 28494 5408 28500
rect 5446 28520 5502 28529
rect 5446 28455 5448 28464
rect 5500 28455 5502 28464
rect 5814 28520 5870 28529
rect 5814 28455 5870 28464
rect 5448 28426 5500 28432
rect 5724 28416 5776 28422
rect 5724 28358 5776 28364
rect 5264 28008 5316 28014
rect 5000 27934 5212 27962
rect 5264 27950 5316 27956
rect 4988 27872 5040 27878
rect 4988 27814 5040 27820
rect 5080 27872 5132 27878
rect 5080 27814 5132 27820
rect 5000 27282 5028 27814
rect 5092 27470 5120 27814
rect 5080 27464 5132 27470
rect 5080 27406 5132 27412
rect 5000 27254 5120 27282
rect 4988 26852 5040 26858
rect 4988 26794 5040 26800
rect 4896 25832 4948 25838
rect 4896 25774 4948 25780
rect 4896 25696 4948 25702
rect 4896 25638 4948 25644
rect 4908 25362 4936 25638
rect 4896 25356 4948 25362
rect 4896 25298 4948 25304
rect 4804 24812 4856 24818
rect 4804 24754 4856 24760
rect 4804 24064 4856 24070
rect 4724 24024 4804 24052
rect 4804 24006 4856 24012
rect 4620 23792 4672 23798
rect 4620 23734 4672 23740
rect 4712 23724 4764 23730
rect 4712 23666 4764 23672
rect 4080 23480 4200 23508
rect 4620 23520 4672 23526
rect 3976 23316 4028 23322
rect 3976 23258 4028 23264
rect 4080 23202 4108 23480
rect 4620 23462 4672 23468
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4080 23174 4200 23202
rect 4172 23118 4200 23174
rect 4632 23118 4660 23462
rect 4160 23112 4212 23118
rect 4160 23054 4212 23060
rect 4620 23112 4672 23118
rect 4620 23054 4672 23060
rect 4724 22778 4752 23666
rect 4816 23186 4844 24006
rect 4804 23180 4856 23186
rect 4804 23122 4856 23128
rect 4896 23112 4948 23118
rect 4896 23054 4948 23060
rect 4712 22772 4764 22778
rect 4712 22714 4764 22720
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4620 22092 4672 22098
rect 4620 22034 4672 22040
rect 3976 21888 4028 21894
rect 3976 21830 4028 21836
rect 4344 21888 4396 21894
rect 4344 21830 4396 21836
rect 3988 21622 4016 21830
rect 3976 21616 4028 21622
rect 3976 21558 4028 21564
rect 2780 21548 2832 21554
rect 2780 21490 2832 21496
rect 2792 21010 2820 21490
rect 4356 21418 4384 21830
rect 4632 21486 4660 22034
rect 4724 22030 4752 22714
rect 4908 22642 4936 23054
rect 4896 22636 4948 22642
rect 4896 22578 4948 22584
rect 4712 22024 4764 22030
rect 4712 21966 4764 21972
rect 4620 21480 4672 21486
rect 4620 21422 4672 21428
rect 4344 21412 4396 21418
rect 4344 21354 4396 21360
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 2780 21004 2832 21010
rect 2780 20946 2832 20952
rect 3976 21004 4028 21010
rect 3976 20946 4028 20952
rect 3988 20330 4016 20946
rect 4632 20398 4660 21422
rect 5000 20602 5028 26794
rect 5092 26466 5120 27254
rect 5184 27169 5212 27934
rect 5632 27600 5684 27606
rect 5632 27542 5684 27548
rect 5264 27464 5316 27470
rect 5264 27406 5316 27412
rect 5448 27464 5500 27470
rect 5448 27406 5500 27412
rect 5170 27160 5226 27169
rect 5170 27095 5226 27104
rect 5172 27056 5224 27062
rect 5172 26998 5224 27004
rect 5184 26586 5212 26998
rect 5172 26580 5224 26586
rect 5172 26522 5224 26528
rect 5276 26518 5304 27406
rect 5356 26920 5408 26926
rect 5356 26862 5408 26868
rect 5264 26512 5316 26518
rect 5092 26438 5212 26466
rect 5264 26454 5316 26460
rect 5184 26382 5212 26438
rect 5172 26376 5224 26382
rect 5224 26324 5304 26330
rect 5172 26318 5304 26324
rect 5184 26302 5304 26318
rect 5276 26246 5304 26302
rect 5172 26240 5224 26246
rect 5172 26182 5224 26188
rect 5264 26240 5316 26246
rect 5264 26182 5316 26188
rect 5080 26036 5132 26042
rect 5080 25978 5132 25984
rect 5092 24886 5120 25978
rect 5184 25702 5212 26182
rect 5172 25696 5224 25702
rect 5172 25638 5224 25644
rect 5184 25430 5212 25638
rect 5172 25424 5224 25430
rect 5172 25366 5224 25372
rect 5080 24880 5132 24886
rect 5080 24822 5132 24828
rect 5184 24698 5212 25366
rect 5368 25294 5396 26862
rect 5460 25362 5488 27406
rect 5540 26784 5592 26790
rect 5540 26726 5592 26732
rect 5552 26586 5580 26726
rect 5540 26580 5592 26586
rect 5540 26522 5592 26528
rect 5540 26376 5592 26382
rect 5540 26318 5592 26324
rect 5448 25356 5500 25362
rect 5448 25298 5500 25304
rect 5356 25288 5408 25294
rect 5356 25230 5408 25236
rect 5092 24670 5212 24698
rect 5092 22710 5120 24670
rect 5172 24608 5224 24614
rect 5172 24550 5224 24556
rect 5184 23798 5212 24550
rect 5172 23792 5224 23798
rect 5172 23734 5224 23740
rect 5368 23526 5396 25230
rect 5460 24954 5488 25298
rect 5552 25158 5580 26318
rect 5644 25498 5672 27542
rect 5736 27402 5764 28358
rect 5724 27396 5776 27402
rect 5724 27338 5776 27344
rect 5736 26994 5764 27338
rect 5724 26988 5776 26994
rect 5724 26930 5776 26936
rect 5632 25492 5684 25498
rect 5632 25434 5684 25440
rect 5540 25152 5592 25158
rect 5540 25094 5592 25100
rect 5448 24948 5500 24954
rect 5448 24890 5500 24896
rect 5552 23866 5580 25094
rect 5644 24818 5672 25434
rect 5632 24812 5684 24818
rect 5632 24754 5684 24760
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 5828 23730 5856 28455
rect 6012 26489 6040 29650
rect 6104 27470 6132 30602
rect 6368 30252 6420 30258
rect 6368 30194 6420 30200
rect 6276 30184 6328 30190
rect 6276 30126 6328 30132
rect 6288 29782 6316 30126
rect 6380 29850 6408 30194
rect 6368 29844 6420 29850
rect 6368 29786 6420 29792
rect 6276 29776 6328 29782
rect 6328 29724 6408 29730
rect 6276 29718 6408 29724
rect 6288 29702 6408 29718
rect 6288 29653 6316 29702
rect 6380 29578 6408 29702
rect 6368 29572 6420 29578
rect 6368 29514 6420 29520
rect 6184 29504 6236 29510
rect 6184 29446 6236 29452
rect 6196 28762 6224 29446
rect 6184 28756 6236 28762
rect 6184 28698 6236 28704
rect 6472 28490 6500 31640
rect 6644 31622 6696 31628
rect 6644 31340 6696 31346
rect 6644 31282 6696 31288
rect 6552 30932 6604 30938
rect 6552 30874 6604 30880
rect 6564 30394 6592 30874
rect 6656 30802 6684 31282
rect 6644 30796 6696 30802
rect 6644 30738 6696 30744
rect 6552 30388 6604 30394
rect 6552 30330 6604 30336
rect 6552 30184 6604 30190
rect 6552 30126 6604 30132
rect 6564 29782 6592 30126
rect 6552 29776 6604 29782
rect 6552 29718 6604 29724
rect 6656 29646 6684 30738
rect 6840 30410 6868 31894
rect 6932 30870 6960 32370
rect 7012 31816 7064 31822
rect 7012 31758 7064 31764
rect 7024 30938 7052 31758
rect 7012 30932 7064 30938
rect 7012 30874 7064 30880
rect 6920 30864 6972 30870
rect 6920 30806 6972 30812
rect 6748 30382 6868 30410
rect 6748 29714 6776 30382
rect 6840 30258 6960 30274
rect 6840 30252 6972 30258
rect 6840 30246 6920 30252
rect 6736 29708 6788 29714
rect 6736 29650 6788 29656
rect 6644 29640 6696 29646
rect 6644 29582 6696 29588
rect 6748 28966 6776 29650
rect 6840 29510 6868 30246
rect 6920 30194 6972 30200
rect 7116 30190 7144 33476
rect 7392 32910 7420 33526
rect 7472 33448 7524 33454
rect 7472 33390 7524 33396
rect 7380 32904 7432 32910
rect 7380 32846 7432 32852
rect 7484 32842 7512 33390
rect 7760 32910 7788 33934
rect 8116 33516 8168 33522
rect 8116 33458 8168 33464
rect 8128 33046 8156 33458
rect 8116 33040 8168 33046
rect 8116 32982 8168 32988
rect 7748 32904 7800 32910
rect 7748 32846 7800 32852
rect 7472 32836 7524 32842
rect 7472 32778 7524 32784
rect 7380 30864 7432 30870
rect 7380 30806 7432 30812
rect 7196 30796 7248 30802
rect 7196 30738 7248 30744
rect 7104 30184 7156 30190
rect 7104 30126 7156 30132
rect 7012 29640 7064 29646
rect 7012 29582 7064 29588
rect 7104 29640 7156 29646
rect 7104 29582 7156 29588
rect 6828 29504 6880 29510
rect 6828 29446 6880 29452
rect 7024 29238 7052 29582
rect 7012 29232 7064 29238
rect 7012 29174 7064 29180
rect 7116 29034 7144 29582
rect 7104 29028 7156 29034
rect 7104 28970 7156 28976
rect 6736 28960 6788 28966
rect 6736 28902 6788 28908
rect 6748 28490 6776 28902
rect 6920 28552 6972 28558
rect 6920 28494 6972 28500
rect 6460 28484 6512 28490
rect 6460 28426 6512 28432
rect 6736 28484 6788 28490
rect 6736 28426 6788 28432
rect 6368 28008 6420 28014
rect 6368 27950 6420 27956
rect 6092 27464 6144 27470
rect 6092 27406 6144 27412
rect 6276 26512 6328 26518
rect 5998 26480 6054 26489
rect 6276 26454 6328 26460
rect 5998 26415 6054 26424
rect 5816 23724 5868 23730
rect 5816 23666 5868 23672
rect 5356 23520 5408 23526
rect 5356 23462 5408 23468
rect 5080 22704 5132 22710
rect 5080 22646 5132 22652
rect 5828 21554 5856 23666
rect 5908 23520 5960 23526
rect 5908 23462 5960 23468
rect 5920 23322 5948 23462
rect 5908 23316 5960 23322
rect 5908 23258 5960 23264
rect 6012 23186 6040 26415
rect 6288 26382 6316 26454
rect 6276 26376 6328 26382
rect 6276 26318 6328 26324
rect 6380 25974 6408 27950
rect 6472 26994 6500 28426
rect 6748 27878 6776 28426
rect 6736 27872 6788 27878
rect 6736 27814 6788 27820
rect 6932 27606 6960 28494
rect 7012 28484 7064 28490
rect 7012 28426 7064 28432
rect 6920 27600 6972 27606
rect 6920 27542 6972 27548
rect 6460 26988 6512 26994
rect 6460 26930 6512 26936
rect 6828 26920 6880 26926
rect 6828 26862 6880 26868
rect 6840 26790 6868 26862
rect 6828 26784 6880 26790
rect 6828 26726 6880 26732
rect 6840 26466 6868 26726
rect 6748 26438 6868 26466
rect 6748 26382 6776 26438
rect 6736 26376 6788 26382
rect 6736 26318 6788 26324
rect 6368 25968 6420 25974
rect 6368 25910 6420 25916
rect 6736 25900 6788 25906
rect 6736 25842 6788 25848
rect 6460 25696 6512 25702
rect 6460 25638 6512 25644
rect 6472 25362 6500 25638
rect 6460 25356 6512 25362
rect 6460 25298 6512 25304
rect 6748 24818 6776 25842
rect 6932 25514 6960 27542
rect 7024 27470 7052 28426
rect 7116 28218 7144 28970
rect 7104 28212 7156 28218
rect 7104 28154 7156 28160
rect 7104 27940 7156 27946
rect 7104 27882 7156 27888
rect 7012 27464 7064 27470
rect 7012 27406 7064 27412
rect 7024 26450 7052 27406
rect 7012 26444 7064 26450
rect 7012 26386 7064 26392
rect 6932 25486 7052 25514
rect 6920 25356 6972 25362
rect 6920 25298 6972 25304
rect 6932 24818 6960 25298
rect 6736 24812 6788 24818
rect 6736 24754 6788 24760
rect 6920 24812 6972 24818
rect 6920 24754 6972 24760
rect 6644 24744 6696 24750
rect 6644 24686 6696 24692
rect 6656 24154 6684 24686
rect 6656 24138 6868 24154
rect 6656 24132 6880 24138
rect 6656 24126 6828 24132
rect 6828 24074 6880 24080
rect 7024 23798 7052 25486
rect 7012 23792 7064 23798
rect 7012 23734 7064 23740
rect 7116 23730 7144 27882
rect 7208 26382 7236 30738
rect 7288 29504 7340 29510
rect 7288 29446 7340 29452
rect 7196 26376 7248 26382
rect 7196 26318 7248 26324
rect 7208 24818 7236 26318
rect 7196 24812 7248 24818
rect 7196 24754 7248 24760
rect 7208 24342 7236 24754
rect 7196 24336 7248 24342
rect 7196 24278 7248 24284
rect 7196 23792 7248 23798
rect 7196 23734 7248 23740
rect 6828 23724 6880 23730
rect 6828 23666 6880 23672
rect 7104 23724 7156 23730
rect 7104 23666 7156 23672
rect 6644 23656 6696 23662
rect 6644 23598 6696 23604
rect 6000 23180 6052 23186
rect 6000 23122 6052 23128
rect 6656 23118 6684 23598
rect 6644 23112 6696 23118
rect 6644 23054 6696 23060
rect 6736 23112 6788 23118
rect 6840 23100 6868 23666
rect 7116 23610 7144 23666
rect 7024 23582 7144 23610
rect 6920 23520 6972 23526
rect 6920 23462 6972 23468
rect 6932 23254 6960 23462
rect 6920 23248 6972 23254
rect 6920 23190 6972 23196
rect 6920 23112 6972 23118
rect 6840 23072 6920 23100
rect 6736 23054 6788 23060
rect 6920 23054 6972 23060
rect 6656 22778 6684 23054
rect 6644 22772 6696 22778
rect 6644 22714 6696 22720
rect 5908 22500 5960 22506
rect 5908 22442 5960 22448
rect 5920 21690 5948 22442
rect 6748 21962 6776 23054
rect 6736 21956 6788 21962
rect 6736 21898 6788 21904
rect 6644 21888 6696 21894
rect 6644 21830 6696 21836
rect 5908 21684 5960 21690
rect 5908 21626 5960 21632
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 5920 21146 5948 21626
rect 6656 21622 6684 21830
rect 6644 21616 6696 21622
rect 6644 21558 6696 21564
rect 6736 21548 6788 21554
rect 6736 21490 6788 21496
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 6000 21344 6052 21350
rect 6000 21286 6052 21292
rect 5908 21140 5960 21146
rect 5908 21082 5960 21088
rect 6012 20942 6040 21286
rect 6000 20936 6052 20942
rect 6000 20878 6052 20884
rect 6552 20800 6604 20806
rect 6552 20742 6604 20748
rect 4988 20596 5040 20602
rect 4988 20538 5040 20544
rect 5356 20460 5408 20466
rect 5356 20402 5408 20408
rect 4620 20392 4672 20398
rect 4620 20334 4672 20340
rect 3976 20324 4028 20330
rect 3976 20266 4028 20272
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 3896 19854 3924 20198
rect 3988 19922 4016 20266
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3976 19916 4028 19922
rect 3976 19858 4028 19864
rect 3884 19848 3936 19854
rect 3884 19790 3936 19796
rect 3988 18834 4016 19858
rect 4632 19378 4660 20334
rect 5368 19990 5396 20402
rect 5356 19984 5408 19990
rect 5356 19926 5408 19932
rect 6564 19854 6592 20742
rect 6552 19848 6604 19854
rect 6552 19790 6604 19796
rect 6748 19786 6776 21490
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 6840 19854 6868 20198
rect 6932 19854 6960 21490
rect 7024 20942 7052 23582
rect 7208 23186 7236 23734
rect 7196 23180 7248 23186
rect 7196 23122 7248 23128
rect 7196 22976 7248 22982
rect 7196 22918 7248 22924
rect 7104 22772 7156 22778
rect 7104 22714 7156 22720
rect 7116 22030 7144 22714
rect 7208 22438 7236 22918
rect 7300 22574 7328 29446
rect 7392 28762 7420 30806
rect 7484 30394 7512 32778
rect 8220 32502 8248 34002
rect 8484 33924 8536 33930
rect 8484 33866 8536 33872
rect 8496 33590 8524 33866
rect 8484 33584 8536 33590
rect 8484 33526 8536 33532
rect 8392 33516 8444 33522
rect 8392 33458 8444 33464
rect 8404 32978 8432 33458
rect 8392 32972 8444 32978
rect 8392 32914 8444 32920
rect 8404 32502 8432 32914
rect 7748 32496 7800 32502
rect 7748 32438 7800 32444
rect 8208 32496 8260 32502
rect 8208 32438 8260 32444
rect 8392 32496 8444 32502
rect 8392 32438 8444 32444
rect 7656 31680 7708 31686
rect 7656 31622 7708 31628
rect 7668 31346 7696 31622
rect 7656 31340 7708 31346
rect 7656 31282 7708 31288
rect 7564 30660 7616 30666
rect 7564 30602 7616 30608
rect 7472 30388 7524 30394
rect 7472 30330 7524 30336
rect 7472 29232 7524 29238
rect 7472 29174 7524 29180
rect 7380 28756 7432 28762
rect 7380 28698 7432 28704
rect 7392 28150 7420 28698
rect 7380 28144 7432 28150
rect 7380 28086 7432 28092
rect 7392 27606 7420 28086
rect 7380 27600 7432 27606
rect 7380 27542 7432 27548
rect 7392 26790 7420 27542
rect 7380 26784 7432 26790
rect 7380 26726 7432 26732
rect 7484 25770 7512 29174
rect 7576 29170 7604 30602
rect 7760 29730 7788 32438
rect 8208 32292 8260 32298
rect 8208 32234 8260 32240
rect 8220 31822 8248 32234
rect 8300 32224 8352 32230
rect 8300 32166 8352 32172
rect 8312 32026 8340 32166
rect 8300 32020 8352 32026
rect 8300 31962 8352 31968
rect 8312 31822 8340 31962
rect 8208 31816 8260 31822
rect 8208 31758 8260 31764
rect 8300 31816 8352 31822
rect 8300 31758 8352 31764
rect 7840 31408 7892 31414
rect 7840 31350 7892 31356
rect 7668 29714 7788 29730
rect 7656 29708 7788 29714
rect 7708 29702 7788 29708
rect 7656 29650 7708 29656
rect 7852 29578 7880 31350
rect 8220 31278 8248 31758
rect 8208 31272 8260 31278
rect 8208 31214 8260 31220
rect 7932 31204 7984 31210
rect 7932 31146 7984 31152
rect 7944 30938 7972 31146
rect 7932 30932 7984 30938
rect 7932 30874 7984 30880
rect 8208 30796 8260 30802
rect 8208 30738 8260 30744
rect 8116 30728 8168 30734
rect 8116 30670 8168 30676
rect 7932 30660 7984 30666
rect 7932 30602 7984 30608
rect 7944 30394 7972 30602
rect 7932 30388 7984 30394
rect 7932 30330 7984 30336
rect 7840 29572 7892 29578
rect 7840 29514 7892 29520
rect 7564 29164 7616 29170
rect 7564 29106 7616 29112
rect 7576 28082 7604 29106
rect 7564 28076 7616 28082
rect 7564 28018 7616 28024
rect 7576 27946 7604 28018
rect 7852 28014 7880 29514
rect 7840 28008 7892 28014
rect 7840 27950 7892 27956
rect 7564 27940 7616 27946
rect 7564 27882 7616 27888
rect 7840 27328 7892 27334
rect 7840 27270 7892 27276
rect 7656 26512 7708 26518
rect 7656 26454 7708 26460
rect 7472 25764 7524 25770
rect 7472 25706 7524 25712
rect 7484 25158 7512 25706
rect 7472 25152 7524 25158
rect 7472 25094 7524 25100
rect 7484 23798 7512 25094
rect 7668 24614 7696 26454
rect 7748 24812 7800 24818
rect 7748 24754 7800 24760
rect 7760 24682 7788 24754
rect 7748 24676 7800 24682
rect 7748 24618 7800 24624
rect 7656 24608 7708 24614
rect 7656 24550 7708 24556
rect 7472 23792 7524 23798
rect 7472 23734 7524 23740
rect 7564 22976 7616 22982
rect 7564 22918 7616 22924
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7288 22568 7340 22574
rect 7288 22510 7340 22516
rect 7196 22432 7248 22438
rect 7196 22374 7248 22380
rect 7300 22094 7328 22510
rect 7484 22234 7512 22578
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7300 22066 7420 22094
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 7116 20806 7144 21966
rect 7196 21956 7248 21962
rect 7196 21898 7248 21904
rect 7208 20942 7236 21898
rect 7196 20936 7248 20942
rect 7196 20878 7248 20884
rect 7104 20800 7156 20806
rect 7104 20742 7156 20748
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7116 20058 7144 20402
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 6920 19848 6972 19854
rect 6920 19790 6972 19796
rect 6736 19780 6788 19786
rect 6736 19722 6788 19728
rect 5632 19440 5684 19446
rect 5632 19382 5684 19388
rect 4620 19372 4672 19378
rect 4620 19314 4672 19320
rect 5080 19168 5132 19174
rect 5080 19110 5132 19116
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3976 18828 4028 18834
rect 3976 18770 4028 18776
rect 5092 18698 5120 19110
rect 5644 18902 5672 19382
rect 6748 19378 6776 19722
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 5632 18896 5684 18902
rect 5632 18838 5684 18844
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 5080 18692 5132 18698
rect 5080 18634 5132 18640
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 5828 17746 5856 18702
rect 6092 18624 6144 18630
rect 6092 18566 6144 18572
rect 5816 17740 5868 17746
rect 5816 17682 5868 17688
rect 6104 17678 6132 18566
rect 6472 18426 6500 18702
rect 6828 18692 6880 18698
rect 6932 18680 6960 19790
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 6880 18652 6960 18680
rect 6828 18634 6880 18640
rect 6460 18420 6512 18426
rect 6460 18362 6512 18368
rect 7116 18290 7144 19246
rect 7392 19242 7420 22066
rect 7472 22024 7524 22030
rect 7472 21966 7524 21972
rect 7484 21690 7512 21966
rect 7576 21894 7604 22918
rect 7564 21888 7616 21894
rect 7564 21830 7616 21836
rect 7472 21684 7524 21690
rect 7472 21626 7524 21632
rect 7668 21434 7696 24550
rect 7852 22710 7880 27270
rect 7944 26042 7972 30330
rect 8128 30190 8156 30670
rect 8116 30184 8168 30190
rect 8116 30126 8168 30132
rect 8128 29646 8156 30126
rect 8220 30054 8248 30738
rect 8208 30048 8260 30054
rect 8208 29990 8260 29996
rect 8116 29640 8168 29646
rect 8116 29582 8168 29588
rect 8588 28626 8616 36246
rect 9324 35766 9352 36246
rect 9312 35760 9364 35766
rect 9312 35702 9364 35708
rect 9416 35562 9444 37266
rect 11716 37262 11744 39200
rect 12164 37324 12216 37330
rect 12164 37266 12216 37272
rect 11704 37256 11756 37262
rect 11704 37198 11756 37204
rect 9496 37188 9548 37194
rect 9496 37130 9548 37136
rect 9508 36242 9536 37130
rect 9588 37120 9640 37126
rect 9588 37062 9640 37068
rect 9600 36922 9628 37062
rect 9588 36916 9640 36922
rect 9588 36858 9640 36864
rect 9496 36236 9548 36242
rect 9496 36178 9548 36184
rect 9600 36038 9628 36858
rect 11520 36780 11572 36786
rect 11520 36722 11572 36728
rect 11532 36310 11560 36722
rect 11520 36304 11572 36310
rect 11520 36246 11572 36252
rect 9680 36168 9732 36174
rect 9680 36110 9732 36116
rect 9588 36032 9640 36038
rect 9588 35974 9640 35980
rect 9404 35556 9456 35562
rect 9404 35498 9456 35504
rect 9588 35488 9640 35494
rect 9588 35430 9640 35436
rect 9600 35018 9628 35430
rect 9692 35086 9720 36110
rect 11704 36100 11756 36106
rect 11704 36042 11756 36048
rect 11716 35834 11744 36042
rect 11888 36032 11940 36038
rect 11888 35974 11940 35980
rect 11900 35834 11928 35974
rect 11704 35828 11756 35834
rect 11704 35770 11756 35776
rect 11888 35828 11940 35834
rect 11888 35770 11940 35776
rect 9956 35692 10008 35698
rect 9956 35634 10008 35640
rect 11612 35692 11664 35698
rect 11612 35634 11664 35640
rect 9680 35080 9732 35086
rect 9680 35022 9732 35028
rect 9588 35012 9640 35018
rect 9588 34954 9640 34960
rect 9692 34066 9720 35022
rect 9968 34678 9996 35634
rect 10048 35624 10100 35630
rect 10048 35566 10100 35572
rect 10060 35290 10088 35566
rect 10048 35284 10100 35290
rect 10048 35226 10100 35232
rect 10060 34746 10088 35226
rect 11336 35216 11388 35222
rect 11336 35158 11388 35164
rect 10048 34740 10100 34746
rect 10048 34682 10100 34688
rect 9956 34672 10008 34678
rect 9956 34614 10008 34620
rect 10232 34196 10284 34202
rect 10232 34138 10284 34144
rect 9680 34060 9732 34066
rect 9680 34002 9732 34008
rect 9128 33924 9180 33930
rect 9128 33866 9180 33872
rect 9140 31414 9168 33866
rect 9312 33584 9364 33590
rect 9312 33526 9364 33532
rect 9220 32904 9272 32910
rect 9220 32846 9272 32852
rect 9232 32570 9260 32846
rect 9220 32564 9272 32570
rect 9220 32506 9272 32512
rect 9220 32428 9272 32434
rect 9220 32370 9272 32376
rect 9232 31793 9260 32370
rect 9218 31784 9274 31793
rect 9218 31719 9274 31728
rect 9128 31408 9180 31414
rect 9128 31350 9180 31356
rect 9220 30728 9272 30734
rect 9220 30670 9272 30676
rect 8668 30252 8720 30258
rect 8668 30194 8720 30200
rect 9036 30252 9088 30258
rect 9036 30194 9088 30200
rect 8680 29510 8708 30194
rect 9048 29850 9076 30194
rect 8760 29844 8812 29850
rect 8760 29786 8812 29792
rect 9036 29844 9088 29850
rect 9036 29786 9088 29792
rect 8668 29504 8720 29510
rect 8668 29446 8720 29452
rect 8772 29170 8800 29786
rect 8760 29164 8812 29170
rect 8760 29106 8812 29112
rect 8576 28620 8628 28626
rect 8576 28562 8628 28568
rect 8300 28552 8352 28558
rect 8300 28494 8352 28500
rect 8482 28520 8538 28529
rect 8116 28484 8168 28490
rect 8116 28426 8168 28432
rect 8024 28416 8076 28422
rect 8024 28358 8076 28364
rect 8036 27538 8064 28358
rect 8128 27674 8156 28426
rect 8312 28082 8340 28494
rect 8482 28455 8484 28464
rect 8536 28455 8538 28464
rect 8484 28426 8536 28432
rect 8484 28212 8536 28218
rect 8484 28154 8536 28160
rect 8300 28076 8352 28082
rect 8300 28018 8352 28024
rect 8300 27872 8352 27878
rect 8300 27814 8352 27820
rect 8116 27668 8168 27674
rect 8116 27610 8168 27616
rect 8024 27532 8076 27538
rect 8024 27474 8076 27480
rect 8116 27396 8168 27402
rect 8116 27338 8168 27344
rect 8128 26994 8156 27338
rect 8116 26988 8168 26994
rect 8116 26930 8168 26936
rect 7932 26036 7984 26042
rect 7932 25978 7984 25984
rect 8208 26036 8260 26042
rect 8208 25978 8260 25984
rect 8116 25696 8168 25702
rect 8116 25638 8168 25644
rect 8024 25424 8076 25430
rect 8024 25366 8076 25372
rect 7932 24336 7984 24342
rect 7932 24278 7984 24284
rect 7840 22704 7892 22710
rect 7840 22646 7892 22652
rect 7944 22094 7972 24278
rect 8036 22574 8064 25366
rect 8128 25294 8156 25638
rect 8116 25288 8168 25294
rect 8116 25230 8168 25236
rect 8128 23730 8156 25230
rect 8220 24886 8248 25978
rect 8208 24880 8260 24886
rect 8208 24822 8260 24828
rect 8312 24154 8340 27814
rect 8496 26994 8524 28154
rect 9048 28082 9076 29786
rect 9232 29646 9260 30670
rect 9324 30258 9352 33526
rect 9956 33312 10008 33318
rect 9956 33254 10008 33260
rect 9680 33040 9732 33046
rect 9968 32994 9996 33254
rect 10244 33114 10272 34138
rect 11348 34066 11376 35158
rect 11624 35018 11652 35634
rect 11900 35578 11928 35770
rect 12176 35698 12204 37266
rect 15028 37244 15056 39200
rect 18340 37262 18368 39200
rect 21652 39114 21680 39200
rect 21744 39114 21772 39222
rect 21652 39086 21772 39114
rect 15200 37256 15252 37262
rect 15028 37216 15200 37244
rect 15200 37198 15252 37204
rect 18328 37256 18380 37262
rect 22020 37244 22048 39222
rect 24950 39200 25006 40000
rect 28262 39200 28318 40000
rect 31574 39200 31630 40000
rect 34886 39200 34942 40000
rect 38198 39200 38254 40000
rect 24964 37262 24992 39200
rect 26516 37324 26568 37330
rect 26516 37266 26568 37272
rect 28080 37324 28132 37330
rect 28080 37266 28132 37272
rect 22100 37256 22152 37262
rect 22020 37216 22100 37244
rect 18328 37198 18380 37204
rect 22100 37198 22152 37204
rect 24952 37256 25004 37262
rect 24952 37198 25004 37204
rect 26240 37256 26292 37262
rect 26240 37198 26292 37204
rect 16028 37188 16080 37194
rect 16028 37130 16080 37136
rect 18604 37188 18656 37194
rect 18604 37130 18656 37136
rect 24308 37188 24360 37194
rect 24308 37130 24360 37136
rect 12992 37120 13044 37126
rect 12992 37062 13044 37068
rect 12624 36780 12676 36786
rect 12624 36722 12676 36728
rect 12636 36378 12664 36722
rect 12624 36372 12676 36378
rect 12624 36314 12676 36320
rect 13004 36174 13032 37062
rect 15292 36848 15344 36854
rect 15292 36790 15344 36796
rect 15844 36848 15896 36854
rect 15844 36790 15896 36796
rect 13360 36780 13412 36786
rect 13360 36722 13412 36728
rect 13084 36576 13136 36582
rect 13084 36518 13136 36524
rect 13096 36242 13124 36518
rect 13084 36236 13136 36242
rect 13084 36178 13136 36184
rect 13268 36236 13320 36242
rect 13268 36178 13320 36184
rect 12716 36168 12768 36174
rect 12716 36110 12768 36116
rect 12992 36168 13044 36174
rect 12992 36110 13044 36116
rect 12164 35692 12216 35698
rect 12164 35634 12216 35640
rect 11808 35550 11928 35578
rect 11808 35018 11836 35550
rect 11888 35216 11940 35222
rect 11888 35158 11940 35164
rect 11900 35018 11928 35158
rect 12728 35154 12756 36110
rect 13096 35154 13124 36178
rect 13280 35834 13308 36178
rect 13268 35828 13320 35834
rect 13268 35770 13320 35776
rect 13280 35562 13308 35770
rect 13372 35698 13400 36722
rect 14556 36712 14608 36718
rect 14556 36654 14608 36660
rect 14004 36304 14056 36310
rect 14004 36246 14056 36252
rect 13544 36236 13596 36242
rect 13544 36178 13596 36184
rect 13360 35692 13412 35698
rect 13360 35634 13412 35640
rect 13268 35556 13320 35562
rect 13268 35498 13320 35504
rect 12716 35148 12768 35154
rect 12716 35090 12768 35096
rect 13084 35148 13136 35154
rect 13084 35090 13136 35096
rect 11612 35012 11664 35018
rect 11612 34954 11664 34960
rect 11796 35012 11848 35018
rect 11796 34954 11848 34960
rect 11888 35012 11940 35018
rect 11888 34954 11940 34960
rect 11336 34060 11388 34066
rect 11336 34002 11388 34008
rect 10600 33992 10652 33998
rect 10600 33934 10652 33940
rect 11152 33992 11204 33998
rect 11152 33934 11204 33940
rect 10232 33108 10284 33114
rect 10232 33050 10284 33056
rect 9680 32982 9732 32988
rect 9588 32768 9640 32774
rect 9588 32710 9640 32716
rect 9600 32570 9628 32710
rect 9588 32564 9640 32570
rect 9588 32506 9640 32512
rect 9496 32428 9548 32434
rect 9496 32370 9548 32376
rect 9508 32337 9536 32370
rect 9494 32328 9550 32337
rect 9494 32263 9550 32272
rect 9692 32230 9720 32982
rect 9784 32978 9996 32994
rect 9772 32972 9996 32978
rect 9824 32966 9996 32972
rect 9772 32914 9824 32920
rect 9864 32904 9916 32910
rect 9864 32846 9916 32852
rect 9680 32224 9732 32230
rect 9680 32166 9732 32172
rect 9588 31272 9640 31278
rect 9588 31214 9640 31220
rect 9404 30932 9456 30938
rect 9404 30874 9456 30880
rect 9312 30252 9364 30258
rect 9312 30194 9364 30200
rect 9220 29640 9272 29646
rect 9220 29582 9272 29588
rect 9232 29102 9260 29582
rect 9220 29096 9272 29102
rect 9220 29038 9272 29044
rect 9128 28960 9180 28966
rect 9128 28902 9180 28908
rect 9220 28960 9272 28966
rect 9220 28902 9272 28908
rect 9140 28558 9168 28902
rect 9232 28762 9260 28902
rect 9220 28756 9272 28762
rect 9220 28698 9272 28704
rect 9128 28552 9180 28558
rect 9128 28494 9180 28500
rect 9128 28416 9180 28422
rect 9128 28358 9180 28364
rect 9036 28076 9088 28082
rect 9036 28018 9088 28024
rect 9036 27396 9088 27402
rect 9140 27384 9168 28358
rect 9312 28144 9364 28150
rect 9312 28086 9364 28092
rect 9220 27464 9272 27470
rect 9220 27406 9272 27412
rect 9088 27356 9168 27384
rect 9036 27338 9088 27344
rect 8484 26988 8536 26994
rect 8484 26930 8536 26936
rect 8496 26314 8524 26930
rect 8668 26852 8720 26858
rect 8668 26794 8720 26800
rect 8484 26308 8536 26314
rect 8484 26250 8536 26256
rect 8392 26240 8444 26246
rect 8392 26182 8444 26188
rect 8404 25498 8432 26182
rect 8484 25900 8536 25906
rect 8484 25842 8536 25848
rect 8392 25492 8444 25498
rect 8392 25434 8444 25440
rect 8392 25288 8444 25294
rect 8496 25276 8524 25842
rect 8444 25248 8524 25276
rect 8392 25230 8444 25236
rect 8404 24954 8432 25230
rect 8392 24948 8444 24954
rect 8392 24890 8444 24896
rect 8404 24410 8432 24890
rect 8576 24744 8628 24750
rect 8576 24686 8628 24692
rect 8392 24404 8444 24410
rect 8392 24346 8444 24352
rect 8220 24138 8340 24154
rect 8208 24132 8340 24138
rect 8260 24126 8340 24132
rect 8208 24074 8260 24080
rect 8300 24064 8352 24070
rect 8220 24012 8300 24018
rect 8220 24006 8352 24012
rect 8220 23990 8340 24006
rect 8116 23724 8168 23730
rect 8116 23666 8168 23672
rect 8220 23594 8248 23990
rect 8392 23724 8444 23730
rect 8392 23666 8444 23672
rect 8208 23588 8260 23594
rect 8208 23530 8260 23536
rect 8024 22568 8076 22574
rect 8024 22510 8076 22516
rect 8116 22432 8168 22438
rect 8116 22374 8168 22380
rect 7852 22066 7972 22094
rect 7852 22030 7880 22066
rect 7840 22024 7892 22030
rect 7840 21966 7892 21972
rect 7932 22024 7984 22030
rect 7932 21966 7984 21972
rect 7576 21406 7696 21434
rect 7852 21418 7880 21966
rect 7944 21486 7972 21966
rect 8128 21486 8156 22374
rect 8220 21554 8248 23530
rect 8404 22030 8432 23666
rect 8588 23526 8616 24686
rect 8680 23662 8708 26794
rect 9048 25140 9076 27338
rect 9128 26920 9180 26926
rect 9128 26862 9180 26868
rect 9140 26586 9168 26862
rect 9232 26790 9260 27406
rect 9220 26784 9272 26790
rect 9218 26752 9220 26761
rect 9272 26752 9274 26761
rect 9218 26687 9274 26696
rect 9324 26602 9352 28086
rect 9416 28082 9444 30874
rect 9600 30326 9628 31214
rect 9692 30394 9720 32166
rect 9876 32026 9904 32846
rect 9864 32020 9916 32026
rect 9864 31962 9916 31968
rect 9968 31822 9996 32966
rect 10140 32972 10192 32978
rect 10140 32914 10192 32920
rect 10152 32026 10180 32914
rect 10244 32910 10272 33050
rect 10232 32904 10284 32910
rect 10232 32846 10284 32852
rect 10244 32434 10272 32846
rect 10612 32842 10640 33934
rect 11164 32910 11192 33934
rect 11348 33454 11376 34002
rect 11336 33448 11388 33454
rect 11336 33390 11388 33396
rect 11348 32994 11376 33390
rect 11256 32978 11376 32994
rect 11244 32972 11376 32978
rect 11296 32966 11376 32972
rect 11244 32914 11296 32920
rect 11152 32904 11204 32910
rect 11152 32846 11204 32852
rect 10600 32836 10652 32842
rect 10600 32778 10652 32784
rect 10416 32768 10468 32774
rect 10416 32710 10468 32716
rect 10428 32570 10456 32710
rect 10416 32564 10468 32570
rect 10416 32506 10468 32512
rect 10232 32428 10284 32434
rect 10232 32370 10284 32376
rect 10324 32292 10376 32298
rect 10324 32234 10376 32240
rect 10140 32020 10192 32026
rect 10140 31962 10192 31968
rect 10048 31884 10100 31890
rect 10048 31826 10100 31832
rect 9772 31816 9824 31822
rect 9772 31758 9824 31764
rect 9956 31816 10008 31822
rect 9956 31758 10008 31764
rect 9784 31142 9812 31758
rect 9864 31680 9916 31686
rect 9864 31622 9916 31628
rect 9772 31136 9824 31142
rect 9772 31078 9824 31084
rect 9876 30954 9904 31622
rect 9784 30926 9904 30954
rect 9680 30388 9732 30394
rect 9680 30330 9732 30336
rect 9588 30320 9640 30326
rect 9640 30268 9720 30274
rect 9588 30262 9720 30268
rect 9600 30246 9720 30262
rect 9600 30197 9628 30246
rect 9588 29164 9640 29170
rect 9588 29106 9640 29112
rect 9600 28150 9628 29106
rect 9588 28144 9640 28150
rect 9588 28086 9640 28092
rect 9404 28076 9456 28082
rect 9404 28018 9456 28024
rect 9416 27538 9444 28018
rect 9404 27532 9456 27538
rect 9404 27474 9456 27480
rect 9586 27432 9642 27441
rect 9128 26580 9180 26586
rect 9128 26522 9180 26528
rect 9232 26574 9352 26602
rect 9416 27376 9586 27384
rect 9416 27356 9588 27376
rect 9232 25906 9260 26574
rect 9416 26058 9444 27356
rect 9640 27367 9642 27376
rect 9588 27338 9640 27344
rect 9588 26852 9640 26858
rect 9588 26794 9640 26800
rect 9494 26480 9550 26489
rect 9494 26415 9550 26424
rect 9508 26360 9536 26415
rect 9496 26354 9548 26360
rect 9600 26314 9628 26794
rect 9692 26518 9720 30246
rect 9784 29102 9812 30926
rect 9864 30592 9916 30598
rect 9864 30534 9916 30540
rect 9876 29170 9904 30534
rect 10060 30258 10088 31826
rect 10232 31816 10284 31822
rect 10232 31758 10284 31764
rect 10244 30938 10272 31758
rect 10336 31346 10364 32234
rect 10612 31822 10640 32778
rect 11060 32768 11112 32774
rect 11060 32710 11112 32716
rect 11072 32230 11100 32710
rect 11060 32224 11112 32230
rect 11060 32166 11112 32172
rect 10600 31816 10652 31822
rect 10414 31784 10470 31793
rect 10600 31758 10652 31764
rect 10414 31719 10470 31728
rect 10324 31340 10376 31346
rect 10324 31282 10376 31288
rect 10232 30932 10284 30938
rect 10232 30874 10284 30880
rect 10324 30388 10376 30394
rect 10324 30330 10376 30336
rect 10048 30252 10100 30258
rect 10048 30194 10100 30200
rect 10140 30252 10192 30258
rect 10140 30194 10192 30200
rect 9956 29640 10008 29646
rect 9956 29582 10008 29588
rect 9864 29164 9916 29170
rect 9864 29106 9916 29112
rect 9772 29096 9824 29102
rect 9772 29038 9824 29044
rect 9876 28014 9904 29106
rect 9864 28008 9916 28014
rect 9864 27950 9916 27956
rect 9968 27606 9996 29582
rect 9956 27600 10008 27606
rect 9956 27542 10008 27548
rect 9864 27396 9916 27402
rect 9864 27338 9916 27344
rect 9876 26858 9904 27338
rect 9968 26994 9996 27542
rect 9956 26988 10008 26994
rect 9956 26930 10008 26936
rect 9864 26852 9916 26858
rect 9864 26794 9916 26800
rect 9680 26512 9732 26518
rect 9680 26454 9732 26460
rect 9772 26512 9824 26518
rect 9772 26454 9824 26460
rect 9496 26296 9548 26302
rect 9588 26308 9640 26314
rect 9588 26250 9640 26256
rect 9324 26030 9444 26058
rect 9220 25900 9272 25906
rect 9220 25842 9272 25848
rect 9324 25702 9352 26030
rect 9404 25968 9456 25974
rect 9404 25910 9456 25916
rect 9312 25696 9364 25702
rect 9312 25638 9364 25644
rect 9220 25152 9272 25158
rect 9048 25112 9220 25140
rect 9220 25094 9272 25100
rect 9232 24206 9260 25094
rect 9312 24812 9364 24818
rect 9312 24754 9364 24760
rect 9324 24614 9352 24754
rect 9312 24608 9364 24614
rect 9312 24550 9364 24556
rect 8760 24200 8812 24206
rect 8760 24142 8812 24148
rect 9220 24200 9272 24206
rect 9220 24142 9272 24148
rect 8668 23656 8720 23662
rect 8668 23598 8720 23604
rect 8576 23520 8628 23526
rect 8576 23462 8628 23468
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8588 21894 8616 23462
rect 8680 23118 8708 23598
rect 8668 23112 8720 23118
rect 8668 23054 8720 23060
rect 8680 22642 8708 23054
rect 8668 22636 8720 22642
rect 8668 22578 8720 22584
rect 8576 21888 8628 21894
rect 8576 21830 8628 21836
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 7932 21480 7984 21486
rect 7932 21422 7984 21428
rect 8116 21480 8168 21486
rect 8116 21422 8168 21428
rect 7840 21412 7892 21418
rect 7380 19236 7432 19242
rect 7380 19178 7432 19184
rect 7576 18766 7604 21406
rect 7840 21354 7892 21360
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7196 18692 7248 18698
rect 7196 18634 7248 18640
rect 7380 18692 7432 18698
rect 7380 18634 7432 18640
rect 7104 18284 7156 18290
rect 7104 18226 7156 18232
rect 6092 17672 6144 17678
rect 6092 17614 6144 17620
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 6552 16516 6604 16522
rect 6552 16458 6604 16464
rect 6564 16250 6592 16458
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 6932 15706 6960 16526
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7024 16182 7052 16390
rect 7012 16176 7064 16182
rect 7012 16118 7064 16124
rect 7116 16046 7144 18226
rect 7208 17542 7236 18634
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7208 17338 7236 17478
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 6932 14482 6960 15642
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 7392 14414 7420 18634
rect 7668 17270 7696 21286
rect 7932 18216 7984 18222
rect 7932 18158 7984 18164
rect 7656 17264 7708 17270
rect 7656 17206 7708 17212
rect 7840 17128 7892 17134
rect 7840 17070 7892 17076
rect 7852 16658 7880 17070
rect 7944 16726 7972 18158
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 8036 16794 8064 17138
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 7932 16720 7984 16726
rect 7932 16662 7984 16668
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 8128 16114 8156 21422
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 8220 19242 8248 19790
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8208 19236 8260 19242
rect 8208 19178 8260 19184
rect 8220 17202 8248 19178
rect 8404 18698 8432 19654
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8392 18692 8444 18698
rect 8392 18634 8444 18640
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8220 16590 8248 16730
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 8404 16250 8432 18634
rect 8588 18358 8616 19110
rect 8772 18426 8800 24142
rect 9324 24138 9352 24550
rect 9416 24410 9444 25910
rect 9680 25356 9732 25362
rect 9680 25298 9732 25304
rect 9496 25152 9548 25158
rect 9496 25094 9548 25100
rect 9404 24404 9456 24410
rect 9404 24346 9456 24352
rect 9312 24132 9364 24138
rect 9312 24074 9364 24080
rect 9312 23588 9364 23594
rect 9312 23530 9364 23536
rect 9128 23112 9180 23118
rect 9128 23054 9180 23060
rect 8944 23044 8996 23050
rect 8944 22986 8996 22992
rect 8956 22778 8984 22986
rect 8944 22772 8996 22778
rect 8944 22714 8996 22720
rect 9140 20942 9168 23054
rect 9324 22574 9352 23530
rect 9312 22568 9364 22574
rect 9312 22510 9364 22516
rect 9324 22166 9352 22510
rect 9312 22160 9364 22166
rect 9312 22102 9364 22108
rect 9220 22024 9272 22030
rect 9220 21966 9272 21972
rect 9232 21486 9260 21966
rect 9404 21684 9456 21690
rect 9404 21626 9456 21632
rect 9220 21480 9272 21486
rect 9220 21422 9272 21428
rect 9220 21344 9272 21350
rect 9220 21286 9272 21292
rect 9232 21010 9260 21286
rect 9220 21004 9272 21010
rect 9220 20946 9272 20952
rect 9128 20936 9180 20942
rect 9128 20878 9180 20884
rect 9140 19378 9168 20878
rect 9232 20534 9260 20946
rect 9220 20528 9272 20534
rect 9220 20470 9272 20476
rect 9416 20466 9444 21626
rect 9404 20460 9456 20466
rect 9404 20402 9456 20408
rect 9508 19514 9536 25094
rect 9692 24750 9720 25298
rect 9784 24818 9812 26454
rect 9864 26376 9916 26382
rect 9864 26318 9916 26324
rect 9876 26042 9904 26318
rect 9864 26036 9916 26042
rect 9864 25978 9916 25984
rect 9968 25906 9996 26930
rect 9956 25900 10008 25906
rect 9956 25842 10008 25848
rect 9772 24812 9824 24818
rect 9772 24754 9824 24760
rect 9680 24744 9732 24750
rect 9680 24686 9732 24692
rect 9692 23730 9720 24686
rect 9864 24608 9916 24614
rect 9864 24550 9916 24556
rect 9680 23724 9732 23730
rect 9680 23666 9732 23672
rect 9876 22982 9904 24550
rect 9864 22976 9916 22982
rect 9864 22918 9916 22924
rect 9876 22681 9904 22918
rect 9862 22672 9918 22681
rect 9862 22607 9918 22616
rect 10060 21962 10088 30194
rect 10152 29306 10180 30194
rect 10140 29300 10192 29306
rect 10140 29242 10192 29248
rect 10232 29164 10284 29170
rect 10232 29106 10284 29112
rect 10140 29096 10192 29102
rect 10140 29038 10192 29044
rect 10152 28014 10180 29038
rect 10244 28082 10272 29106
rect 10232 28076 10284 28082
rect 10232 28018 10284 28024
rect 10140 28008 10192 28014
rect 10140 27950 10192 27956
rect 10152 27334 10180 27950
rect 10336 27878 10364 30330
rect 10428 28490 10456 31719
rect 10600 31680 10652 31686
rect 10600 31622 10652 31628
rect 10612 31346 10640 31622
rect 10600 31340 10652 31346
rect 10600 31282 10652 31288
rect 10508 31136 10560 31142
rect 10508 31078 10560 31084
rect 10520 29850 10548 31078
rect 10612 30870 10640 31282
rect 11072 31278 11100 32166
rect 11164 31754 11192 32846
rect 11520 32292 11572 32298
rect 11520 32234 11572 32240
rect 11532 32026 11560 32234
rect 11520 32020 11572 32026
rect 11520 31962 11572 31968
rect 11624 31793 11652 34954
rect 11900 34542 11928 34954
rect 12716 34944 12768 34950
rect 12716 34886 12768 34892
rect 11888 34536 11940 34542
rect 11888 34478 11940 34484
rect 11888 33992 11940 33998
rect 11888 33934 11940 33940
rect 12256 33992 12308 33998
rect 12256 33934 12308 33940
rect 11900 32502 11928 33934
rect 12268 33522 12296 33934
rect 12072 33516 12124 33522
rect 12072 33458 12124 33464
rect 12256 33516 12308 33522
rect 12256 33458 12308 33464
rect 11980 32836 12032 32842
rect 11980 32778 12032 32784
rect 11888 32496 11940 32502
rect 11888 32438 11940 32444
rect 11704 31816 11756 31822
rect 11610 31784 11666 31793
rect 11152 31748 11204 31754
rect 11152 31690 11204 31696
rect 11520 31748 11572 31754
rect 11756 31776 11836 31804
rect 11704 31758 11756 31764
rect 11610 31719 11666 31728
rect 11520 31690 11572 31696
rect 11060 31272 11112 31278
rect 11060 31214 11112 31220
rect 10600 30864 10652 30870
rect 10600 30806 10652 30812
rect 11072 30802 11100 31214
rect 11060 30796 11112 30802
rect 11060 30738 11112 30744
rect 11152 30592 11204 30598
rect 11152 30534 11204 30540
rect 10508 29844 10560 29850
rect 10508 29786 10560 29792
rect 11164 29034 11192 30534
rect 11532 29170 11560 31690
rect 11808 31346 11836 31776
rect 11900 31482 11928 32438
rect 11992 32366 12020 32778
rect 12084 32434 12112 33458
rect 12268 32910 12296 33458
rect 12256 32904 12308 32910
rect 12532 32904 12584 32910
rect 12308 32864 12480 32892
rect 12256 32846 12308 32852
rect 12256 32496 12308 32502
rect 12256 32438 12308 32444
rect 12072 32428 12124 32434
rect 12072 32370 12124 32376
rect 11980 32360 12032 32366
rect 11980 32302 12032 32308
rect 11980 31952 12032 31958
rect 11980 31894 12032 31900
rect 11888 31476 11940 31482
rect 11888 31418 11940 31424
rect 11796 31340 11848 31346
rect 11796 31282 11848 31288
rect 11704 31136 11756 31142
rect 11704 31078 11756 31084
rect 11716 30734 11744 31078
rect 11704 30728 11756 30734
rect 11704 30670 11756 30676
rect 11808 30394 11836 31282
rect 11888 31204 11940 31210
rect 11888 31146 11940 31152
rect 11796 30388 11848 30394
rect 11796 30330 11848 30336
rect 11900 30138 11928 31146
rect 11992 30734 12020 31894
rect 12084 30938 12112 32370
rect 12164 32360 12216 32366
rect 12164 32302 12216 32308
rect 12176 31929 12204 32302
rect 12162 31920 12218 31929
rect 12162 31855 12218 31864
rect 12162 31784 12218 31793
rect 12162 31719 12218 31728
rect 12072 30932 12124 30938
rect 12072 30874 12124 30880
rect 11980 30728 12032 30734
rect 11980 30670 12032 30676
rect 11992 30326 12020 30670
rect 11980 30320 12032 30326
rect 11980 30262 12032 30268
rect 11980 30184 12032 30190
rect 11900 30132 11980 30138
rect 11900 30126 12032 30132
rect 11900 30110 12020 30126
rect 11796 29844 11848 29850
rect 11796 29786 11848 29792
rect 11704 29572 11756 29578
rect 11704 29514 11756 29520
rect 11520 29164 11572 29170
rect 11520 29106 11572 29112
rect 11612 29164 11664 29170
rect 11612 29106 11664 29112
rect 11152 29028 11204 29034
rect 11152 28970 11204 28976
rect 11060 28756 11112 28762
rect 11060 28698 11112 28704
rect 10416 28484 10468 28490
rect 10416 28426 10468 28432
rect 10968 28484 11020 28490
rect 10968 28426 11020 28432
rect 10324 27872 10376 27878
rect 10324 27814 10376 27820
rect 10140 27328 10192 27334
rect 10140 27270 10192 27276
rect 10152 26518 10180 27270
rect 10140 26512 10192 26518
rect 10140 26454 10192 26460
rect 10336 25498 10364 27814
rect 10600 27328 10652 27334
rect 10600 27270 10652 27276
rect 10508 26444 10560 26450
rect 10508 26386 10560 26392
rect 10324 25492 10376 25498
rect 10324 25434 10376 25440
rect 10232 24744 10284 24750
rect 10232 24686 10284 24692
rect 10140 24608 10192 24614
rect 10140 24550 10192 24556
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 10048 21956 10100 21962
rect 10048 21898 10100 21904
rect 9588 21344 9640 21350
rect 9588 21286 9640 21292
rect 9600 21146 9628 21286
rect 9588 21140 9640 21146
rect 9588 21082 9640 21088
rect 9692 19922 9720 21898
rect 9772 21548 9824 21554
rect 9772 21490 9824 21496
rect 9784 20466 9812 21490
rect 9956 20868 10008 20874
rect 9956 20810 10008 20816
rect 9968 20602 9996 20810
rect 9956 20596 10008 20602
rect 9956 20538 10008 20544
rect 9772 20460 9824 20466
rect 9772 20402 9824 20408
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9772 19780 9824 19786
rect 9772 19722 9824 19728
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 9312 19440 9364 19446
rect 9312 19382 9364 19388
rect 9128 19372 9180 19378
rect 9128 19314 9180 19320
rect 9140 18834 9168 19314
rect 9324 18902 9352 19382
rect 9312 18896 9364 18902
rect 9312 18838 9364 18844
rect 9128 18828 9180 18834
rect 9128 18770 9180 18776
rect 8760 18420 8812 18426
rect 8760 18362 8812 18368
rect 8576 18352 8628 18358
rect 8576 18294 8628 18300
rect 9140 17746 9168 18770
rect 9324 18426 9352 18838
rect 9508 18766 9536 19450
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9692 18222 9720 19110
rect 9784 18766 9812 19722
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 9968 18970 9996 19314
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 8668 16992 8720 16998
rect 8668 16934 8720 16940
rect 8680 16590 8708 16934
rect 8668 16584 8720 16590
rect 8668 16526 8720 16532
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 7760 15502 7788 15846
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 8312 14958 8340 15846
rect 8404 15706 8432 15982
rect 8392 15700 8444 15706
rect 8392 15642 8444 15648
rect 10048 15428 10100 15434
rect 10048 15370 10100 15376
rect 8850 15192 8906 15201
rect 10060 15162 10088 15370
rect 8850 15127 8852 15136
rect 8904 15127 8906 15136
rect 10048 15156 10100 15162
rect 8852 15098 8904 15104
rect 10048 15098 10100 15104
rect 10152 15026 10180 24550
rect 10244 24070 10272 24686
rect 10416 24404 10468 24410
rect 10416 24346 10468 24352
rect 10232 24064 10284 24070
rect 10232 24006 10284 24012
rect 10244 19854 10272 24006
rect 10428 22710 10456 24346
rect 10520 24274 10548 26386
rect 10612 25906 10640 27270
rect 10980 26926 11008 28426
rect 11072 28218 11100 28698
rect 11164 28626 11192 28970
rect 11152 28620 11204 28626
rect 11152 28562 11204 28568
rect 11624 28422 11652 29106
rect 11716 28472 11744 29514
rect 11808 29306 11836 29786
rect 11992 29646 12020 30110
rect 12072 29776 12124 29782
rect 12072 29718 12124 29724
rect 11980 29640 12032 29646
rect 11980 29582 12032 29588
rect 11980 29504 12032 29510
rect 11980 29446 12032 29452
rect 11796 29300 11848 29306
rect 11796 29242 11848 29248
rect 11888 29164 11940 29170
rect 11888 29106 11940 29112
rect 11900 28762 11928 29106
rect 11992 28762 12020 29446
rect 11888 28756 11940 28762
rect 11888 28698 11940 28704
rect 11980 28756 12032 28762
rect 11980 28698 12032 28704
rect 11796 28484 11848 28490
rect 11716 28444 11796 28472
rect 11796 28426 11848 28432
rect 11612 28416 11664 28422
rect 11612 28358 11664 28364
rect 11808 28218 11836 28426
rect 11060 28212 11112 28218
rect 11060 28154 11112 28160
rect 11796 28212 11848 28218
rect 11796 28154 11848 28160
rect 11428 27940 11480 27946
rect 11428 27882 11480 27888
rect 11440 27470 11468 27882
rect 11428 27464 11480 27470
rect 11992 27418 12020 28698
rect 12084 28014 12112 29718
rect 12072 28008 12124 28014
rect 12072 27950 12124 27956
rect 11428 27406 11480 27412
rect 11796 27396 11848 27402
rect 11796 27338 11848 27344
rect 11900 27390 12020 27418
rect 11244 27328 11296 27334
rect 11244 27270 11296 27276
rect 10968 26920 11020 26926
rect 10968 26862 11020 26868
rect 10784 26852 10836 26858
rect 10784 26794 10836 26800
rect 10600 25900 10652 25906
rect 10600 25842 10652 25848
rect 10600 25696 10652 25702
rect 10600 25638 10652 25644
rect 10612 25294 10640 25638
rect 10600 25288 10652 25294
rect 10600 25230 10652 25236
rect 10612 24818 10640 25230
rect 10600 24812 10652 24818
rect 10600 24754 10652 24760
rect 10796 24698 10824 26794
rect 10876 26784 10928 26790
rect 10876 26726 10928 26732
rect 10888 26382 10916 26726
rect 11256 26586 11284 27270
rect 11244 26580 11296 26586
rect 11244 26522 11296 26528
rect 11808 26450 11836 27338
rect 11900 26858 11928 27390
rect 11980 26988 12032 26994
rect 11980 26930 12032 26936
rect 11888 26852 11940 26858
rect 11888 26794 11940 26800
rect 11992 26586 12020 26930
rect 11980 26580 12032 26586
rect 11980 26522 12032 26528
rect 11796 26444 11848 26450
rect 11796 26386 11848 26392
rect 10876 26376 10928 26382
rect 10876 26318 10928 26324
rect 10876 25900 10928 25906
rect 10876 25842 10928 25848
rect 10888 25294 10916 25842
rect 10876 25288 10928 25294
rect 10876 25230 10928 25236
rect 10888 24818 10916 25230
rect 10876 24812 10928 24818
rect 10876 24754 10928 24760
rect 11152 24812 11204 24818
rect 11152 24754 11204 24760
rect 10796 24670 10916 24698
rect 10508 24268 10560 24274
rect 10508 24210 10560 24216
rect 10600 23520 10652 23526
rect 10600 23462 10652 23468
rect 10692 23520 10744 23526
rect 10692 23462 10744 23468
rect 10416 22704 10468 22710
rect 10416 22646 10468 22652
rect 10612 22642 10640 23462
rect 10704 23322 10732 23462
rect 10692 23316 10744 23322
rect 10692 23258 10744 23264
rect 10600 22636 10652 22642
rect 10600 22578 10652 22584
rect 10600 22432 10652 22438
rect 10600 22374 10652 22380
rect 10612 21962 10640 22374
rect 10600 21956 10652 21962
rect 10600 21898 10652 21904
rect 10692 21140 10744 21146
rect 10692 21082 10744 21088
rect 10414 20360 10470 20369
rect 10414 20295 10470 20304
rect 10428 19990 10456 20295
rect 10416 19984 10468 19990
rect 10416 19926 10468 19932
rect 10232 19848 10284 19854
rect 10600 19848 10652 19854
rect 10232 19790 10284 19796
rect 10336 19796 10600 19802
rect 10336 19790 10652 19796
rect 10244 18426 10272 19790
rect 10336 19786 10640 19790
rect 10324 19780 10640 19786
rect 10376 19774 10640 19780
rect 10324 19722 10376 19728
rect 10612 19378 10640 19774
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 10428 18290 10456 18702
rect 10416 18284 10468 18290
rect 10416 18226 10468 18232
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 10612 17678 10640 18022
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10508 17264 10560 17270
rect 10508 17206 10560 17212
rect 10520 16794 10548 17206
rect 10508 16788 10560 16794
rect 10508 16730 10560 16736
rect 10520 15042 10548 16730
rect 10704 16522 10732 21082
rect 10784 19236 10836 19242
rect 10784 19178 10836 19184
rect 10796 18698 10824 19178
rect 10784 18692 10836 18698
rect 10784 18634 10836 18640
rect 10888 16726 10916 24670
rect 10968 24608 11020 24614
rect 10968 24550 11020 24556
rect 10980 24206 11008 24550
rect 10968 24200 11020 24206
rect 10968 24142 11020 24148
rect 11164 23730 11192 24754
rect 12072 24744 12124 24750
rect 12072 24686 12124 24692
rect 12084 24410 12112 24686
rect 12072 24404 12124 24410
rect 12072 24346 12124 24352
rect 11152 23724 11204 23730
rect 11152 23666 11204 23672
rect 11164 22642 11192 23666
rect 12072 22976 12124 22982
rect 12072 22918 12124 22924
rect 12084 22710 12112 22918
rect 11704 22704 11756 22710
rect 12072 22704 12124 22710
rect 11704 22646 11756 22652
rect 11794 22672 11850 22681
rect 11152 22636 11204 22642
rect 11152 22578 11204 22584
rect 11716 22234 11744 22646
rect 12072 22646 12124 22652
rect 11794 22607 11796 22616
rect 11848 22607 11850 22616
rect 11796 22578 11848 22584
rect 11704 22228 11756 22234
rect 11704 22170 11756 22176
rect 11888 22228 11940 22234
rect 11888 22170 11940 22176
rect 11900 21622 11928 22170
rect 12176 22094 12204 31719
rect 12268 31278 12296 32438
rect 12348 32224 12400 32230
rect 12348 32166 12400 32172
rect 12360 32026 12388 32166
rect 12348 32020 12400 32026
rect 12348 31962 12400 31968
rect 12346 31920 12402 31929
rect 12346 31855 12402 31864
rect 12360 31822 12388 31855
rect 12348 31816 12400 31822
rect 12348 31758 12400 31764
rect 12360 31346 12388 31758
rect 12452 31346 12480 32864
rect 12532 32846 12584 32852
rect 12348 31340 12400 31346
rect 12348 31282 12400 31288
rect 12440 31340 12492 31346
rect 12440 31282 12492 31288
rect 12256 31272 12308 31278
rect 12256 31214 12308 31220
rect 12268 29850 12296 31214
rect 12360 30734 12388 31282
rect 12452 30870 12480 31282
rect 12440 30864 12492 30870
rect 12440 30806 12492 30812
rect 12348 30728 12400 30734
rect 12348 30670 12400 30676
rect 12256 29844 12308 29850
rect 12256 29786 12308 29792
rect 12360 29628 12388 30670
rect 12544 30598 12572 32846
rect 12622 32464 12678 32473
rect 12622 32399 12678 32408
rect 12636 32366 12664 32399
rect 12624 32360 12676 32366
rect 12624 32302 12676 32308
rect 12624 31816 12676 31822
rect 12624 31758 12676 31764
rect 12636 31686 12664 31758
rect 12624 31680 12676 31686
rect 12624 31622 12676 31628
rect 12532 30592 12584 30598
rect 12532 30534 12584 30540
rect 12532 29640 12584 29646
rect 12360 29600 12532 29628
rect 12532 29582 12584 29588
rect 12440 28960 12492 28966
rect 12440 28902 12492 28908
rect 12256 26444 12308 26450
rect 12256 26386 12308 26392
rect 12268 22642 12296 26386
rect 12452 23526 12480 28902
rect 12728 28422 12756 34886
rect 13372 32978 13400 35634
rect 13556 35086 13584 36178
rect 13636 35624 13688 35630
rect 13636 35566 13688 35572
rect 13544 35080 13596 35086
rect 13544 35022 13596 35028
rect 13648 33658 13676 35566
rect 13636 33652 13688 33658
rect 13636 33594 13688 33600
rect 13544 33448 13596 33454
rect 13544 33390 13596 33396
rect 13556 33114 13584 33390
rect 14016 33130 14044 36246
rect 14096 33856 14148 33862
rect 14096 33798 14148 33804
rect 14108 33318 14136 33798
rect 14568 33522 14596 36654
rect 15304 36378 15332 36790
rect 15292 36372 15344 36378
rect 15292 36314 15344 36320
rect 15856 36242 15884 36790
rect 15844 36236 15896 36242
rect 15844 36178 15896 36184
rect 15200 36168 15252 36174
rect 15200 36110 15252 36116
rect 14740 35692 14792 35698
rect 14740 35634 14792 35640
rect 14752 35290 14780 35634
rect 14832 35488 14884 35494
rect 14832 35430 14884 35436
rect 14740 35284 14792 35290
rect 14740 35226 14792 35232
rect 14648 33992 14700 33998
rect 14648 33934 14700 33940
rect 14660 33658 14688 33934
rect 14844 33844 14872 35430
rect 15212 35086 15240 36110
rect 15856 35170 15884 36178
rect 15764 35154 15884 35170
rect 15752 35148 15884 35154
rect 15804 35142 15884 35148
rect 15752 35090 15804 35096
rect 15200 35080 15252 35086
rect 15200 35022 15252 35028
rect 15936 35012 15988 35018
rect 15936 34954 15988 34960
rect 15844 33992 15896 33998
rect 15844 33934 15896 33940
rect 14752 33816 14872 33844
rect 15476 33856 15528 33862
rect 14648 33652 14700 33658
rect 14648 33594 14700 33600
rect 14188 33516 14240 33522
rect 14188 33458 14240 33464
rect 14556 33516 14608 33522
rect 14556 33458 14608 33464
rect 14200 33318 14228 33458
rect 14372 33448 14424 33454
rect 14372 33390 14424 33396
rect 14648 33448 14700 33454
rect 14648 33390 14700 33396
rect 14096 33312 14148 33318
rect 14096 33254 14148 33260
rect 14188 33312 14240 33318
rect 14188 33254 14240 33260
rect 13544 33108 13596 33114
rect 13544 33050 13596 33056
rect 13728 33108 13780 33114
rect 14016 33102 14136 33130
rect 13728 33050 13780 33056
rect 13360 32972 13412 32978
rect 13360 32914 13412 32920
rect 13556 32910 13584 33050
rect 13740 32910 13768 33050
rect 13544 32904 13596 32910
rect 13544 32846 13596 32852
rect 13728 32904 13780 32910
rect 13728 32846 13780 32852
rect 12808 32836 12860 32842
rect 12808 32778 12860 32784
rect 13820 32836 13872 32842
rect 13820 32778 13872 32784
rect 12820 32230 12848 32778
rect 12900 32360 12952 32366
rect 12900 32302 12952 32308
rect 13542 32328 13598 32337
rect 12808 32224 12860 32230
rect 12808 32166 12860 32172
rect 12912 31822 12940 32302
rect 13542 32263 13598 32272
rect 12900 31816 12952 31822
rect 12900 31758 12952 31764
rect 12808 31680 12860 31686
rect 12808 31622 12860 31628
rect 12820 30666 12848 31622
rect 12912 31482 12940 31758
rect 12900 31476 12952 31482
rect 12900 31418 12952 31424
rect 12992 31340 13044 31346
rect 12992 31282 13044 31288
rect 13004 30938 13032 31282
rect 12992 30932 13044 30938
rect 12992 30874 13044 30880
rect 13360 30728 13412 30734
rect 13360 30670 13412 30676
rect 12808 30660 12860 30666
rect 12808 30602 12860 30608
rect 13176 30184 13228 30190
rect 13176 30126 13228 30132
rect 13268 30184 13320 30190
rect 13268 30126 13320 30132
rect 12808 30116 12860 30122
rect 12808 30058 12860 30064
rect 12820 29170 12848 30058
rect 13188 29578 13216 30126
rect 13176 29572 13228 29578
rect 13176 29514 13228 29520
rect 12808 29164 12860 29170
rect 12808 29106 12860 29112
rect 13084 29028 13136 29034
rect 13280 29016 13308 30126
rect 13372 29646 13400 30670
rect 13556 30666 13584 32263
rect 13832 31754 13860 32778
rect 13648 31726 13860 31754
rect 13648 31414 13676 31726
rect 13636 31408 13688 31414
rect 13636 31350 13688 31356
rect 13544 30660 13596 30666
rect 13544 30602 13596 30608
rect 13360 29640 13412 29646
rect 13360 29582 13412 29588
rect 13136 28988 13308 29016
rect 13084 28970 13136 28976
rect 13372 28626 13400 29582
rect 13648 29170 13676 31350
rect 13820 31204 13872 31210
rect 13820 31146 13872 31152
rect 13728 30796 13780 30802
rect 13728 30738 13780 30744
rect 13740 30705 13768 30738
rect 13726 30696 13782 30705
rect 13726 30631 13782 30640
rect 13832 30054 13860 31146
rect 13912 30252 13964 30258
rect 13912 30194 13964 30200
rect 13820 30048 13872 30054
rect 13820 29990 13872 29996
rect 13636 29164 13688 29170
rect 13636 29106 13688 29112
rect 13544 28688 13596 28694
rect 13544 28630 13596 28636
rect 13360 28620 13412 28626
rect 13360 28562 13412 28568
rect 12716 28416 12768 28422
rect 12716 28358 12768 28364
rect 13268 28416 13320 28422
rect 13268 28358 13320 28364
rect 12728 28082 12756 28358
rect 13280 28150 13308 28358
rect 13268 28144 13320 28150
rect 13268 28086 13320 28092
rect 12716 28076 12768 28082
rect 12716 28018 12768 28024
rect 13280 27674 13308 28086
rect 13268 27668 13320 27674
rect 13268 27610 13320 27616
rect 13268 26988 13320 26994
rect 13268 26930 13320 26936
rect 13176 26784 13228 26790
rect 13176 26726 13228 26732
rect 13188 25974 13216 26726
rect 13280 26586 13308 26930
rect 13268 26580 13320 26586
rect 13268 26522 13320 26528
rect 13556 26382 13584 28630
rect 13544 26376 13596 26382
rect 13544 26318 13596 26324
rect 13176 25968 13228 25974
rect 13176 25910 13228 25916
rect 13176 25832 13228 25838
rect 13176 25774 13228 25780
rect 13188 25294 13216 25774
rect 13176 25288 13228 25294
rect 13176 25230 13228 25236
rect 13556 25226 13584 26318
rect 13544 25220 13596 25226
rect 13544 25162 13596 25168
rect 12440 23520 12492 23526
rect 12440 23462 12492 23468
rect 12348 23044 12400 23050
rect 12348 22986 12400 22992
rect 12360 22778 12388 22986
rect 12348 22772 12400 22778
rect 12348 22714 12400 22720
rect 12256 22636 12308 22642
rect 12256 22578 12308 22584
rect 12268 22522 12296 22578
rect 12268 22494 12388 22522
rect 12176 22066 12296 22094
rect 12164 22024 12216 22030
rect 12164 21966 12216 21972
rect 11888 21616 11940 21622
rect 11888 21558 11940 21564
rect 11888 21480 11940 21486
rect 11888 21422 11940 21428
rect 10968 21412 11020 21418
rect 10968 21354 11020 21360
rect 10980 21146 11008 21354
rect 10968 21140 11020 21146
rect 10968 21082 11020 21088
rect 10980 20534 11008 21082
rect 10968 20528 11020 20534
rect 10968 20470 11020 20476
rect 11704 20392 11756 20398
rect 11704 20334 11756 20340
rect 11716 19786 11744 20334
rect 11900 20330 11928 21422
rect 12176 20398 12204 21966
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 11888 20324 11940 20330
rect 11888 20266 11940 20272
rect 11704 19780 11756 19786
rect 11704 19722 11756 19728
rect 11428 18828 11480 18834
rect 11428 18770 11480 18776
rect 11440 18358 11468 18770
rect 11428 18352 11480 18358
rect 11428 18294 11480 18300
rect 11440 17882 11468 18294
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11716 17134 11744 19722
rect 11704 17128 11756 17134
rect 11704 17070 11756 17076
rect 10876 16720 10928 16726
rect 10876 16662 10928 16668
rect 11716 16658 11744 17070
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11900 16590 11928 20266
rect 12268 19174 12296 22066
rect 12360 19446 12388 22494
rect 12452 21690 12480 23462
rect 12440 21684 12492 21690
rect 12440 21626 12492 21632
rect 13648 21418 13676 29106
rect 13728 28076 13780 28082
rect 13728 28018 13780 28024
rect 13740 27441 13768 28018
rect 13832 27606 13860 29990
rect 13924 29646 13952 30194
rect 13912 29640 13964 29646
rect 13912 29582 13964 29588
rect 14004 28756 14056 28762
rect 14004 28698 14056 28704
rect 14016 27674 14044 28698
rect 14004 27668 14056 27674
rect 14004 27610 14056 27616
rect 13820 27600 13872 27606
rect 13820 27542 13872 27548
rect 13726 27432 13782 27441
rect 13726 27367 13782 27376
rect 13740 25362 13768 27367
rect 13728 25356 13780 25362
rect 13728 25298 13780 25304
rect 14108 22094 14136 33102
rect 14188 32768 14240 32774
rect 14188 32710 14240 32716
rect 14200 32502 14228 32710
rect 14384 32570 14412 33390
rect 14372 32564 14424 32570
rect 14372 32506 14424 32512
rect 14188 32496 14240 32502
rect 14188 32438 14240 32444
rect 14556 32428 14608 32434
rect 14556 32370 14608 32376
rect 14372 32360 14424 32366
rect 14370 32328 14372 32337
rect 14424 32328 14426 32337
rect 14370 32263 14426 32272
rect 14188 32224 14240 32230
rect 14188 32166 14240 32172
rect 14200 30938 14228 32166
rect 14568 31754 14596 32370
rect 14556 31748 14608 31754
rect 14556 31690 14608 31696
rect 14556 31340 14608 31346
rect 14556 31282 14608 31288
rect 14188 30932 14240 30938
rect 14188 30874 14240 30880
rect 14200 30326 14228 30874
rect 14464 30388 14516 30394
rect 14464 30330 14516 30336
rect 14188 30320 14240 30326
rect 14188 30262 14240 30268
rect 14476 30258 14504 30330
rect 14568 30297 14596 31282
rect 14554 30288 14610 30297
rect 14464 30252 14516 30258
rect 14554 30223 14610 30232
rect 14464 30194 14516 30200
rect 14660 30122 14688 33390
rect 14648 30116 14700 30122
rect 14648 30058 14700 30064
rect 14464 29776 14516 29782
rect 14464 29718 14516 29724
rect 14280 29708 14332 29714
rect 14280 29650 14332 29656
rect 14188 29096 14240 29102
rect 14188 29038 14240 29044
rect 14200 27470 14228 29038
rect 14292 28558 14320 29650
rect 14372 28620 14424 28626
rect 14372 28562 14424 28568
rect 14280 28552 14332 28558
rect 14280 28494 14332 28500
rect 14188 27464 14240 27470
rect 14188 27406 14240 27412
rect 14200 25294 14228 27406
rect 14292 26926 14320 28494
rect 14384 28082 14412 28562
rect 14476 28558 14504 29718
rect 14648 29028 14700 29034
rect 14648 28970 14700 28976
rect 14660 28558 14688 28970
rect 14464 28552 14516 28558
rect 14464 28494 14516 28500
rect 14648 28552 14700 28558
rect 14648 28494 14700 28500
rect 14372 28076 14424 28082
rect 14372 28018 14424 28024
rect 14556 27872 14608 27878
rect 14556 27814 14608 27820
rect 14568 27470 14596 27814
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 14464 26988 14516 26994
rect 14464 26930 14516 26936
rect 14280 26920 14332 26926
rect 14280 26862 14332 26868
rect 14188 25288 14240 25294
rect 14188 25230 14240 25236
rect 14200 24732 14228 25230
rect 14280 24744 14332 24750
rect 14200 24704 14280 24732
rect 14280 24686 14332 24692
rect 14292 24206 14320 24686
rect 14372 24608 14424 24614
rect 14372 24550 14424 24556
rect 14384 24206 14412 24550
rect 14280 24200 14332 24206
rect 14280 24142 14332 24148
rect 14372 24200 14424 24206
rect 14372 24142 14424 24148
rect 14292 23186 14320 24142
rect 14476 23730 14504 26930
rect 14648 26920 14700 26926
rect 14648 26862 14700 26868
rect 14660 26382 14688 26862
rect 14648 26376 14700 26382
rect 14648 26318 14700 26324
rect 14660 25294 14688 26318
rect 14648 25288 14700 25294
rect 14648 25230 14700 25236
rect 14464 23724 14516 23730
rect 14464 23666 14516 23672
rect 14280 23180 14332 23186
rect 14280 23122 14332 23128
rect 14280 22704 14332 22710
rect 14280 22646 14332 22652
rect 14016 22066 14136 22094
rect 13728 21888 13780 21894
rect 13728 21830 13780 21836
rect 13544 21412 13596 21418
rect 13544 21354 13596 21360
rect 13636 21412 13688 21418
rect 13636 21354 13688 21360
rect 13556 20942 13584 21354
rect 13544 20936 13596 20942
rect 13544 20878 13596 20884
rect 12348 19440 12400 19446
rect 12400 19388 12480 19394
rect 12348 19382 12480 19388
rect 12360 19366 12480 19382
rect 12360 19317 12388 19366
rect 12256 19168 12308 19174
rect 12256 19110 12308 19116
rect 12268 18426 12296 19110
rect 12452 18698 12480 19366
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 12440 18692 12492 18698
rect 12440 18634 12492 18640
rect 13084 18692 13136 18698
rect 13084 18634 13136 18640
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12728 17746 12756 18022
rect 12716 17740 12768 17746
rect 12716 17682 12768 17688
rect 13096 17678 13124 18634
rect 13372 18154 13400 18702
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13464 18290 13492 18566
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 13360 18148 13412 18154
rect 13360 18090 13412 18096
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 12360 17270 12388 17478
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 13096 17066 13124 17478
rect 13084 17060 13136 17066
rect 13084 17002 13136 17008
rect 13544 17060 13596 17066
rect 13544 17002 13596 17008
rect 13096 16726 13124 17002
rect 13084 16720 13136 16726
rect 13084 16662 13136 16668
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 10692 16516 10744 16522
rect 10692 16458 10744 16464
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 12084 16182 12112 16390
rect 12072 16176 12124 16182
rect 12072 16118 12124 16124
rect 12164 16040 12216 16046
rect 12164 15982 12216 15988
rect 11152 15632 11204 15638
rect 11152 15574 11204 15580
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 10140 15020 10192 15026
rect 10520 15014 10640 15042
rect 11164 15026 11192 15574
rect 12176 15502 12204 15982
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 10140 14962 10192 14968
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8392 14816 8444 14822
rect 8392 14758 8444 14764
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7944 13938 7972 14418
rect 8404 14006 8432 14758
rect 9324 14074 9352 14962
rect 10612 14958 10640 15014
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 8392 14000 8444 14006
rect 8392 13942 8444 13948
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 7944 12986 7972 13874
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 7944 11694 7972 12922
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9232 12306 9260 12582
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9324 11898 9352 12174
rect 9784 11898 9812 12718
rect 10612 12442 10640 13874
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10704 13530 10732 13806
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10796 13326 10824 13466
rect 11164 13394 11192 14758
rect 11900 14414 11928 14962
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 11900 13938 11928 14350
rect 12084 14006 12112 14350
rect 12072 14000 12124 14006
rect 12072 13942 12124 13948
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 10784 13320 10836 13326
rect 10704 13280 10784 13308
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 7944 10130 7972 11630
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10336 11150 10364 11494
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10520 11014 10548 11630
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10704 10266 10732 13280
rect 10784 13262 10836 13268
rect 11164 12918 11192 13330
rect 12176 12918 12204 15438
rect 12452 14482 12480 16526
rect 13556 16522 13584 17002
rect 13648 16590 13676 21354
rect 13740 21078 13768 21830
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13728 21072 13780 21078
rect 13728 21014 13780 21020
rect 13832 20058 13860 21490
rect 13912 20868 13964 20874
rect 13912 20810 13964 20816
rect 13924 20602 13952 20810
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 14016 20262 14044 22066
rect 14292 21350 14320 22646
rect 14372 22636 14424 22642
rect 14372 22578 14424 22584
rect 14556 22636 14608 22642
rect 14556 22578 14608 22584
rect 14384 22234 14412 22578
rect 14464 22432 14516 22438
rect 14464 22374 14516 22380
rect 14372 22228 14424 22234
rect 14372 22170 14424 22176
rect 14476 22030 14504 22374
rect 14464 22024 14516 22030
rect 14464 21966 14516 21972
rect 14568 21570 14596 22578
rect 14648 21956 14700 21962
rect 14648 21898 14700 21904
rect 14476 21542 14596 21570
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 14476 20874 14504 21542
rect 14556 21480 14608 21486
rect 14556 21422 14608 21428
rect 14568 21146 14596 21422
rect 14556 21140 14608 21146
rect 14556 21082 14608 21088
rect 14464 20868 14516 20874
rect 14464 20810 14516 20816
rect 14280 20800 14332 20806
rect 14280 20742 14332 20748
rect 14292 20534 14320 20742
rect 14280 20528 14332 20534
rect 14280 20470 14332 20476
rect 14464 20460 14516 20466
rect 14464 20402 14516 20408
rect 14476 20262 14504 20402
rect 14556 20392 14608 20398
rect 14556 20334 14608 20340
rect 14004 20256 14056 20262
rect 14004 20198 14056 20204
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14568 20058 14596 20334
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 14280 18624 14332 18630
rect 14280 18566 14332 18572
rect 14292 18426 14320 18566
rect 14280 18420 14332 18426
rect 14280 18362 14332 18368
rect 14004 18080 14056 18086
rect 14004 18022 14056 18028
rect 14016 17746 14044 18022
rect 14004 17740 14056 17746
rect 14004 17682 14056 17688
rect 13820 17604 13872 17610
rect 13820 17546 13872 17552
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13544 16516 13596 16522
rect 13544 16458 13596 16464
rect 13556 16250 13584 16458
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 12532 14884 12584 14890
rect 12532 14826 12584 14832
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12452 13326 12480 14418
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12544 13172 12572 14826
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 12992 14340 13044 14346
rect 12992 14282 13044 14288
rect 13004 13938 13032 14282
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 13188 13870 13216 14350
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 12452 13144 12572 13172
rect 11152 12912 11204 12918
rect 11152 12854 11204 12860
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 11796 12368 11848 12374
rect 11796 12310 11848 12316
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10796 11354 10824 11698
rect 11072 11354 11100 11766
rect 11704 11620 11756 11626
rect 11704 11562 11756 11568
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11256 11150 11284 11494
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 10888 9178 10916 9998
rect 11072 9450 11100 11086
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11256 10062 11284 10406
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11256 9518 11284 9998
rect 11428 9988 11480 9994
rect 11428 9930 11480 9936
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 11348 9518 11376 9862
rect 11440 9586 11468 9930
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 11072 9042 11100 9386
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 11348 8974 11376 9454
rect 11716 9450 11744 11562
rect 11808 10674 11836 12310
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12360 11830 12388 12174
rect 12452 12170 12480 13144
rect 12728 12850 12756 13806
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 12912 12918 12940 13194
rect 12900 12912 12952 12918
rect 12900 12854 12952 12860
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12728 12714 12756 12786
rect 12716 12708 12768 12714
rect 12716 12650 12768 12656
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11992 10674 12020 11494
rect 12360 11150 12388 11766
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12452 11014 12480 12106
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 12544 10266 12572 12582
rect 12912 12434 12940 12854
rect 13188 12442 13216 13806
rect 13280 13190 13308 13874
rect 13268 13184 13320 13190
rect 13268 13126 13320 13132
rect 13280 12918 13308 13126
rect 13372 12986 13400 14962
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 13464 14618 13492 14894
rect 13544 14884 13596 14890
rect 13544 14826 13596 14832
rect 13452 14612 13504 14618
rect 13452 14554 13504 14560
rect 13556 13938 13584 14826
rect 13636 14000 13688 14006
rect 13636 13942 13688 13948
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13268 12912 13320 12918
rect 13268 12854 13320 12860
rect 13452 12912 13504 12918
rect 13452 12854 13504 12860
rect 13464 12714 13492 12854
rect 13648 12714 13676 13942
rect 13832 13818 13860 17546
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 14200 16114 14228 16594
rect 14188 16108 14240 16114
rect 14188 16050 14240 16056
rect 14464 16040 14516 16046
rect 14464 15982 14516 15988
rect 14476 15162 14504 15982
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 14660 14414 14688 21898
rect 14752 21350 14780 33816
rect 15476 33798 15528 33804
rect 15016 33516 15068 33522
rect 15016 33458 15068 33464
rect 15384 33516 15436 33522
rect 15384 33458 15436 33464
rect 14832 33312 14884 33318
rect 14832 33254 14884 33260
rect 14844 32366 14872 33254
rect 14924 32428 14976 32434
rect 14924 32370 14976 32376
rect 14832 32360 14884 32366
rect 14832 32302 14884 32308
rect 14936 32026 14964 32370
rect 14924 32020 14976 32026
rect 14924 31962 14976 31968
rect 14832 31816 14884 31822
rect 14832 31758 14884 31764
rect 14844 28762 14872 31758
rect 15028 31686 15056 33458
rect 15200 33380 15252 33386
rect 15200 33322 15252 33328
rect 15108 32904 15160 32910
rect 15108 32846 15160 32852
rect 15120 32026 15148 32846
rect 15212 32842 15240 33322
rect 15396 33130 15424 33458
rect 15488 33318 15516 33798
rect 15856 33386 15884 33934
rect 15844 33380 15896 33386
rect 15844 33322 15896 33328
rect 15476 33312 15528 33318
rect 15476 33254 15528 33260
rect 15396 33102 15516 33130
rect 15856 33114 15884 33322
rect 15948 33114 15976 34954
rect 16040 34678 16068 37130
rect 16488 36780 16540 36786
rect 16488 36722 16540 36728
rect 16500 36242 16528 36722
rect 18052 36712 18104 36718
rect 18052 36654 18104 36660
rect 17684 36644 17736 36650
rect 17684 36586 17736 36592
rect 16948 36576 17000 36582
rect 16948 36518 17000 36524
rect 16488 36236 16540 36242
rect 16488 36178 16540 36184
rect 16212 36168 16264 36174
rect 16212 36110 16264 36116
rect 16120 36032 16172 36038
rect 16120 35974 16172 35980
rect 16028 34672 16080 34678
rect 16028 34614 16080 34620
rect 16040 34105 16068 34614
rect 16026 34096 16082 34105
rect 16026 34031 16082 34040
rect 15384 32972 15436 32978
rect 15384 32914 15436 32920
rect 15200 32836 15252 32842
rect 15200 32778 15252 32784
rect 15396 32366 15424 32914
rect 15488 32366 15516 33102
rect 15660 33108 15712 33114
rect 15660 33050 15712 33056
rect 15844 33108 15896 33114
rect 15844 33050 15896 33056
rect 15936 33108 15988 33114
rect 15936 33050 15988 33056
rect 15672 32774 15700 33050
rect 15660 32768 15712 32774
rect 15660 32710 15712 32716
rect 15384 32360 15436 32366
rect 15384 32302 15436 32308
rect 15476 32360 15528 32366
rect 15476 32302 15528 32308
rect 15108 32020 15160 32026
rect 15108 31962 15160 31968
rect 15200 32020 15252 32026
rect 15200 31962 15252 31968
rect 15016 31680 15068 31686
rect 15016 31622 15068 31628
rect 15016 30932 15068 30938
rect 15016 30874 15068 30880
rect 15028 30734 15056 30874
rect 15016 30728 15068 30734
rect 15212 30682 15240 31962
rect 15396 31482 15424 32302
rect 15488 32230 15516 32302
rect 15476 32224 15528 32230
rect 15476 32166 15528 32172
rect 15752 31816 15804 31822
rect 15752 31758 15804 31764
rect 15384 31476 15436 31482
rect 15384 31418 15436 31424
rect 15384 31272 15436 31278
rect 15384 31214 15436 31220
rect 15476 31272 15528 31278
rect 15476 31214 15528 31220
rect 15016 30670 15068 30676
rect 15120 30654 15240 30682
rect 15016 30592 15068 30598
rect 15016 30534 15068 30540
rect 14924 30048 14976 30054
rect 14924 29990 14976 29996
rect 14936 29102 14964 29990
rect 14924 29096 14976 29102
rect 14924 29038 14976 29044
rect 14832 28756 14884 28762
rect 14832 28698 14884 28704
rect 15028 28422 15056 30534
rect 15120 30138 15148 30654
rect 15200 30592 15252 30598
rect 15200 30534 15252 30540
rect 15212 30258 15240 30534
rect 15200 30252 15252 30258
rect 15200 30194 15252 30200
rect 15120 30110 15240 30138
rect 15212 28694 15240 30110
rect 15396 29714 15424 31214
rect 15488 30870 15516 31214
rect 15476 30864 15528 30870
rect 15476 30806 15528 30812
rect 15764 30818 15792 31758
rect 15844 31748 15896 31754
rect 15844 31690 15896 31696
rect 15856 31210 15884 31690
rect 15844 31204 15896 31210
rect 15844 31146 15896 31152
rect 15764 30790 15976 30818
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 15844 30728 15896 30734
rect 15844 30670 15896 30676
rect 15488 29850 15516 30670
rect 15752 30388 15804 30394
rect 15752 30330 15804 30336
rect 15764 30190 15792 30330
rect 15752 30184 15804 30190
rect 15752 30126 15804 30132
rect 15568 30048 15620 30054
rect 15568 29990 15620 29996
rect 15660 30048 15712 30054
rect 15660 29990 15712 29996
rect 15476 29844 15528 29850
rect 15476 29786 15528 29792
rect 15384 29708 15436 29714
rect 15384 29650 15436 29656
rect 15580 28762 15608 29990
rect 15672 29782 15700 29990
rect 15660 29776 15712 29782
rect 15660 29718 15712 29724
rect 15672 29306 15700 29718
rect 15752 29640 15804 29646
rect 15750 29608 15752 29617
rect 15804 29608 15806 29617
rect 15750 29543 15806 29552
rect 15660 29300 15712 29306
rect 15660 29242 15712 29248
rect 15856 28966 15884 30670
rect 15948 30054 15976 30790
rect 16028 30252 16080 30258
rect 16028 30194 16080 30200
rect 15936 30048 15988 30054
rect 15936 29990 15988 29996
rect 16040 29730 16068 30194
rect 15948 29702 16068 29730
rect 15948 29510 15976 29702
rect 16028 29572 16080 29578
rect 16028 29514 16080 29520
rect 15936 29504 15988 29510
rect 15936 29446 15988 29452
rect 15844 28960 15896 28966
rect 15844 28902 15896 28908
rect 15568 28756 15620 28762
rect 15568 28698 15620 28704
rect 15200 28688 15252 28694
rect 15200 28630 15252 28636
rect 15016 28416 15068 28422
rect 15016 28358 15068 28364
rect 15660 27940 15712 27946
rect 15660 27882 15712 27888
rect 15672 27606 15700 27882
rect 15660 27600 15712 27606
rect 15660 27542 15712 27548
rect 15568 26784 15620 26790
rect 15568 26726 15620 26732
rect 15580 26382 15608 26726
rect 15568 26376 15620 26382
rect 15568 26318 15620 26324
rect 15016 26308 15068 26314
rect 15016 26250 15068 26256
rect 15108 26308 15160 26314
rect 15108 26250 15160 26256
rect 14832 25152 14884 25158
rect 14832 25094 14884 25100
rect 14844 24818 14872 25094
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14924 21480 14976 21486
rect 14924 21422 14976 21428
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 14752 20602 14780 20742
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 14752 18358 14780 20334
rect 14936 19242 14964 21422
rect 14924 19236 14976 19242
rect 14924 19178 14976 19184
rect 14936 18766 14964 19178
rect 14924 18760 14976 18766
rect 14924 18702 14976 18708
rect 14740 18352 14792 18358
rect 14740 18294 14792 18300
rect 14924 17604 14976 17610
rect 14924 17546 14976 17552
rect 14936 17338 14964 17546
rect 14924 17332 14976 17338
rect 14924 17274 14976 17280
rect 15028 17218 15056 26250
rect 15120 26042 15148 26250
rect 15108 26036 15160 26042
rect 15108 25978 15160 25984
rect 15106 25528 15162 25537
rect 15672 25514 15700 27542
rect 16040 26382 16068 29514
rect 16028 26376 16080 26382
rect 16028 26318 16080 26324
rect 15106 25463 15162 25472
rect 15580 25486 15700 25514
rect 15120 22642 15148 25463
rect 15580 24750 15608 25486
rect 15660 25220 15712 25226
rect 15660 25162 15712 25168
rect 15568 24744 15620 24750
rect 15568 24686 15620 24692
rect 15200 23248 15252 23254
rect 15200 23190 15252 23196
rect 15108 22636 15160 22642
rect 15108 22578 15160 22584
rect 15212 22098 15240 23190
rect 15384 23112 15436 23118
rect 15384 23054 15436 23060
rect 15292 22704 15344 22710
rect 15292 22646 15344 22652
rect 15304 22506 15332 22646
rect 15292 22500 15344 22506
rect 15292 22442 15344 22448
rect 15396 22098 15424 23054
rect 15476 22432 15528 22438
rect 15476 22374 15528 22380
rect 15200 22092 15252 22098
rect 15200 22034 15252 22040
rect 15384 22092 15436 22098
rect 15384 22034 15436 22040
rect 15488 22030 15516 22374
rect 15476 22024 15528 22030
rect 15476 21966 15528 21972
rect 15200 21344 15252 21350
rect 15200 21286 15252 21292
rect 15384 21344 15436 21350
rect 15384 21286 15436 21292
rect 15212 20806 15240 21286
rect 15292 21004 15344 21010
rect 15292 20946 15344 20952
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 15304 20534 15332 20946
rect 15396 20534 15424 21286
rect 15580 20942 15608 24686
rect 15672 24614 15700 25162
rect 15660 24608 15712 24614
rect 15660 24550 15712 24556
rect 15672 23322 15700 24550
rect 16040 23798 16068 26318
rect 15844 23792 15896 23798
rect 15844 23734 15896 23740
rect 16028 23792 16080 23798
rect 16028 23734 16080 23740
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15752 23112 15804 23118
rect 15752 23054 15804 23060
rect 15672 22778 15700 23054
rect 15660 22772 15712 22778
rect 15660 22714 15712 22720
rect 15764 21622 15792 23054
rect 15752 21616 15804 21622
rect 15752 21558 15804 21564
rect 15660 21548 15712 21554
rect 15660 21490 15712 21496
rect 15672 21298 15700 21490
rect 15856 21434 15884 23734
rect 16028 22976 16080 22982
rect 16028 22918 16080 22924
rect 16040 22706 16068 22918
rect 16132 22760 16160 35974
rect 16224 33658 16252 36110
rect 16500 35698 16528 36178
rect 16960 36106 16988 36518
rect 16948 36100 17000 36106
rect 16948 36042 17000 36048
rect 17696 35698 17724 36586
rect 16488 35692 16540 35698
rect 16488 35634 16540 35640
rect 17684 35692 17736 35698
rect 17684 35634 17736 35640
rect 17960 35624 18012 35630
rect 17960 35566 18012 35572
rect 16580 35488 16632 35494
rect 16580 35430 16632 35436
rect 16948 35488 17000 35494
rect 16948 35430 17000 35436
rect 16592 33930 16620 35430
rect 16960 35018 16988 35430
rect 16948 35012 17000 35018
rect 16948 34954 17000 34960
rect 17972 34542 18000 35566
rect 17408 34536 17460 34542
rect 17408 34478 17460 34484
rect 17960 34536 18012 34542
rect 17960 34478 18012 34484
rect 16580 33924 16632 33930
rect 16580 33866 16632 33872
rect 16212 33652 16264 33658
rect 16212 33594 16264 33600
rect 17420 33522 17448 34478
rect 17960 34400 18012 34406
rect 17960 34342 18012 34348
rect 17684 34060 17736 34066
rect 17684 34002 17736 34008
rect 17592 33856 17644 33862
rect 17592 33798 17644 33804
rect 17500 33652 17552 33658
rect 17500 33594 17552 33600
rect 17408 33516 17460 33522
rect 17408 33458 17460 33464
rect 16948 33448 17000 33454
rect 16948 33390 17000 33396
rect 16304 32564 16356 32570
rect 16304 32506 16356 32512
rect 16316 32434 16344 32506
rect 16856 32496 16908 32502
rect 16856 32438 16908 32444
rect 16304 32428 16356 32434
rect 16304 32370 16356 32376
rect 16212 32224 16264 32230
rect 16212 32166 16264 32172
rect 16224 31346 16252 32166
rect 16316 31754 16344 32370
rect 16316 31726 16436 31754
rect 16212 31340 16264 31346
rect 16212 31282 16264 31288
rect 16304 30116 16356 30122
rect 16304 30058 16356 30064
rect 16212 29504 16264 29510
rect 16212 29446 16264 29452
rect 16224 29238 16252 29446
rect 16212 29232 16264 29238
rect 16212 29174 16264 29180
rect 16224 28490 16252 29174
rect 16316 29102 16344 30058
rect 16304 29096 16356 29102
rect 16304 29038 16356 29044
rect 16304 28960 16356 28966
rect 16304 28902 16356 28908
rect 16316 28558 16344 28902
rect 16304 28552 16356 28558
rect 16304 28494 16356 28500
rect 16212 28484 16264 28490
rect 16212 28426 16264 28432
rect 16408 26994 16436 31726
rect 16868 31414 16896 32438
rect 16960 32230 16988 33390
rect 17512 33386 17540 33594
rect 17500 33380 17552 33386
rect 17500 33322 17552 33328
rect 17604 32910 17632 33798
rect 17592 32904 17644 32910
rect 17592 32846 17644 32852
rect 17316 32428 17368 32434
rect 17316 32370 17368 32376
rect 16948 32224 17000 32230
rect 16948 32166 17000 32172
rect 17224 31952 17276 31958
rect 17224 31894 17276 31900
rect 16948 31816 17000 31822
rect 16948 31758 17000 31764
rect 16960 31414 16988 31758
rect 16856 31408 16908 31414
rect 16856 31350 16908 31356
rect 16948 31408 17000 31414
rect 16948 31350 17000 31356
rect 17236 31278 17264 31894
rect 17328 31822 17356 32370
rect 17604 32337 17632 32846
rect 17696 32434 17724 34002
rect 17972 33930 18000 34342
rect 17960 33924 18012 33930
rect 17960 33866 18012 33872
rect 17776 33448 17828 33454
rect 17972 33436 18000 33866
rect 17828 33408 18000 33436
rect 17776 33390 17828 33396
rect 17776 32972 17828 32978
rect 17776 32914 17828 32920
rect 17684 32428 17736 32434
rect 17684 32370 17736 32376
rect 17590 32328 17646 32337
rect 17590 32263 17646 32272
rect 17408 32224 17460 32230
rect 17406 32192 17408 32201
rect 17500 32224 17552 32230
rect 17460 32192 17462 32201
rect 17500 32166 17552 32172
rect 17682 32192 17738 32201
rect 17406 32127 17462 32136
rect 17408 32020 17460 32026
rect 17408 31962 17460 31968
rect 17316 31816 17368 31822
rect 17314 31784 17316 31793
rect 17368 31784 17370 31793
rect 17314 31719 17370 31728
rect 17420 31482 17448 31962
rect 17512 31890 17540 32166
rect 17682 32127 17738 32136
rect 17500 31884 17552 31890
rect 17500 31826 17552 31832
rect 17408 31476 17460 31482
rect 17408 31418 17460 31424
rect 17224 31272 17276 31278
rect 17224 31214 17276 31220
rect 17408 31272 17460 31278
rect 17408 31214 17460 31220
rect 16580 30728 16632 30734
rect 16580 30670 16632 30676
rect 17224 30728 17276 30734
rect 17224 30670 17276 30676
rect 16592 30394 16620 30670
rect 16580 30388 16632 30394
rect 16580 30330 16632 30336
rect 16488 29640 16540 29646
rect 16592 29628 16620 30330
rect 16856 30116 16908 30122
rect 16856 30058 16908 30064
rect 16868 29646 16896 30058
rect 16540 29600 16620 29628
rect 16856 29640 16908 29646
rect 16670 29608 16726 29617
rect 16488 29582 16540 29588
rect 16856 29582 16908 29588
rect 16670 29543 16726 29552
rect 16488 29096 16540 29102
rect 16488 29038 16540 29044
rect 16396 26988 16448 26994
rect 16396 26930 16448 26936
rect 16500 23526 16528 29038
rect 16580 27124 16632 27130
rect 16580 27066 16632 27072
rect 16592 25430 16620 27066
rect 16684 26586 16712 29543
rect 16764 29504 16816 29510
rect 16764 29446 16816 29452
rect 16776 28694 16804 29446
rect 16868 28762 16896 29582
rect 16948 29164 17000 29170
rect 16948 29106 17000 29112
rect 16856 28756 16908 28762
rect 16856 28698 16908 28704
rect 16764 28688 16816 28694
rect 16764 28630 16816 28636
rect 16764 28552 16816 28558
rect 16764 28494 16816 28500
rect 16776 28150 16804 28494
rect 16960 28218 16988 29106
rect 17040 28484 17092 28490
rect 17040 28426 17092 28432
rect 16948 28212 17000 28218
rect 16948 28154 17000 28160
rect 16764 28144 16816 28150
rect 16764 28086 16816 28092
rect 17052 28082 17080 28426
rect 17040 28076 17092 28082
rect 17040 28018 17092 28024
rect 17040 27600 17092 27606
rect 17040 27542 17092 27548
rect 17052 26994 17080 27542
rect 17040 26988 17092 26994
rect 16960 26948 17040 26976
rect 16672 26580 16724 26586
rect 16672 26522 16724 26528
rect 16960 26382 16988 26948
rect 17040 26930 17092 26936
rect 17236 26926 17264 30670
rect 17420 30054 17448 31214
rect 17592 31204 17644 31210
rect 17592 31146 17644 31152
rect 17500 31136 17552 31142
rect 17500 31078 17552 31084
rect 17512 30666 17540 31078
rect 17604 30666 17632 31146
rect 17500 30660 17552 30666
rect 17500 30602 17552 30608
rect 17592 30660 17644 30666
rect 17592 30602 17644 30608
rect 17512 30190 17540 30602
rect 17500 30184 17552 30190
rect 17500 30126 17552 30132
rect 17408 30048 17460 30054
rect 17408 29990 17460 29996
rect 17316 29572 17368 29578
rect 17316 29514 17368 29520
rect 17328 28762 17356 29514
rect 17408 29096 17460 29102
rect 17406 29064 17408 29073
rect 17460 29064 17462 29073
rect 17406 28999 17462 29008
rect 17316 28756 17368 28762
rect 17316 28698 17368 28704
rect 17604 28218 17632 30602
rect 17696 30122 17724 32127
rect 17684 30116 17736 30122
rect 17684 30058 17736 30064
rect 17788 29850 17816 32914
rect 17868 32904 17920 32910
rect 17868 32846 17920 32852
rect 17880 30682 17908 32846
rect 17972 31822 18000 33408
rect 18064 33114 18092 36654
rect 18420 36168 18472 36174
rect 18420 36110 18472 36116
rect 18236 36100 18288 36106
rect 18236 36042 18288 36048
rect 18248 35086 18276 36042
rect 18432 35562 18460 36110
rect 18420 35556 18472 35562
rect 18420 35498 18472 35504
rect 18432 35290 18460 35498
rect 18420 35284 18472 35290
rect 18420 35226 18472 35232
rect 18236 35080 18288 35086
rect 18236 35022 18288 35028
rect 18248 34610 18276 35022
rect 18420 35012 18472 35018
rect 18420 34954 18472 34960
rect 18236 34604 18288 34610
rect 18236 34546 18288 34552
rect 18248 34406 18276 34546
rect 18432 34474 18460 34954
rect 18420 34468 18472 34474
rect 18420 34410 18472 34416
rect 18144 34400 18196 34406
rect 18144 34342 18196 34348
rect 18236 34400 18288 34406
rect 18236 34342 18288 34348
rect 18156 33114 18184 34342
rect 18248 33522 18276 34342
rect 18616 34134 18644 37130
rect 22468 37120 22520 37126
rect 22468 37062 22520 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19524 36780 19576 36786
rect 19524 36722 19576 36728
rect 19984 36780 20036 36786
rect 19984 36722 20036 36728
rect 22100 36780 22152 36786
rect 22100 36722 22152 36728
rect 19536 36378 19564 36722
rect 19892 36576 19944 36582
rect 19892 36518 19944 36524
rect 19524 36372 19576 36378
rect 19524 36314 19576 36320
rect 19904 36174 19932 36518
rect 19892 36168 19944 36174
rect 19892 36110 19944 36116
rect 18788 36032 18840 36038
rect 18788 35974 18840 35980
rect 18800 35698 18828 35974
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 18788 35692 18840 35698
rect 18788 35634 18840 35640
rect 19892 35692 19944 35698
rect 19996 35680 20024 36722
rect 20812 36712 20864 36718
rect 20812 36654 20864 36660
rect 20076 36644 20128 36650
rect 20076 36586 20128 36592
rect 19944 35652 20024 35680
rect 19892 35634 19944 35640
rect 19156 35624 19208 35630
rect 20088 35578 20116 36586
rect 20628 36236 20680 36242
rect 20628 36178 20680 36184
rect 20444 36168 20496 36174
rect 20444 36110 20496 36116
rect 20456 35698 20484 36110
rect 20640 35766 20668 36178
rect 20824 36106 20852 36654
rect 20812 36100 20864 36106
rect 20812 36042 20864 36048
rect 20996 36100 21048 36106
rect 20996 36042 21048 36048
rect 20628 35760 20680 35766
rect 20628 35702 20680 35708
rect 20444 35692 20496 35698
rect 20444 35634 20496 35640
rect 19156 35566 19208 35572
rect 19064 35012 19116 35018
rect 19064 34954 19116 34960
rect 19076 34542 19104 34954
rect 19168 34950 19196 35566
rect 19708 35556 19760 35562
rect 19708 35498 19760 35504
rect 19812 35550 20392 35578
rect 19340 35216 19392 35222
rect 19340 35158 19392 35164
rect 19156 34944 19208 34950
rect 19156 34886 19208 34892
rect 19168 34746 19196 34886
rect 19156 34740 19208 34746
rect 19156 34682 19208 34688
rect 19064 34536 19116 34542
rect 19064 34478 19116 34484
rect 18604 34128 18656 34134
rect 18604 34070 18656 34076
rect 19076 33930 19104 34478
rect 19064 33924 19116 33930
rect 19064 33866 19116 33872
rect 18236 33516 18288 33522
rect 18236 33458 18288 33464
rect 18052 33108 18104 33114
rect 18052 33050 18104 33056
rect 18144 33108 18196 33114
rect 18144 33050 18196 33056
rect 18144 32836 18196 32842
rect 18144 32778 18196 32784
rect 18156 32434 18184 32778
rect 18144 32428 18196 32434
rect 18144 32370 18196 32376
rect 17960 31816 18012 31822
rect 17960 31758 18012 31764
rect 17880 30654 18000 30682
rect 17868 30592 17920 30598
rect 17868 30534 17920 30540
rect 17776 29844 17828 29850
rect 17776 29786 17828 29792
rect 17776 29640 17828 29646
rect 17880 29628 17908 30534
rect 17972 30190 18000 30654
rect 18052 30592 18104 30598
rect 18052 30534 18104 30540
rect 18144 30592 18196 30598
rect 18144 30534 18196 30540
rect 18064 30258 18092 30534
rect 18156 30326 18184 30534
rect 18144 30320 18196 30326
rect 18144 30262 18196 30268
rect 18052 30252 18104 30258
rect 18052 30194 18104 30200
rect 17960 30184 18012 30190
rect 18248 30172 18276 33458
rect 18328 33108 18380 33114
rect 18328 33050 18380 33056
rect 17960 30126 18012 30132
rect 18156 30144 18276 30172
rect 17828 29600 17908 29628
rect 17776 29582 17828 29588
rect 17684 28688 17736 28694
rect 17684 28630 17736 28636
rect 17592 28212 17644 28218
rect 17592 28154 17644 28160
rect 17696 27470 17724 28630
rect 17684 27464 17736 27470
rect 17684 27406 17736 27412
rect 17696 26994 17724 27406
rect 17316 26988 17368 26994
rect 17316 26930 17368 26936
rect 17684 26988 17736 26994
rect 17684 26930 17736 26936
rect 17224 26920 17276 26926
rect 17224 26862 17276 26868
rect 17132 26852 17184 26858
rect 17132 26794 17184 26800
rect 17144 26382 17172 26794
rect 17236 26382 17264 26862
rect 17328 26518 17356 26930
rect 17500 26852 17552 26858
rect 17500 26794 17552 26800
rect 17316 26512 17368 26518
rect 17316 26454 17368 26460
rect 16948 26376 17000 26382
rect 16948 26318 17000 26324
rect 17132 26376 17184 26382
rect 17132 26318 17184 26324
rect 17224 26376 17276 26382
rect 17224 26318 17276 26324
rect 16960 26042 16988 26318
rect 16948 26036 17000 26042
rect 16948 25978 17000 25984
rect 17144 25922 17172 26318
rect 17052 25906 17172 25922
rect 17040 25900 17172 25906
rect 17092 25894 17172 25900
rect 17040 25842 17092 25848
rect 17224 25696 17276 25702
rect 17224 25638 17276 25644
rect 16580 25424 16632 25430
rect 16580 25366 16632 25372
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 16764 24608 16816 24614
rect 16764 24550 16816 24556
rect 16776 24274 16804 24550
rect 16764 24268 16816 24274
rect 16764 24210 16816 24216
rect 16868 23866 16896 24754
rect 17236 24274 17264 25638
rect 17316 25152 17368 25158
rect 17316 25094 17368 25100
rect 17224 24268 17276 24274
rect 17224 24210 17276 24216
rect 17328 24206 17356 25094
rect 17316 24200 17368 24206
rect 17316 24142 17368 24148
rect 16856 23860 16908 23866
rect 16856 23802 16908 23808
rect 16304 23520 16356 23526
rect 16304 23462 16356 23468
rect 16488 23520 16540 23526
rect 16488 23462 16540 23468
rect 16132 22732 16252 22760
rect 16040 22642 16069 22706
rect 16029 22636 16081 22642
rect 16029 22578 16081 22584
rect 15936 22160 15988 22166
rect 15936 22102 15988 22108
rect 15948 21962 15976 22102
rect 15936 21956 15988 21962
rect 15936 21898 15988 21904
rect 15948 21706 15976 21898
rect 16040 21894 16068 22578
rect 16224 22506 16252 22732
rect 16212 22500 16264 22506
rect 16212 22442 16264 22448
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 16028 21888 16080 21894
rect 16028 21830 16080 21836
rect 15948 21678 16068 21706
rect 15856 21406 15976 21434
rect 15844 21344 15896 21350
rect 15672 21270 15792 21298
rect 15844 21286 15896 21292
rect 15568 20936 15620 20942
rect 15568 20878 15620 20884
rect 15764 20874 15792 21270
rect 15856 21146 15884 21286
rect 15844 21140 15896 21146
rect 15844 21082 15896 21088
rect 15948 20992 15976 21406
rect 15856 20964 15976 20992
rect 15752 20868 15804 20874
rect 15752 20810 15804 20816
rect 15660 20800 15712 20806
rect 15660 20742 15712 20748
rect 15292 20528 15344 20534
rect 15292 20470 15344 20476
rect 15384 20528 15436 20534
rect 15384 20470 15436 20476
rect 15672 20398 15700 20742
rect 15752 20528 15804 20534
rect 15752 20470 15804 20476
rect 15384 20392 15436 20398
rect 15384 20334 15436 20340
rect 15660 20392 15712 20398
rect 15764 20369 15792 20470
rect 15660 20334 15712 20340
rect 15750 20360 15806 20369
rect 15200 19780 15252 19786
rect 15200 19722 15252 19728
rect 15212 19394 15240 19722
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15304 19514 15332 19654
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15212 19366 15332 19394
rect 15200 18216 15252 18222
rect 15200 18158 15252 18164
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 15120 17678 15148 17818
rect 15212 17814 15240 18158
rect 15200 17808 15252 17814
rect 15200 17750 15252 17756
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 14936 17190 15056 17218
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 13740 13802 13860 13818
rect 13728 13796 13860 13802
rect 13780 13790 13860 13796
rect 13728 13738 13780 13744
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14568 12850 14596 13126
rect 14660 12986 14688 14350
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 13452 12708 13504 12714
rect 13452 12650 13504 12656
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13176 12436 13228 12442
rect 12912 12406 13032 12434
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 12636 11830 12664 12242
rect 12624 11824 12676 11830
rect 12624 11766 12676 11772
rect 12636 11150 12664 11766
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12452 9722 12480 9862
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12452 9602 12480 9658
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 12164 9580 12216 9586
rect 12452 9574 12572 9602
rect 12164 9522 12216 9528
rect 11704 9444 11756 9450
rect 11704 9386 11756 9392
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11808 8498 11836 9522
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 11808 8090 11836 8434
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11992 7342 12020 9318
rect 12176 9042 12204 9522
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 12452 8634 12480 9454
rect 12544 9042 12572 9574
rect 12912 9042 12940 10202
rect 13004 9518 13032 12406
rect 13176 12378 13228 12384
rect 13464 12238 13492 12650
rect 14016 12345 14044 12786
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14002 12336 14058 12345
rect 14200 12306 14228 12582
rect 14002 12271 14058 12280
rect 14188 12300 14240 12306
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13188 10062 13216 10610
rect 13280 10130 13308 12174
rect 14016 11150 14044 12271
rect 14188 12242 14240 12248
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13372 10674 13400 10950
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12728 7886 12756 8774
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12820 8090 12848 8434
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 11992 6866 12020 7278
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 12268 6798 12296 7822
rect 12900 7812 12952 7818
rect 12900 7754 12952 7760
rect 12912 7274 12940 7754
rect 13004 7410 13032 9454
rect 13372 7478 13400 10202
rect 13556 9042 13584 10406
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 14476 8974 14504 10066
rect 14752 9654 14780 16934
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14844 11354 14872 12718
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14832 10192 14884 10198
rect 14832 10134 14884 10140
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14660 8974 14688 9318
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 14476 8634 14504 8910
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14844 8498 14872 10134
rect 14936 9654 14964 17190
rect 15120 16998 15148 17614
rect 15212 17202 15240 17750
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 15198 15056 15254 15065
rect 15198 14991 15200 15000
rect 15252 14991 15254 15000
rect 15200 14962 15252 14968
rect 15212 14328 15240 14962
rect 15304 14822 15332 19366
rect 15396 18884 15424 20334
rect 15750 20295 15806 20304
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 15672 18970 15700 19314
rect 15660 18964 15712 18970
rect 15660 18906 15712 18912
rect 15476 18896 15528 18902
rect 15396 18856 15476 18884
rect 15396 18290 15424 18856
rect 15476 18838 15528 18844
rect 15384 18284 15436 18290
rect 15384 18226 15436 18232
rect 15764 18154 15792 19314
rect 15856 18902 15884 20964
rect 15936 20868 15988 20874
rect 15936 20810 15988 20816
rect 15948 19854 15976 20810
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15948 19310 15976 19790
rect 15936 19304 15988 19310
rect 15936 19246 15988 19252
rect 15844 18896 15896 18902
rect 15844 18838 15896 18844
rect 15856 18290 15884 18838
rect 15948 18358 15976 19246
rect 15936 18352 15988 18358
rect 15936 18294 15988 18300
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15752 18148 15804 18154
rect 15752 18090 15804 18096
rect 15476 17604 15528 17610
rect 15476 17546 15528 17552
rect 15488 17338 15516 17546
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15672 17202 15700 17478
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15568 17128 15620 17134
rect 15568 17070 15620 17076
rect 15384 17060 15436 17066
rect 15384 17002 15436 17008
rect 15396 16590 15424 17002
rect 15476 16720 15528 16726
rect 15476 16662 15528 16668
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 15384 14884 15436 14890
rect 15384 14826 15436 14832
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15292 14340 15344 14346
rect 15212 14300 15292 14328
rect 15292 14282 15344 14288
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 15028 13326 15056 13874
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15108 13796 15160 13802
rect 15108 13738 15160 13744
rect 15120 13530 15148 13738
rect 15212 13530 15240 13806
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 15028 12442 15056 13262
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 15304 11014 15332 14282
rect 15396 13938 15424 14826
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15396 13394 15424 13874
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15384 12368 15436 12374
rect 15384 12310 15436 12316
rect 15396 11694 15424 12310
rect 15488 12186 15516 16662
rect 15580 16590 15608 17070
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15764 16182 15792 18090
rect 15856 17202 15884 18226
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 15752 16176 15804 16182
rect 15752 16118 15804 16124
rect 16040 15502 16068 21678
rect 16224 21486 16252 21966
rect 16212 21480 16264 21486
rect 16212 21422 16264 21428
rect 16316 19786 16344 23462
rect 17224 23044 17276 23050
rect 17224 22986 17276 22992
rect 16856 22704 16908 22710
rect 17236 22681 17264 22986
rect 16856 22646 16908 22652
rect 17222 22672 17278 22681
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 16488 22568 16540 22574
rect 16488 22510 16540 22516
rect 16500 22234 16528 22510
rect 16488 22228 16540 22234
rect 16488 22170 16540 22176
rect 16500 20330 16528 22170
rect 16592 22098 16620 22578
rect 16868 22438 16896 22646
rect 17132 22636 17184 22642
rect 17512 22642 17540 26794
rect 17592 26580 17644 26586
rect 17592 26522 17644 26528
rect 17604 26382 17632 26522
rect 17592 26376 17644 26382
rect 17592 26318 17644 26324
rect 17604 24206 17632 26318
rect 17696 25906 17724 26930
rect 17684 25900 17736 25906
rect 17684 25842 17736 25848
rect 17684 25288 17736 25294
rect 17684 25230 17736 25236
rect 17696 24818 17724 25230
rect 17788 25158 17816 29582
rect 17868 29300 17920 29306
rect 17868 29242 17920 29248
rect 17880 28558 17908 29242
rect 18156 29170 18184 30144
rect 18236 30048 18288 30054
rect 18236 29990 18288 29996
rect 18248 29714 18276 29990
rect 18236 29708 18288 29714
rect 18236 29650 18288 29656
rect 18340 29578 18368 33050
rect 18420 32768 18472 32774
rect 18420 32710 18472 32716
rect 18696 32768 18748 32774
rect 18696 32710 18748 32716
rect 18432 32298 18460 32710
rect 18420 32292 18472 32298
rect 18420 32234 18472 32240
rect 18512 32224 18564 32230
rect 18512 32166 18564 32172
rect 18420 31816 18472 31822
rect 18420 31758 18472 31764
rect 18328 29572 18380 29578
rect 18328 29514 18380 29520
rect 18144 29164 18196 29170
rect 18144 29106 18196 29112
rect 18432 29084 18460 31758
rect 18524 31346 18552 32166
rect 18708 31822 18736 32710
rect 18788 32224 18840 32230
rect 18788 32166 18840 32172
rect 18800 31890 18828 32166
rect 19076 31958 19104 33866
rect 19168 33454 19196 34682
rect 19248 33992 19300 33998
rect 19248 33934 19300 33940
rect 19156 33448 19208 33454
rect 19156 33390 19208 33396
rect 19064 31952 19116 31958
rect 19064 31894 19116 31900
rect 18788 31884 18840 31890
rect 18972 31884 19024 31890
rect 18788 31826 18840 31832
rect 18892 31844 18972 31872
rect 18696 31816 18748 31822
rect 18696 31758 18748 31764
rect 18512 31340 18564 31346
rect 18512 31282 18564 31288
rect 18708 30802 18736 31758
rect 18892 31482 18920 31844
rect 18972 31826 19024 31832
rect 18972 31680 19024 31686
rect 18972 31622 19024 31628
rect 18880 31476 18932 31482
rect 18880 31418 18932 31424
rect 18984 31346 19012 31622
rect 18788 31340 18840 31346
rect 18788 31282 18840 31288
rect 18972 31340 19024 31346
rect 18972 31282 19024 31288
rect 18800 31142 18828 31282
rect 18788 31136 18840 31142
rect 18788 31078 18840 31084
rect 18696 30796 18748 30802
rect 18696 30738 18748 30744
rect 18604 30252 18656 30258
rect 18604 30194 18656 30200
rect 18512 29096 18564 29102
rect 18432 29056 18512 29084
rect 18512 29038 18564 29044
rect 18524 28762 18552 29038
rect 18512 28756 18564 28762
rect 18512 28698 18564 28704
rect 17868 28552 17920 28558
rect 17868 28494 17920 28500
rect 18616 28082 18644 30194
rect 18800 29458 18828 31078
rect 18984 29510 19012 31282
rect 18708 29430 18828 29458
rect 18972 29504 19024 29510
rect 18972 29446 19024 29452
rect 18604 28076 18656 28082
rect 18604 28018 18656 28024
rect 18420 27940 18472 27946
rect 18420 27882 18472 27888
rect 18328 27396 18380 27402
rect 18328 27338 18380 27344
rect 18144 26444 18196 26450
rect 18144 26386 18196 26392
rect 17868 26240 17920 26246
rect 17868 26182 17920 26188
rect 17880 25226 17908 26182
rect 18156 26042 18184 26386
rect 18144 26036 18196 26042
rect 18144 25978 18196 25984
rect 17868 25220 17920 25226
rect 17868 25162 17920 25168
rect 17776 25152 17828 25158
rect 17776 25094 17828 25100
rect 17880 24818 17908 25162
rect 17684 24812 17736 24818
rect 17684 24754 17736 24760
rect 17868 24812 17920 24818
rect 17868 24754 17920 24760
rect 17696 24342 17724 24754
rect 18156 24614 18184 25978
rect 18340 25362 18368 27338
rect 18432 27334 18460 27882
rect 18420 27328 18472 27334
rect 18420 27270 18472 27276
rect 18512 27328 18564 27334
rect 18512 27270 18564 27276
rect 18432 26586 18460 27270
rect 18420 26580 18472 26586
rect 18420 26522 18472 26528
rect 18524 25430 18552 27270
rect 18708 26926 18736 29430
rect 18788 29096 18840 29102
rect 18788 29038 18840 29044
rect 18800 28150 18828 29038
rect 18880 28552 18932 28558
rect 18880 28494 18932 28500
rect 18788 28144 18840 28150
rect 18788 28086 18840 28092
rect 18696 26920 18748 26926
rect 18696 26862 18748 26868
rect 18604 25900 18656 25906
rect 18604 25842 18656 25848
rect 18512 25424 18564 25430
rect 18512 25366 18564 25372
rect 18328 25356 18380 25362
rect 18328 25298 18380 25304
rect 18524 24818 18552 25366
rect 18616 25294 18644 25842
rect 18800 25430 18828 28086
rect 18892 28082 18920 28494
rect 18984 28082 19012 29446
rect 19076 29034 19104 31894
rect 19168 31414 19196 33390
rect 19260 33318 19288 33934
rect 19352 33658 19380 35158
rect 19720 35057 19748 35498
rect 19812 35086 19840 35550
rect 19892 35488 19944 35494
rect 19892 35430 19944 35436
rect 20168 35488 20220 35494
rect 20168 35430 20220 35436
rect 19904 35154 19932 35430
rect 19984 35284 20036 35290
rect 19984 35226 20036 35232
rect 19892 35148 19944 35154
rect 19892 35090 19944 35096
rect 19800 35080 19852 35086
rect 19706 35048 19762 35057
rect 19800 35022 19852 35028
rect 19996 35018 20024 35226
rect 19706 34983 19762 34992
rect 19984 35012 20036 35018
rect 19984 34954 20036 34960
rect 19432 34944 19484 34950
rect 19432 34886 19484 34892
rect 19444 34678 19472 34886
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19432 34672 19484 34678
rect 19432 34614 19484 34620
rect 19892 34536 19944 34542
rect 19892 34478 19944 34484
rect 19904 34406 19932 34478
rect 19892 34400 19944 34406
rect 19892 34342 19944 34348
rect 19522 34232 19578 34241
rect 19522 34167 19578 34176
rect 19536 34066 19564 34167
rect 19524 34060 19576 34066
rect 19524 34002 19576 34008
rect 19996 33862 20024 34954
rect 20076 34672 20128 34678
rect 20076 34614 20128 34620
rect 19432 33856 19484 33862
rect 19432 33798 19484 33804
rect 19984 33856 20036 33862
rect 19984 33798 20036 33804
rect 19340 33652 19392 33658
rect 19340 33594 19392 33600
rect 19352 33522 19380 33594
rect 19340 33516 19392 33522
rect 19340 33458 19392 33464
rect 19444 33454 19472 33798
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19800 33516 19852 33522
rect 19800 33458 19852 33464
rect 19432 33448 19484 33454
rect 19432 33390 19484 33396
rect 19248 33312 19300 33318
rect 19248 33254 19300 33260
rect 19260 31754 19288 33254
rect 19812 32774 19840 33458
rect 19432 32768 19484 32774
rect 19432 32710 19484 32716
rect 19800 32768 19852 32774
rect 19800 32710 19852 32716
rect 19984 32768 20036 32774
rect 19984 32710 20036 32716
rect 19260 31726 19380 31754
rect 19352 31686 19380 31726
rect 19340 31680 19392 31686
rect 19340 31622 19392 31628
rect 19156 31408 19208 31414
rect 19156 31350 19208 31356
rect 19340 30932 19392 30938
rect 19444 30920 19472 32710
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19708 32496 19760 32502
rect 19708 32438 19760 32444
rect 19720 31793 19748 32438
rect 19996 32366 20024 32710
rect 19984 32360 20036 32366
rect 19984 32302 20036 32308
rect 19706 31784 19762 31793
rect 19706 31719 19762 31728
rect 19984 31680 20036 31686
rect 19984 31622 20036 31628
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19996 31482 20024 31622
rect 19984 31476 20036 31482
rect 19984 31418 20036 31424
rect 19524 31408 19576 31414
rect 19524 31350 19576 31356
rect 19392 30892 19472 30920
rect 19340 30874 19392 30880
rect 19536 30818 19564 31350
rect 19892 31272 19944 31278
rect 19892 31214 19944 31220
rect 19904 30977 19932 31214
rect 19890 30968 19946 30977
rect 19708 30932 19760 30938
rect 19890 30903 19946 30912
rect 19708 30874 19760 30880
rect 19720 30841 19748 30874
rect 19352 30790 19564 30818
rect 19706 30832 19762 30841
rect 19156 30252 19208 30258
rect 19156 30194 19208 30200
rect 19168 29510 19196 30194
rect 19248 29572 19300 29578
rect 19248 29514 19300 29520
rect 19156 29504 19208 29510
rect 19156 29446 19208 29452
rect 19260 29186 19288 29514
rect 19168 29170 19288 29186
rect 19168 29164 19300 29170
rect 19168 29158 19248 29164
rect 19064 29028 19116 29034
rect 19064 28970 19116 28976
rect 18880 28076 18932 28082
rect 18880 28018 18932 28024
rect 18972 28076 19024 28082
rect 18972 28018 19024 28024
rect 18984 27538 19012 28018
rect 18972 27532 19024 27538
rect 18972 27474 19024 27480
rect 18880 27464 18932 27470
rect 18880 27406 18932 27412
rect 19064 27464 19116 27470
rect 19064 27406 19116 27412
rect 18892 26908 18920 27406
rect 18972 26920 19024 26926
rect 18892 26880 18972 26908
rect 18788 25424 18840 25430
rect 18788 25366 18840 25372
rect 18892 25294 18920 26880
rect 18972 26862 19024 26868
rect 19076 26790 19104 27406
rect 19168 27402 19196 29158
rect 19248 29106 19300 29112
rect 19352 28966 19380 30790
rect 19706 30767 19762 30776
rect 19904 30580 19932 30903
rect 19996 30734 20024 31418
rect 19984 30728 20036 30734
rect 19984 30670 20036 30676
rect 19904 30552 20024 30580
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19996 30258 20024 30552
rect 19984 30252 20036 30258
rect 19984 30194 20036 30200
rect 19984 29708 20036 29714
rect 19984 29650 20036 29656
rect 19432 29504 19484 29510
rect 19432 29446 19484 29452
rect 19444 29306 19472 29446
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19432 29300 19484 29306
rect 19432 29242 19484 29248
rect 19430 29200 19486 29209
rect 19430 29135 19432 29144
rect 19484 29135 19486 29144
rect 19432 29106 19484 29112
rect 19996 29102 20024 29650
rect 19616 29096 19668 29102
rect 19616 29038 19668 29044
rect 19984 29096 20036 29102
rect 19984 29038 20036 29044
rect 19340 28960 19392 28966
rect 19340 28902 19392 28908
rect 19340 28688 19392 28694
rect 19340 28630 19392 28636
rect 19156 27396 19208 27402
rect 19156 27338 19208 27344
rect 19168 26994 19196 27338
rect 19156 26988 19208 26994
rect 19156 26930 19208 26936
rect 19064 26784 19116 26790
rect 19064 26726 19116 26732
rect 19352 26353 19380 28630
rect 19628 28558 19656 29038
rect 19982 28928 20038 28937
rect 19982 28863 20038 28872
rect 19432 28552 19484 28558
rect 19432 28494 19484 28500
rect 19616 28552 19668 28558
rect 19616 28494 19668 28500
rect 19338 26344 19394 26353
rect 19338 26279 19394 26288
rect 19340 25764 19392 25770
rect 19340 25706 19392 25712
rect 19156 25492 19208 25498
rect 19156 25434 19208 25440
rect 18604 25288 18656 25294
rect 18604 25230 18656 25236
rect 18880 25288 18932 25294
rect 18880 25230 18932 25236
rect 18892 24954 18920 25230
rect 18972 25152 19024 25158
rect 18972 25094 19024 25100
rect 18880 24948 18932 24954
rect 18880 24890 18932 24896
rect 18512 24812 18564 24818
rect 18512 24754 18564 24760
rect 18144 24608 18196 24614
rect 18144 24550 18196 24556
rect 17684 24336 17736 24342
rect 17684 24278 17736 24284
rect 17592 24200 17644 24206
rect 17592 24142 17644 24148
rect 17592 24064 17644 24070
rect 17592 24006 17644 24012
rect 18144 24064 18196 24070
rect 18144 24006 18196 24012
rect 18788 24064 18840 24070
rect 18788 24006 18840 24012
rect 17222 22607 17278 22616
rect 17500 22636 17552 22642
rect 17132 22578 17184 22584
rect 17500 22578 17552 22584
rect 16856 22432 16908 22438
rect 16856 22374 16908 22380
rect 16580 22092 16632 22098
rect 16580 22034 16632 22040
rect 16764 22024 16816 22030
rect 16764 21966 16816 21972
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 16592 20466 16620 21830
rect 16672 21548 16724 21554
rect 16672 21490 16724 21496
rect 16580 20460 16632 20466
rect 16580 20402 16632 20408
rect 16488 20324 16540 20330
rect 16488 20266 16540 20272
rect 16500 20058 16528 20266
rect 16488 20052 16540 20058
rect 16488 19994 16540 20000
rect 16592 19922 16620 20402
rect 16684 19922 16712 21490
rect 16776 21010 16804 21966
rect 16948 21616 17000 21622
rect 16948 21558 17000 21564
rect 16764 21004 16816 21010
rect 16764 20946 16816 20952
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16672 19916 16724 19922
rect 16672 19858 16724 19864
rect 16304 19780 16356 19786
rect 16304 19722 16356 19728
rect 16580 19780 16632 19786
rect 16580 19722 16632 19728
rect 16592 19514 16620 19722
rect 16580 19508 16632 19514
rect 16580 19450 16632 19456
rect 16684 19446 16712 19858
rect 16672 19440 16724 19446
rect 16672 19382 16724 19388
rect 16684 18222 16712 19382
rect 16776 19242 16804 20946
rect 16764 19236 16816 19242
rect 16764 19178 16816 19184
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 16856 18080 16908 18086
rect 16856 18022 16908 18028
rect 16868 17746 16896 18022
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 16132 16590 16160 17478
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 15936 15360 15988 15366
rect 15936 15302 15988 15308
rect 15948 15026 15976 15302
rect 16040 15162 16068 15438
rect 16028 15156 16080 15162
rect 16028 15098 16080 15104
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 16580 15088 16632 15094
rect 16580 15030 16632 15036
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 15948 14550 15976 14962
rect 16592 14618 16620 15030
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 15936 14544 15988 14550
rect 15936 14486 15988 14492
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15764 12850 15792 13262
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15580 12306 15608 12786
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15672 12442 15700 12582
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15488 12158 15608 12186
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15488 11898 15516 12038
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15396 11150 15424 11630
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15396 10062 15424 10406
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15396 9722 15424 9998
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 14924 9648 14976 9654
rect 14924 9590 14976 9596
rect 15488 9194 15516 10610
rect 15580 9382 15608 12158
rect 15660 12164 15712 12170
rect 15660 12106 15712 12112
rect 15672 11762 15700 12106
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15672 10674 15700 11698
rect 15764 11286 15792 12786
rect 15752 11280 15804 11286
rect 15752 11222 15804 11228
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15672 9926 15700 10610
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 15672 9586 15700 9862
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15488 9166 15608 9194
rect 14924 8900 14976 8906
rect 14924 8842 14976 8848
rect 14936 8566 14964 8842
rect 14924 8560 14976 8566
rect 14924 8502 14976 8508
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14188 8288 14240 8294
rect 14188 8230 14240 8236
rect 14200 7886 14228 8230
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 13360 7472 13412 7478
rect 13360 7414 13412 7420
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 14200 7342 14228 7822
rect 14476 7410 14504 8366
rect 14844 7954 14872 8434
rect 14832 7948 14884 7954
rect 14832 7890 14884 7896
rect 14936 7886 14964 8502
rect 15580 8362 15608 9166
rect 15672 8974 15700 9522
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15568 8356 15620 8362
rect 15568 8298 15620 8304
rect 15580 8090 15608 8298
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 14740 7812 14792 7818
rect 14740 7754 14792 7760
rect 14752 7410 14780 7754
rect 15936 7472 15988 7478
rect 15936 7414 15988 7420
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 14200 6730 14228 7278
rect 14384 6769 14412 7346
rect 14476 7002 14504 7346
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14752 6934 14780 7346
rect 14740 6928 14792 6934
rect 14740 6870 14792 6876
rect 14740 6792 14792 6798
rect 14370 6760 14426 6769
rect 14188 6724 14240 6730
rect 14370 6695 14426 6704
rect 14738 6760 14740 6769
rect 14792 6760 14794 6769
rect 14738 6695 14794 6704
rect 14188 6666 14240 6672
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 15488 5710 15516 6054
rect 15476 5704 15528 5710
rect 15476 5646 15528 5652
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 15948 4622 15976 7414
rect 16040 6798 16068 13670
rect 16408 12306 16436 14418
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16500 12918 16528 13262
rect 16488 12912 16540 12918
rect 16488 12854 16540 12860
rect 16396 12300 16448 12306
rect 16396 12242 16448 12248
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 16316 7886 16344 8774
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16500 7886 16528 8366
rect 16684 8090 16712 14758
rect 16776 12714 16804 15098
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16868 14414 16896 14962
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16868 12986 16896 13262
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16764 12708 16816 12714
rect 16764 12650 16816 12656
rect 16960 12306 16988 21558
rect 17040 18828 17092 18834
rect 17040 18770 17092 18776
rect 17052 18290 17080 18770
rect 17144 18766 17172 22578
rect 17408 22568 17460 22574
rect 17408 22510 17460 22516
rect 17420 22166 17448 22510
rect 17408 22160 17460 22166
rect 17408 22102 17460 22108
rect 17224 21956 17276 21962
rect 17224 21898 17276 21904
rect 17236 20874 17264 21898
rect 17604 20942 17632 24006
rect 18052 23724 18104 23730
rect 18052 23666 18104 23672
rect 17592 20936 17644 20942
rect 17592 20878 17644 20884
rect 17224 20868 17276 20874
rect 17224 20810 17276 20816
rect 17868 20868 17920 20874
rect 17868 20810 17920 20816
rect 17960 20868 18012 20874
rect 17960 20810 18012 20816
rect 17592 20528 17644 20534
rect 17592 20470 17644 20476
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17316 19236 17368 19242
rect 17316 19178 17368 19184
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 17144 17134 17172 18702
rect 17328 18290 17356 19178
rect 17316 18284 17368 18290
rect 17316 18226 17368 18232
rect 17316 18080 17368 18086
rect 17316 18022 17368 18028
rect 17222 17912 17278 17921
rect 17222 17847 17278 17856
rect 17132 17128 17184 17134
rect 17132 17070 17184 17076
rect 17236 16250 17264 17847
rect 17328 17270 17356 18022
rect 17316 17264 17368 17270
rect 17316 17206 17368 17212
rect 17420 17082 17448 19790
rect 17604 19378 17632 20470
rect 17776 19780 17828 19786
rect 17776 19722 17828 19728
rect 17788 19378 17816 19722
rect 17592 19372 17644 19378
rect 17592 19314 17644 19320
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17880 18408 17908 20810
rect 17972 19394 18000 20810
rect 18064 20330 18092 23666
rect 18052 20324 18104 20330
rect 18052 20266 18104 20272
rect 18156 19854 18184 24006
rect 18800 23866 18828 24006
rect 18788 23860 18840 23866
rect 18788 23802 18840 23808
rect 18984 23118 19012 25094
rect 19168 24818 19196 25434
rect 19248 25424 19300 25430
rect 19248 25366 19300 25372
rect 19260 24886 19288 25366
rect 19248 24880 19300 24886
rect 19248 24822 19300 24828
rect 19156 24812 19208 24818
rect 19156 24754 19208 24760
rect 19064 24676 19116 24682
rect 19064 24618 19116 24624
rect 18420 23112 18472 23118
rect 18420 23054 18472 23060
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 18328 22976 18380 22982
rect 18328 22918 18380 22924
rect 18340 22642 18368 22918
rect 18432 22642 18460 23054
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 18420 22636 18472 22642
rect 18420 22578 18472 22584
rect 18512 22568 18564 22574
rect 18512 22510 18564 22516
rect 18420 21480 18472 21486
rect 18420 21422 18472 21428
rect 18236 20460 18288 20466
rect 18236 20402 18288 20408
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 17972 19366 18092 19394
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 17972 18970 18000 19246
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 17960 18420 18012 18426
rect 17880 18380 17960 18408
rect 17960 18362 18012 18368
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17512 17814 17540 18226
rect 17500 17808 17552 17814
rect 17500 17750 17552 17756
rect 18064 17728 18092 19366
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 18156 18970 18184 19110
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 18144 18080 18196 18086
rect 18144 18022 18196 18028
rect 17972 17700 18092 17728
rect 17972 17542 18000 17700
rect 18052 17604 18104 17610
rect 18052 17546 18104 17552
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 17328 17054 17448 17082
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 17052 14278 17080 14962
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 17236 13938 17264 14350
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 17236 12850 17264 13874
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 17040 12436 17092 12442
rect 17328 12434 17356 17054
rect 17972 16726 18000 17478
rect 18064 17202 18092 17546
rect 18156 17270 18184 18022
rect 18144 17264 18196 17270
rect 18144 17206 18196 17212
rect 18248 17202 18276 20402
rect 18432 19854 18460 21422
rect 18524 21146 18552 22510
rect 19076 22094 19104 24618
rect 19168 24206 19196 24754
rect 19248 24676 19300 24682
rect 19248 24618 19300 24624
rect 19260 24410 19288 24618
rect 19248 24404 19300 24410
rect 19248 24346 19300 24352
rect 19156 24200 19208 24206
rect 19156 24142 19208 24148
rect 19076 22066 19288 22094
rect 18512 21140 18564 21146
rect 18512 21082 18564 21088
rect 18512 20392 18564 20398
rect 18512 20334 18564 20340
rect 18524 19990 18552 20334
rect 18512 19984 18564 19990
rect 18512 19926 18564 19932
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18432 18834 18460 19790
rect 18512 19712 18564 19718
rect 18512 19654 18564 19660
rect 18788 19712 18840 19718
rect 18788 19654 18840 19660
rect 18524 19378 18552 19654
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 18420 18828 18472 18834
rect 18420 18770 18472 18776
rect 18524 18698 18552 19314
rect 18512 18692 18564 18698
rect 18512 18634 18564 18640
rect 18616 18630 18644 19314
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 18708 18222 18736 19110
rect 18696 18216 18748 18222
rect 18432 18154 18644 18170
rect 18696 18158 18748 18164
rect 18420 18148 18656 18154
rect 18472 18142 18604 18148
rect 18420 18090 18472 18096
rect 18604 18090 18656 18096
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18248 16794 18276 17138
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 17960 16720 18012 16726
rect 17960 16662 18012 16668
rect 17972 16522 18000 16662
rect 17960 16516 18012 16522
rect 17960 16458 18012 16464
rect 17592 16108 17644 16114
rect 17592 16050 17644 16056
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 17500 15904 17552 15910
rect 17500 15846 17552 15852
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17040 12378 17092 12384
rect 17144 12406 17356 12434
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 17052 12238 17080 12378
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16776 10062 16804 11834
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16776 9110 16804 9998
rect 16764 9104 16816 9110
rect 16764 9046 16816 9052
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16776 8498 16804 8910
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16684 7886 16712 8026
rect 16868 7886 16896 11018
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16960 9994 16988 10950
rect 16948 9988 17000 9994
rect 16948 9930 17000 9936
rect 17144 9178 17172 12406
rect 17222 12336 17278 12345
rect 17222 12271 17224 12280
rect 17276 12271 17278 12280
rect 17224 12242 17276 12248
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 17236 10810 17264 10950
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17420 10554 17448 13806
rect 17512 12850 17540 15846
rect 17604 15502 17632 16050
rect 17788 15706 17816 16050
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17788 15570 17816 15642
rect 17880 15638 17908 16050
rect 17868 15632 17920 15638
rect 17868 15574 17920 15580
rect 17776 15564 17828 15570
rect 17776 15506 17828 15512
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 17776 15428 17828 15434
rect 17776 15370 17828 15376
rect 17684 15360 17736 15366
rect 17684 15302 17736 15308
rect 17592 15020 17644 15026
rect 17592 14962 17644 14968
rect 17604 13394 17632 14962
rect 17696 14346 17724 15302
rect 17788 15026 17816 15370
rect 17868 15088 17920 15094
rect 17866 15056 17868 15065
rect 18052 15088 18104 15094
rect 17920 15056 17922 15065
rect 17776 15020 17828 15026
rect 18052 15030 18104 15036
rect 17866 14991 17922 15000
rect 17776 14962 17828 14968
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 17788 14482 17816 14758
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17684 14340 17736 14346
rect 17684 14282 17736 14288
rect 17880 14074 17908 14894
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 17972 14006 18000 14894
rect 18064 14414 18092 15030
rect 18328 14884 18380 14890
rect 18328 14826 18380 14832
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 17960 14000 18012 14006
rect 17960 13942 18012 13948
rect 18340 13870 18368 14826
rect 18800 14090 18828 19654
rect 19156 18964 19208 18970
rect 19156 18906 19208 18912
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18892 14278 18920 14962
rect 19168 14414 19196 18906
rect 18972 14408 19024 14414
rect 18972 14350 19024 14356
rect 19156 14408 19208 14414
rect 19156 14350 19208 14356
rect 18880 14272 18932 14278
rect 18880 14214 18932 14220
rect 18616 14062 18828 14090
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 18156 13462 18184 13670
rect 18144 13456 18196 13462
rect 18144 13398 18196 13404
rect 17592 13388 17644 13394
rect 17592 13330 17644 13336
rect 18156 13326 18184 13398
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 17776 13252 17828 13258
rect 17776 13194 17828 13200
rect 17788 12986 17816 13194
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17500 12844 17552 12850
rect 17788 12832 17816 12922
rect 17500 12786 17552 12792
rect 17604 12804 17816 12832
rect 17512 11830 17540 12786
rect 17604 12442 17632 12804
rect 17776 12708 17828 12714
rect 17776 12650 17828 12656
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17500 11824 17552 11830
rect 17500 11766 17552 11772
rect 17604 11150 17632 12378
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17696 11626 17724 12038
rect 17788 11762 17816 12650
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 17684 11620 17736 11626
rect 17684 11562 17736 11568
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17696 10742 17724 11562
rect 17788 11286 17816 11698
rect 18616 11286 18644 14062
rect 18696 14000 18748 14006
rect 18696 13942 18748 13948
rect 17776 11280 17828 11286
rect 17776 11222 17828 11228
rect 18052 11280 18104 11286
rect 18052 11222 18104 11228
rect 18604 11280 18656 11286
rect 18604 11222 18656 11228
rect 17684 10736 17736 10742
rect 17684 10678 17736 10684
rect 17328 10526 17448 10554
rect 17788 10538 17816 11222
rect 18064 10674 18092 11222
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 17776 10532 17828 10538
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17328 9042 17356 10526
rect 17776 10474 17828 10480
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17420 10062 17448 10406
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17512 9926 17540 10406
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 18064 9518 18092 10610
rect 18248 10606 18276 10950
rect 18524 10810 18552 11018
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 18708 10062 18736 13942
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18800 12238 18828 12378
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18432 9382 18460 9522
rect 18328 9376 18380 9382
rect 18328 9318 18380 9324
rect 18420 9376 18472 9382
rect 18420 9318 18472 9324
rect 17316 9036 17368 9042
rect 17316 8978 17368 8984
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17880 8838 17908 8910
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16488 7880 16540 7886
rect 16488 7822 16540 7828
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16224 6866 16252 7686
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16040 5710 16068 6734
rect 16224 6322 16252 6802
rect 16592 6730 16620 7686
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 17972 6866 18000 7210
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 16580 6724 16632 6730
rect 16580 6666 16632 6672
rect 16592 6390 16620 6666
rect 16580 6384 16632 6390
rect 16580 6326 16632 6332
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 17420 5914 17448 6734
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 17420 4690 17448 5850
rect 17972 5098 18000 6802
rect 18156 6746 18184 7278
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 18064 6730 18184 6746
rect 18052 6724 18184 6730
rect 18104 6718 18184 6724
rect 18052 6666 18104 6672
rect 18156 6322 18184 6718
rect 18144 6316 18196 6322
rect 18144 6258 18196 6264
rect 18248 5710 18276 7142
rect 18340 6798 18368 9318
rect 18420 9104 18472 9110
rect 18420 9046 18472 9052
rect 18432 7886 18460 9046
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18524 8566 18552 8910
rect 18512 8560 18564 8566
rect 18512 8502 18564 8508
rect 18800 8430 18828 8978
rect 18892 8906 18920 12038
rect 18984 11082 19012 14350
rect 19064 12232 19116 12238
rect 19064 12174 19116 12180
rect 19076 11898 19104 12174
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 18972 11076 19024 11082
rect 18972 11018 19024 11024
rect 19156 9580 19208 9586
rect 19260 9568 19288 22066
rect 19352 21350 19380 25706
rect 19444 25294 19472 28494
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19996 28121 20024 28863
rect 19982 28112 20038 28121
rect 19982 28047 19984 28056
rect 20036 28047 20038 28056
rect 19984 28018 20036 28024
rect 19996 27987 20024 28018
rect 20088 27878 20116 34614
rect 20180 33114 20208 35430
rect 20260 34468 20312 34474
rect 20260 34410 20312 34416
rect 20272 33998 20300 34410
rect 20260 33992 20312 33998
rect 20260 33934 20312 33940
rect 20260 33856 20312 33862
rect 20260 33798 20312 33804
rect 20168 33108 20220 33114
rect 20168 33050 20220 33056
rect 20168 32904 20220 32910
rect 20168 32846 20220 32852
rect 20180 31210 20208 32846
rect 20272 31754 20300 33798
rect 20364 33522 20392 35550
rect 20536 35488 20588 35494
rect 20536 35430 20588 35436
rect 20444 34944 20496 34950
rect 20444 34886 20496 34892
rect 20456 34746 20484 34886
rect 20444 34740 20496 34746
rect 20444 34682 20496 34688
rect 20548 34626 20576 35430
rect 20456 34598 20576 34626
rect 20352 33516 20404 33522
rect 20352 33458 20404 33464
rect 20364 33386 20392 33458
rect 20352 33380 20404 33386
rect 20352 33322 20404 33328
rect 20352 33108 20404 33114
rect 20352 33050 20404 33056
rect 20364 32502 20392 33050
rect 20456 32570 20484 34598
rect 20824 33930 20852 36042
rect 20904 35080 20956 35086
rect 20904 35022 20956 35028
rect 20916 34678 20944 35022
rect 20904 34672 20956 34678
rect 20904 34614 20956 34620
rect 20904 34196 20956 34202
rect 20904 34138 20956 34144
rect 20812 33924 20864 33930
rect 20812 33866 20864 33872
rect 20720 33856 20772 33862
rect 20720 33798 20772 33804
rect 20536 33108 20588 33114
rect 20536 33050 20588 33056
rect 20548 32910 20576 33050
rect 20732 33046 20760 33798
rect 20916 33318 20944 34138
rect 20812 33312 20864 33318
rect 20812 33254 20864 33260
rect 20904 33312 20956 33318
rect 20904 33254 20956 33260
rect 20720 33040 20772 33046
rect 20720 32982 20772 32988
rect 20536 32904 20588 32910
rect 20536 32846 20588 32852
rect 20720 32904 20772 32910
rect 20720 32846 20772 32852
rect 20444 32564 20496 32570
rect 20444 32506 20496 32512
rect 20352 32496 20404 32502
rect 20352 32438 20404 32444
rect 20444 31816 20496 31822
rect 20444 31758 20496 31764
rect 20272 31726 20392 31754
rect 20260 31340 20312 31346
rect 20260 31282 20312 31288
rect 20168 31204 20220 31210
rect 20168 31146 20220 31152
rect 20166 31104 20222 31113
rect 20166 31039 20222 31048
rect 20180 28098 20208 31039
rect 20272 30326 20300 31282
rect 20260 30320 20312 30326
rect 20260 30262 20312 30268
rect 20260 29640 20312 29646
rect 20260 29582 20312 29588
rect 20272 29170 20300 29582
rect 20260 29164 20312 29170
rect 20260 29106 20312 29112
rect 20258 29064 20314 29073
rect 20258 28999 20260 29008
rect 20312 28999 20314 29008
rect 20260 28970 20312 28976
rect 20180 28070 20300 28098
rect 20168 28008 20220 28014
rect 20168 27950 20220 27956
rect 20076 27872 20128 27878
rect 20076 27814 20128 27820
rect 20088 27470 20116 27814
rect 20076 27464 20128 27470
rect 19982 27432 20038 27441
rect 20076 27406 20128 27412
rect 19982 27367 20038 27376
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19996 26994 20024 27367
rect 20180 27130 20208 27950
rect 20168 27124 20220 27130
rect 20168 27066 20220 27072
rect 19984 26988 20036 26994
rect 19984 26930 20036 26936
rect 20168 26988 20220 26994
rect 20168 26930 20220 26936
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19996 25974 20024 26930
rect 20180 26897 20208 26930
rect 20166 26888 20222 26897
rect 20166 26823 20222 26832
rect 20272 26518 20300 28070
rect 20260 26512 20312 26518
rect 20260 26454 20312 26460
rect 19984 25968 20036 25974
rect 19984 25910 20036 25916
rect 20364 25906 20392 31726
rect 20456 30938 20484 31758
rect 20444 30932 20496 30938
rect 20444 30874 20496 30880
rect 20444 30796 20496 30802
rect 20444 30738 20496 30744
rect 20456 30376 20484 30738
rect 20548 30734 20576 32846
rect 20732 32570 20760 32846
rect 20720 32564 20772 32570
rect 20720 32506 20772 32512
rect 20628 32496 20680 32502
rect 20628 32438 20680 32444
rect 20536 30728 20588 30734
rect 20534 30696 20536 30705
rect 20588 30696 20590 30705
rect 20534 30631 20590 30640
rect 20456 30348 20576 30376
rect 20444 30252 20496 30258
rect 20444 30194 20496 30200
rect 20456 28694 20484 30194
rect 20548 29578 20576 30348
rect 20640 30138 20668 32438
rect 20732 31822 20760 32506
rect 20720 31816 20772 31822
rect 20720 31758 20772 31764
rect 20824 30841 20852 33254
rect 20904 32836 20956 32842
rect 20904 32778 20956 32784
rect 20916 32745 20944 32778
rect 20902 32736 20958 32745
rect 20902 32671 20958 32680
rect 20904 32564 20956 32570
rect 20904 32506 20956 32512
rect 20916 32434 20944 32506
rect 20904 32428 20956 32434
rect 20904 32370 20956 32376
rect 20904 31136 20956 31142
rect 20904 31078 20956 31084
rect 20916 30938 20944 31078
rect 20904 30932 20956 30938
rect 20904 30874 20956 30880
rect 20810 30832 20866 30841
rect 20810 30767 20866 30776
rect 20640 30110 20760 30138
rect 20628 30048 20680 30054
rect 20628 29990 20680 29996
rect 20640 29646 20668 29990
rect 20732 29782 20760 30110
rect 20720 29776 20772 29782
rect 20720 29718 20772 29724
rect 20628 29640 20680 29646
rect 20628 29582 20680 29588
rect 20536 29572 20588 29578
rect 20536 29514 20588 29520
rect 20444 28688 20496 28694
rect 20444 28630 20496 28636
rect 20548 28558 20576 29514
rect 20640 28626 20668 29582
rect 20720 29504 20772 29510
rect 20720 29446 20772 29452
rect 20732 29170 20760 29446
rect 20720 29164 20772 29170
rect 20720 29106 20772 29112
rect 20824 28966 20852 30767
rect 20904 30592 20956 30598
rect 20904 30534 20956 30540
rect 20812 28960 20864 28966
rect 20812 28902 20864 28908
rect 20628 28620 20680 28626
rect 20628 28562 20680 28568
rect 20536 28552 20588 28558
rect 20536 28494 20588 28500
rect 20444 28144 20496 28150
rect 20444 28086 20496 28092
rect 20352 25900 20404 25906
rect 20352 25842 20404 25848
rect 20456 25770 20484 28086
rect 20720 28008 20772 28014
rect 20720 27950 20772 27956
rect 20732 27674 20760 27950
rect 20720 27668 20772 27674
rect 20720 27610 20772 27616
rect 20812 26988 20864 26994
rect 20812 26930 20864 26936
rect 20628 26376 20680 26382
rect 20628 26318 20680 26324
rect 20720 26376 20772 26382
rect 20720 26318 20772 26324
rect 20640 25770 20668 26318
rect 20732 25906 20760 26318
rect 20720 25900 20772 25906
rect 20720 25842 20772 25848
rect 20076 25764 20128 25770
rect 20076 25706 20128 25712
rect 20444 25764 20496 25770
rect 20444 25706 20496 25712
rect 20628 25764 20680 25770
rect 20628 25706 20680 25712
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19432 25152 19484 25158
rect 19432 25094 19484 25100
rect 19444 21554 19472 25094
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 20088 24818 20116 25706
rect 20732 25226 20760 25842
rect 20720 25220 20772 25226
rect 20720 25162 20772 25168
rect 20536 25152 20588 25158
rect 20536 25094 20588 25100
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 19984 24744 20036 24750
rect 19984 24686 20036 24692
rect 19892 24676 19944 24682
rect 19892 24618 19944 24624
rect 19904 24342 19932 24618
rect 19892 24336 19944 24342
rect 19892 24278 19944 24284
rect 19904 24138 19932 24278
rect 19892 24132 19944 24138
rect 19892 24074 19944 24080
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19996 23610 20024 24686
rect 20444 24676 20496 24682
rect 20444 24618 20496 24624
rect 20260 24608 20312 24614
rect 20260 24550 20312 24556
rect 20272 24206 20300 24550
rect 20352 24336 20404 24342
rect 20352 24278 20404 24284
rect 20260 24200 20312 24206
rect 20260 24142 20312 24148
rect 20364 23746 20392 24278
rect 19904 23582 20024 23610
rect 20272 23718 20392 23746
rect 19904 23526 19932 23582
rect 19892 23520 19944 23526
rect 19892 23462 19944 23468
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 20088 22710 20116 23462
rect 20076 22704 20128 22710
rect 20076 22646 20128 22652
rect 19800 22500 19852 22506
rect 19800 22442 19852 22448
rect 19812 22234 19840 22442
rect 20168 22432 20220 22438
rect 20168 22374 20220 22380
rect 19800 22228 19852 22234
rect 19800 22170 19852 22176
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19444 20505 19472 21490
rect 20076 20800 20128 20806
rect 20076 20742 20128 20748
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19430 20496 19486 20505
rect 19430 20431 19486 20440
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 19352 19514 19380 20334
rect 19892 20052 19944 20058
rect 19892 19994 19944 20000
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19340 18284 19392 18290
rect 19340 18226 19392 18232
rect 19352 17338 19380 18226
rect 19444 18222 19472 19858
rect 19904 19854 19932 19994
rect 19892 19848 19944 19854
rect 19944 19808 20024 19836
rect 19892 19790 19944 19796
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19996 19378 20024 19808
rect 20088 19446 20116 20742
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 19996 18834 20024 19314
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 20180 18714 20208 22374
rect 20272 20058 20300 23718
rect 20456 23644 20484 24618
rect 20548 24342 20576 25094
rect 20536 24336 20588 24342
rect 20536 24278 20588 24284
rect 20364 23616 20484 23644
rect 20260 20052 20312 20058
rect 20260 19994 20312 20000
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 20272 19310 20300 19858
rect 20364 19360 20392 23616
rect 20536 23520 20588 23526
rect 20536 23462 20588 23468
rect 20548 23186 20576 23462
rect 20720 23316 20772 23322
rect 20720 23258 20772 23264
rect 20732 23225 20760 23258
rect 20718 23216 20774 23225
rect 20536 23180 20588 23186
rect 20536 23122 20588 23128
rect 20628 23180 20680 23186
rect 20718 23151 20774 23160
rect 20628 23122 20680 23128
rect 20444 22976 20496 22982
rect 20444 22918 20496 22924
rect 20456 22234 20484 22918
rect 20444 22228 20496 22234
rect 20444 22170 20496 22176
rect 20640 22094 20668 23122
rect 20720 22228 20772 22234
rect 20720 22170 20772 22176
rect 20456 22066 20668 22094
rect 20456 20534 20484 22066
rect 20534 21992 20590 22001
rect 20534 21927 20590 21936
rect 20548 20942 20576 21927
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 20444 20528 20496 20534
rect 20444 20470 20496 20476
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20548 20097 20576 20198
rect 20534 20088 20590 20097
rect 20534 20023 20590 20032
rect 20536 19984 20588 19990
rect 20536 19926 20588 19932
rect 20548 19514 20576 19926
rect 20536 19508 20588 19514
rect 20536 19450 20588 19456
rect 20536 19372 20588 19378
rect 20364 19332 20536 19360
rect 20536 19314 20588 19320
rect 20260 19304 20312 19310
rect 20260 19246 20312 19252
rect 20180 18686 20300 18714
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 20168 18624 20220 18630
rect 20168 18566 20220 18572
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 18426 20024 18566
rect 20074 18456 20130 18465
rect 19984 18420 20036 18426
rect 20074 18391 20130 18400
rect 19984 18362 20036 18368
rect 20088 18358 20116 18391
rect 20076 18352 20128 18358
rect 20076 18294 20128 18300
rect 19524 18284 19576 18290
rect 19524 18226 19576 18232
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 19432 18080 19484 18086
rect 19536 18068 19564 18226
rect 20180 18086 20208 18566
rect 19484 18040 19564 18068
rect 20168 18080 20220 18086
rect 19432 18022 19484 18028
rect 20168 18022 20220 18028
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19444 15144 19472 18022
rect 20168 17808 20220 17814
rect 20168 17750 20220 17756
rect 19524 17672 19576 17678
rect 19522 17640 19524 17649
rect 19576 17640 19578 17649
rect 19522 17575 19578 17584
rect 20076 17536 20128 17542
rect 20076 17478 20128 17484
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 20088 16590 20116 17478
rect 20076 16584 20128 16590
rect 20076 16526 20128 16532
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 20180 15638 20208 17750
rect 20168 15632 20220 15638
rect 20168 15574 20220 15580
rect 20180 15450 20208 15574
rect 20272 15570 20300 18686
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20088 15422 20208 15450
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19444 15116 19564 15144
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19352 14618 19380 14962
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19352 13938 19380 14214
rect 19444 14074 19472 14962
rect 19536 14385 19564 15116
rect 19708 14952 19760 14958
rect 19708 14894 19760 14900
rect 19720 14618 19748 14894
rect 19708 14612 19760 14618
rect 19708 14554 19760 14560
rect 19522 14376 19578 14385
rect 19522 14311 19578 14320
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19430 13968 19486 13977
rect 19340 13932 19392 13938
rect 19430 13903 19486 13912
rect 19340 13874 19392 13880
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19352 12850 19380 13126
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 19340 12164 19392 12170
rect 19340 12106 19392 12112
rect 19352 11898 19380 12106
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19340 11688 19392 11694
rect 19340 11630 19392 11636
rect 19352 11218 19380 11630
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19208 9540 19288 9568
rect 19156 9522 19208 9528
rect 19260 8906 19288 9540
rect 18880 8900 18932 8906
rect 18880 8842 18932 8848
rect 19248 8900 19300 8906
rect 19248 8842 19300 8848
rect 18892 8498 18920 8842
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18788 8424 18840 8430
rect 18788 8366 18840 8372
rect 18696 8288 18748 8294
rect 18696 8230 18748 8236
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18616 7410 18644 7890
rect 18708 7886 18736 8230
rect 18800 8090 18828 8366
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18708 7478 18736 7822
rect 18696 7472 18748 7478
rect 18696 7414 18748 7420
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18328 6792 18380 6798
rect 18328 6734 18380 6740
rect 18432 6390 18460 6802
rect 18420 6384 18472 6390
rect 18420 6326 18472 6332
rect 18616 6322 18644 7346
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 18694 6760 18750 6769
rect 18694 6695 18750 6704
rect 18708 6662 18736 6695
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 18800 5710 18828 7278
rect 18972 6384 19024 6390
rect 18972 6326 19024 6332
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18328 5568 18380 5574
rect 18328 5510 18380 5516
rect 18340 5302 18368 5510
rect 18328 5296 18380 5302
rect 18328 5238 18380 5244
rect 18984 5166 19012 6326
rect 18972 5160 19024 5166
rect 18972 5102 19024 5108
rect 17960 5092 18012 5098
rect 17960 5034 18012 5040
rect 18512 5024 18564 5030
rect 18512 4966 18564 4972
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 15948 4146 15976 4558
rect 18524 4146 18552 4966
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 19444 4078 19472 13903
rect 19996 13394 20024 14214
rect 20088 13938 20116 15422
rect 20168 15360 20220 15366
rect 20168 15302 20220 15308
rect 20180 14482 20208 15302
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 20272 14006 20300 15506
rect 20364 15162 20392 18566
rect 20548 16114 20576 19314
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20640 15994 20668 18906
rect 20548 15966 20668 15994
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20352 14884 20404 14890
rect 20352 14826 20404 14832
rect 20364 14278 20392 14826
rect 20352 14272 20404 14278
rect 20352 14214 20404 14220
rect 20260 14000 20312 14006
rect 20260 13942 20312 13948
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19706 12880 19762 12889
rect 20258 12880 20314 12889
rect 19706 12815 19708 12824
rect 19760 12815 19762 12824
rect 19984 12844 20036 12850
rect 19708 12786 19760 12792
rect 20258 12815 20314 12824
rect 19984 12786 20036 12792
rect 19708 12640 19760 12646
rect 19708 12582 19760 12588
rect 19720 12238 19748 12582
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 19720 11694 19748 11834
rect 19996 11762 20024 12786
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 20088 12238 20116 12718
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19996 11354 20024 11698
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 20180 11218 20208 12378
rect 20272 11898 20300 12815
rect 20260 11892 20312 11898
rect 20260 11834 20312 11840
rect 20272 11762 20300 11834
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19892 9512 19944 9518
rect 19892 9454 19944 9460
rect 19904 8838 19932 9454
rect 20180 9042 20208 11154
rect 20364 10130 20392 13874
rect 20444 12164 20496 12170
rect 20444 12106 20496 12112
rect 20456 11150 20484 12106
rect 20444 11144 20496 11150
rect 20444 11086 20496 11092
rect 20548 10266 20576 15966
rect 20732 15026 20760 22170
rect 20824 19922 20852 26930
rect 20916 26926 20944 30534
rect 21008 28014 21036 36042
rect 22112 35834 22140 36722
rect 22480 36038 22508 37062
rect 24320 36718 24348 37130
rect 23020 36712 23072 36718
rect 23020 36654 23072 36660
rect 24308 36712 24360 36718
rect 24308 36654 24360 36660
rect 22928 36168 22980 36174
rect 22928 36110 22980 36116
rect 22468 36032 22520 36038
rect 22468 35974 22520 35980
rect 22100 35828 22152 35834
rect 22100 35770 22152 35776
rect 22480 35698 22508 35974
rect 22940 35834 22968 36110
rect 22928 35828 22980 35834
rect 22928 35770 22980 35776
rect 22468 35692 22520 35698
rect 22468 35634 22520 35640
rect 22928 35692 22980 35698
rect 22928 35634 22980 35640
rect 21364 35624 21416 35630
rect 21364 35566 21416 35572
rect 21088 34944 21140 34950
rect 21088 34886 21140 34892
rect 20996 28008 21048 28014
rect 20996 27950 21048 27956
rect 20996 27056 21048 27062
rect 20996 26998 21048 27004
rect 20904 26920 20956 26926
rect 20904 26862 20956 26868
rect 21008 26489 21036 26998
rect 20994 26480 21050 26489
rect 20994 26415 21050 26424
rect 20904 25900 20956 25906
rect 20904 25842 20956 25848
rect 20916 23186 20944 25842
rect 20996 25832 21048 25838
rect 20996 25774 21048 25780
rect 21008 25294 21036 25774
rect 20996 25288 21048 25294
rect 20996 25230 21048 25236
rect 21100 24886 21128 34886
rect 21376 34678 21404 35566
rect 22008 35080 22060 35086
rect 22008 35022 22060 35028
rect 21364 34672 21416 34678
rect 21364 34614 21416 34620
rect 21272 33516 21324 33522
rect 21272 33458 21324 33464
rect 21284 32774 21312 33458
rect 21272 32768 21324 32774
rect 21272 32710 21324 32716
rect 21180 32360 21232 32366
rect 21376 32348 21404 34614
rect 22020 34610 22048 35022
rect 22744 34944 22796 34950
rect 22744 34886 22796 34892
rect 21824 34604 21876 34610
rect 21824 34546 21876 34552
rect 22008 34604 22060 34610
rect 22008 34546 22060 34552
rect 22376 34604 22428 34610
rect 22376 34546 22428 34552
rect 21836 34354 21864 34546
rect 22284 34536 22336 34542
rect 22020 34462 22232 34490
rect 22284 34478 22336 34484
rect 22020 34354 22048 34462
rect 21836 34326 22048 34354
rect 21732 34196 21784 34202
rect 21732 34138 21784 34144
rect 21548 34060 21600 34066
rect 21548 34002 21600 34008
rect 21456 33312 21508 33318
rect 21456 33254 21508 33260
rect 21232 32320 21404 32348
rect 21180 32302 21232 32308
rect 21192 29646 21220 32302
rect 21272 32224 21324 32230
rect 21272 32166 21324 32172
rect 21180 29640 21232 29646
rect 21180 29582 21232 29588
rect 21192 26897 21220 29582
rect 21178 26888 21234 26897
rect 21178 26823 21234 26832
rect 21284 26518 21312 32166
rect 21468 31754 21496 33254
rect 21560 31822 21588 34002
rect 21640 33924 21692 33930
rect 21640 33866 21692 33872
rect 21652 33658 21680 33866
rect 21640 33652 21692 33658
rect 21640 33594 21692 33600
rect 21652 32978 21680 33594
rect 21640 32972 21692 32978
rect 21640 32914 21692 32920
rect 21640 32768 21692 32774
rect 21640 32710 21692 32716
rect 21652 31906 21680 32710
rect 21744 32026 21772 34138
rect 21822 33960 21878 33969
rect 22204 33930 22232 34462
rect 22296 34066 22324 34478
rect 22388 34406 22416 34546
rect 22376 34400 22428 34406
rect 22376 34342 22428 34348
rect 22652 34400 22704 34406
rect 22652 34342 22704 34348
rect 22284 34060 22336 34066
rect 22284 34002 22336 34008
rect 22388 33998 22416 34342
rect 22664 33998 22692 34342
rect 22756 33998 22784 34886
rect 22376 33992 22428 33998
rect 22376 33934 22428 33940
rect 22652 33992 22704 33998
rect 22744 33992 22796 33998
rect 22652 33934 22704 33940
rect 22742 33960 22744 33969
rect 22796 33960 22798 33969
rect 21822 33895 21878 33904
rect 22192 33924 22244 33930
rect 21836 32502 21864 33895
rect 22192 33866 22244 33872
rect 22284 33856 22336 33862
rect 22284 33798 22336 33804
rect 22100 33448 22152 33454
rect 22100 33390 22152 33396
rect 21824 32496 21876 32502
rect 21824 32438 21876 32444
rect 21822 32328 21878 32337
rect 22112 32314 22140 33390
rect 22296 32570 22324 33798
rect 22468 33516 22520 33522
rect 22468 33458 22520 33464
rect 22480 32978 22508 33458
rect 22664 33114 22692 33934
rect 22742 33895 22798 33904
rect 22744 33856 22796 33862
rect 22744 33798 22796 33804
rect 22756 33658 22784 33798
rect 22744 33652 22796 33658
rect 22744 33594 22796 33600
rect 22756 33522 22784 33594
rect 22744 33516 22796 33522
rect 22744 33458 22796 33464
rect 22652 33108 22704 33114
rect 22652 33050 22704 33056
rect 22756 33046 22784 33458
rect 22744 33040 22796 33046
rect 22744 32982 22796 32988
rect 22468 32972 22520 32978
rect 22468 32914 22520 32920
rect 22284 32564 22336 32570
rect 22284 32506 22336 32512
rect 22376 32360 22428 32366
rect 22296 32320 22376 32348
rect 22112 32286 22232 32314
rect 21822 32263 21824 32272
rect 21876 32263 21878 32272
rect 21824 32234 21876 32240
rect 21732 32020 21784 32026
rect 21732 31962 21784 31968
rect 21652 31878 21772 31906
rect 21548 31816 21600 31822
rect 21548 31758 21600 31764
rect 21744 31754 21772 31878
rect 21376 31726 21496 31754
rect 21732 31748 21784 31754
rect 21376 29714 21404 31726
rect 21732 31690 21784 31696
rect 21456 31340 21508 31346
rect 21456 31282 21508 31288
rect 21468 30802 21496 31282
rect 21548 31272 21600 31278
rect 21548 31214 21600 31220
rect 21456 30796 21508 30802
rect 21456 30738 21508 30744
rect 21364 29708 21416 29714
rect 21364 29650 21416 29656
rect 21456 29096 21508 29102
rect 21456 29038 21508 29044
rect 21364 28552 21416 28558
rect 21364 28494 21416 28500
rect 21272 26512 21324 26518
rect 21272 26454 21324 26460
rect 21178 25936 21234 25945
rect 21178 25871 21234 25880
rect 21088 24880 21140 24886
rect 21088 24822 21140 24828
rect 21086 24168 21142 24177
rect 21086 24103 21142 24112
rect 21100 24070 21128 24103
rect 20996 24064 21048 24070
rect 20996 24006 21048 24012
rect 21088 24064 21140 24070
rect 21088 24006 21140 24012
rect 21008 23186 21036 24006
rect 20904 23180 20956 23186
rect 20904 23122 20956 23128
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 21100 22778 21128 24006
rect 21192 23866 21220 25871
rect 21376 25498 21404 28494
rect 21468 27520 21496 29038
rect 21560 28762 21588 31214
rect 21732 28960 21784 28966
rect 21732 28902 21784 28908
rect 21548 28756 21600 28762
rect 21548 28698 21600 28704
rect 21560 28150 21588 28698
rect 21640 28552 21692 28558
rect 21640 28494 21692 28500
rect 21548 28144 21600 28150
rect 21548 28086 21600 28092
rect 21652 27674 21680 28494
rect 21640 27668 21692 27674
rect 21640 27610 21692 27616
rect 21468 27492 21680 27520
rect 21652 26466 21680 27492
rect 21468 26438 21680 26466
rect 21468 25906 21496 26438
rect 21548 26376 21600 26382
rect 21548 26318 21600 26324
rect 21456 25900 21508 25906
rect 21456 25842 21508 25848
rect 21560 25809 21588 26318
rect 21640 26240 21692 26246
rect 21640 26182 21692 26188
rect 21652 26042 21680 26182
rect 21640 26036 21692 26042
rect 21640 25978 21692 25984
rect 21546 25800 21602 25809
rect 21546 25735 21602 25744
rect 21364 25492 21416 25498
rect 21364 25434 21416 25440
rect 21364 24132 21416 24138
rect 21364 24074 21416 24080
rect 21180 23860 21232 23866
rect 21180 23802 21232 23808
rect 21272 23792 21324 23798
rect 21272 23734 21324 23740
rect 21284 23322 21312 23734
rect 21376 23662 21404 24074
rect 21364 23656 21416 23662
rect 21364 23598 21416 23604
rect 21272 23316 21324 23322
rect 21272 23258 21324 23264
rect 21088 22772 21140 22778
rect 21088 22714 21140 22720
rect 21560 22642 21588 25735
rect 21652 25294 21680 25978
rect 21640 25288 21692 25294
rect 21640 25230 21692 25236
rect 21640 22976 21692 22982
rect 21638 22944 21640 22953
rect 21692 22944 21694 22953
rect 21638 22879 21694 22888
rect 21652 22778 21680 22879
rect 21640 22772 21692 22778
rect 21640 22714 21692 22720
rect 21548 22636 21600 22642
rect 21548 22578 21600 22584
rect 21744 22094 21772 28902
rect 21836 28558 21864 32234
rect 21916 31816 21968 31822
rect 21916 31758 21968 31764
rect 21928 29238 21956 31758
rect 22008 31476 22060 31482
rect 22008 31418 22060 31424
rect 22020 30938 22048 31418
rect 22008 30932 22060 30938
rect 22008 30874 22060 30880
rect 22100 30252 22152 30258
rect 22100 30194 22152 30200
rect 22112 29850 22140 30194
rect 22204 29850 22232 32286
rect 22296 31346 22324 32320
rect 22376 32302 22428 32308
rect 22480 31890 22508 32914
rect 22560 32904 22612 32910
rect 22560 32846 22612 32852
rect 22468 31884 22520 31890
rect 22468 31826 22520 31832
rect 22572 31754 22600 32846
rect 22756 32842 22784 32982
rect 22744 32836 22796 32842
rect 22744 32778 22796 32784
rect 22652 32768 22704 32774
rect 22652 32710 22704 32716
rect 22376 31748 22428 31754
rect 22376 31690 22428 31696
rect 22560 31748 22612 31754
rect 22560 31690 22612 31696
rect 22388 31414 22416 31690
rect 22376 31408 22428 31414
rect 22376 31350 22428 31356
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22560 31136 22612 31142
rect 22560 31078 22612 31084
rect 22284 30932 22336 30938
rect 22284 30874 22336 30880
rect 22296 30734 22324 30874
rect 22284 30728 22336 30734
rect 22284 30670 22336 30676
rect 22374 30696 22430 30705
rect 22374 30631 22430 30640
rect 22100 29844 22152 29850
rect 22100 29786 22152 29792
rect 22192 29844 22244 29850
rect 22192 29786 22244 29792
rect 22008 29708 22060 29714
rect 22008 29650 22060 29656
rect 21916 29232 21968 29238
rect 21916 29174 21968 29180
rect 21928 29073 21956 29174
rect 22020 29170 22048 29650
rect 22284 29300 22336 29306
rect 22284 29242 22336 29248
rect 22008 29164 22060 29170
rect 22008 29106 22060 29112
rect 21914 29064 21970 29073
rect 21914 28999 21970 29008
rect 21824 28552 21876 28558
rect 21824 28494 21876 28500
rect 21928 27606 21956 28999
rect 22296 28966 22324 29242
rect 22284 28960 22336 28966
rect 22284 28902 22336 28908
rect 22100 28416 22152 28422
rect 22100 28358 22152 28364
rect 22112 28082 22140 28358
rect 22100 28076 22152 28082
rect 22100 28018 22152 28024
rect 22284 28008 22336 28014
rect 22284 27950 22336 27956
rect 22008 27872 22060 27878
rect 22008 27814 22060 27820
rect 21916 27600 21968 27606
rect 21916 27542 21968 27548
rect 21916 27396 21968 27402
rect 21916 27338 21968 27344
rect 21928 26790 21956 27338
rect 22020 27062 22048 27814
rect 22008 27056 22060 27062
rect 22008 26998 22060 27004
rect 22192 26920 22244 26926
rect 22192 26862 22244 26868
rect 21916 26784 21968 26790
rect 21916 26726 21968 26732
rect 21824 26580 21876 26586
rect 21824 26522 21876 26528
rect 21836 25294 21864 26522
rect 21824 25288 21876 25294
rect 21824 25230 21876 25236
rect 21836 24206 21864 25230
rect 21928 25129 21956 26726
rect 22008 26580 22060 26586
rect 22008 26522 22060 26528
rect 22020 26450 22048 26522
rect 22008 26444 22060 26450
rect 22008 26386 22060 26392
rect 21914 25120 21970 25129
rect 21914 25055 21970 25064
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 21824 22704 21876 22710
rect 21824 22646 21876 22652
rect 21836 22234 21864 22646
rect 22204 22234 22232 26862
rect 21824 22228 21876 22234
rect 21824 22170 21876 22176
rect 22192 22228 22244 22234
rect 22192 22170 22244 22176
rect 22296 22094 22324 27950
rect 22388 27062 22416 30631
rect 22572 30122 22600 31078
rect 22664 30240 22692 32710
rect 22756 30734 22784 32778
rect 22836 32428 22888 32434
rect 22836 32370 22888 32376
rect 22848 32026 22876 32370
rect 22836 32020 22888 32026
rect 22836 31962 22888 31968
rect 22940 31754 22968 35634
rect 23032 34202 23060 36654
rect 23388 36576 23440 36582
rect 23388 36518 23440 36524
rect 23400 36174 23428 36518
rect 23388 36168 23440 36174
rect 23388 36110 23440 36116
rect 23756 36100 23808 36106
rect 23756 36042 23808 36048
rect 23848 36100 23900 36106
rect 23848 36042 23900 36048
rect 23204 35828 23256 35834
rect 23204 35770 23256 35776
rect 23216 35698 23244 35770
rect 23204 35692 23256 35698
rect 23204 35634 23256 35640
rect 23664 35488 23716 35494
rect 23664 35430 23716 35436
rect 23572 35284 23624 35290
rect 23572 35226 23624 35232
rect 23584 35154 23612 35226
rect 23572 35148 23624 35154
rect 23572 35090 23624 35096
rect 23204 35080 23256 35086
rect 23204 35022 23256 35028
rect 23216 34542 23244 35022
rect 23676 35018 23704 35430
rect 23664 35012 23716 35018
rect 23664 34954 23716 34960
rect 23676 34542 23704 34954
rect 23204 34536 23256 34542
rect 23204 34478 23256 34484
rect 23664 34536 23716 34542
rect 23664 34478 23716 34484
rect 23572 34468 23624 34474
rect 23572 34410 23624 34416
rect 23020 34196 23072 34202
rect 23020 34138 23072 34144
rect 23584 33998 23612 34410
rect 23676 34082 23704 34478
rect 23768 34241 23796 36042
rect 23860 35154 23888 36042
rect 23848 35148 23900 35154
rect 23848 35090 23900 35096
rect 23860 34746 23888 35090
rect 23848 34740 23900 34746
rect 23848 34682 23900 34688
rect 23754 34232 23810 34241
rect 23860 34202 23888 34682
rect 23754 34167 23810 34176
rect 23848 34196 23900 34202
rect 23848 34138 23900 34144
rect 23676 34054 23796 34082
rect 23572 33992 23624 33998
rect 23572 33934 23624 33940
rect 23020 33924 23072 33930
rect 23020 33866 23072 33872
rect 23032 32978 23060 33866
rect 23388 33584 23440 33590
rect 23388 33526 23440 33532
rect 23204 33380 23256 33386
rect 23204 33322 23256 33328
rect 23020 32972 23072 32978
rect 23020 32914 23072 32920
rect 23032 32434 23060 32914
rect 23112 32768 23164 32774
rect 23112 32710 23164 32716
rect 23020 32428 23072 32434
rect 23020 32370 23072 32376
rect 23124 32337 23152 32710
rect 23110 32328 23166 32337
rect 23020 32292 23072 32298
rect 23110 32263 23166 32272
rect 23020 32234 23072 32240
rect 22848 31726 22968 31754
rect 22744 30728 22796 30734
rect 22744 30670 22796 30676
rect 22848 30258 22876 31726
rect 23032 30802 23060 32234
rect 23216 31890 23244 33322
rect 23400 33046 23428 33526
rect 23388 33040 23440 33046
rect 23584 32994 23612 33934
rect 23768 33454 23796 34054
rect 23860 33998 23888 34138
rect 23848 33992 23900 33998
rect 23848 33934 23900 33940
rect 24216 33652 24268 33658
rect 24216 33594 24268 33600
rect 24228 33522 24256 33594
rect 24216 33516 24268 33522
rect 24216 33458 24268 33464
rect 23756 33448 23808 33454
rect 23756 33390 23808 33396
rect 24032 33448 24084 33454
rect 24032 33390 24084 33396
rect 23768 33318 23796 33390
rect 23756 33312 23808 33318
rect 23756 33254 23808 33260
rect 23388 32982 23440 32988
rect 23492 32966 23612 32994
rect 23296 32224 23348 32230
rect 23296 32166 23348 32172
rect 23308 31890 23336 32166
rect 23388 31952 23440 31958
rect 23388 31894 23440 31900
rect 23204 31884 23256 31890
rect 23204 31826 23256 31832
rect 23296 31884 23348 31890
rect 23296 31826 23348 31832
rect 23020 30796 23072 30802
rect 23020 30738 23072 30744
rect 23204 30796 23256 30802
rect 23204 30738 23256 30744
rect 22928 30660 22980 30666
rect 22928 30602 22980 30608
rect 22744 30252 22796 30258
rect 22664 30212 22744 30240
rect 22744 30194 22796 30200
rect 22836 30252 22888 30258
rect 22836 30194 22888 30200
rect 22560 30116 22612 30122
rect 22560 30058 22612 30064
rect 22572 29646 22600 30058
rect 22652 29776 22704 29782
rect 22652 29718 22704 29724
rect 22560 29640 22612 29646
rect 22560 29582 22612 29588
rect 22664 29102 22692 29718
rect 22652 29096 22704 29102
rect 22652 29038 22704 29044
rect 22560 29028 22612 29034
rect 22560 28970 22612 28976
rect 22572 28150 22600 28970
rect 22652 28484 22704 28490
rect 22652 28426 22704 28432
rect 22560 28144 22612 28150
rect 22560 28086 22612 28092
rect 22376 27056 22428 27062
rect 22376 26998 22428 27004
rect 22572 26994 22600 28086
rect 22560 26988 22612 26994
rect 22560 26930 22612 26936
rect 22376 26784 22428 26790
rect 22374 26752 22376 26761
rect 22428 26752 22430 26761
rect 22374 26687 22430 26696
rect 22376 26376 22428 26382
rect 22376 26318 22428 26324
rect 22388 24410 22416 26318
rect 22468 26036 22520 26042
rect 22468 25978 22520 25984
rect 22376 24404 22428 24410
rect 22376 24346 22428 24352
rect 22388 24274 22416 24346
rect 22376 24268 22428 24274
rect 22376 24210 22428 24216
rect 22480 24154 22508 25978
rect 22664 24954 22692 28426
rect 22756 27470 22784 30194
rect 22744 27464 22796 27470
rect 22744 27406 22796 27412
rect 22744 26988 22796 26994
rect 22744 26930 22796 26936
rect 22756 26586 22784 26930
rect 22744 26580 22796 26586
rect 22744 26522 22796 26528
rect 22848 26450 22876 30194
rect 22940 30122 22968 30602
rect 23216 30394 23244 30738
rect 23400 30705 23428 31894
rect 23492 31822 23520 32966
rect 23572 32904 23624 32910
rect 23572 32846 23624 32852
rect 23480 31816 23532 31822
rect 23480 31758 23532 31764
rect 23584 31482 23612 32846
rect 23664 32020 23716 32026
rect 23664 31962 23716 31968
rect 23572 31476 23624 31482
rect 23572 31418 23624 31424
rect 23676 31346 23704 31962
rect 23768 31346 23796 33254
rect 23848 32904 23900 32910
rect 23848 32846 23900 32852
rect 23664 31340 23716 31346
rect 23664 31282 23716 31288
rect 23756 31340 23808 31346
rect 23756 31282 23808 31288
rect 23480 31204 23532 31210
rect 23480 31146 23532 31152
rect 23492 30734 23520 31146
rect 23480 30728 23532 30734
rect 23386 30696 23442 30705
rect 23480 30670 23532 30676
rect 23572 30728 23624 30734
rect 23572 30670 23624 30676
rect 23386 30631 23442 30640
rect 23204 30388 23256 30394
rect 23204 30330 23256 30336
rect 23216 30190 23244 30330
rect 23020 30184 23072 30190
rect 23204 30184 23256 30190
rect 23072 30132 23152 30138
rect 23020 30126 23152 30132
rect 23204 30126 23256 30132
rect 22928 30116 22980 30122
rect 23032 30110 23152 30126
rect 22928 30058 22980 30064
rect 22940 29306 22968 30058
rect 23020 29640 23072 29646
rect 23020 29582 23072 29588
rect 22928 29300 22980 29306
rect 22928 29242 22980 29248
rect 23032 29186 23060 29582
rect 22940 29158 23060 29186
rect 22940 28422 22968 29158
rect 22928 28416 22980 28422
rect 22928 28358 22980 28364
rect 22836 26444 22888 26450
rect 22836 26386 22888 26392
rect 22652 24948 22704 24954
rect 22652 24890 22704 24896
rect 22560 24608 22612 24614
rect 22560 24550 22612 24556
rect 21652 22066 21772 22094
rect 22204 22066 22324 22094
rect 22388 24126 22508 24154
rect 20996 20800 21048 20806
rect 20996 20742 21048 20748
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20824 19446 20852 19858
rect 20916 19854 20944 20334
rect 21008 20330 21036 20742
rect 21362 20360 21418 20369
rect 20996 20324 21048 20330
rect 21362 20295 21418 20304
rect 20996 20266 21048 20272
rect 21376 19854 21404 20295
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 20812 19440 20864 19446
rect 20812 19382 20864 19388
rect 20824 19174 20852 19382
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 21376 18698 21404 19790
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 21364 18692 21416 18698
rect 21364 18634 21416 18640
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21284 17513 21312 17614
rect 21270 17504 21326 17513
rect 21270 17439 21326 17448
rect 21086 17232 21142 17241
rect 21086 17167 21142 17176
rect 21100 15094 21128 17167
rect 21088 15088 21140 15094
rect 21088 15030 21140 15036
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20628 12640 20680 12646
rect 20628 12582 20680 12588
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20168 9036 20220 9042
rect 20168 8978 20220 8984
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 20548 8430 20576 9318
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 19984 8356 20036 8362
rect 19984 8298 20036 8304
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19996 6798 20024 8298
rect 20640 7954 20668 12582
rect 20732 12442 20760 14758
rect 20904 14544 20956 14550
rect 20904 14486 20956 14492
rect 20916 13326 20944 14486
rect 21376 13802 21404 18634
rect 21560 17882 21588 18770
rect 21548 17876 21600 17882
rect 21548 17818 21600 17824
rect 21456 17604 21508 17610
rect 21456 17546 21508 17552
rect 21468 15502 21496 17546
rect 21652 16182 21680 22066
rect 22100 21684 22152 21690
rect 22100 21626 22152 21632
rect 21824 21412 21876 21418
rect 21824 21354 21876 21360
rect 21836 21146 21864 21354
rect 21824 21140 21876 21146
rect 21824 21082 21876 21088
rect 21836 16590 21864 21082
rect 22112 20466 22140 21626
rect 22204 21554 22232 22066
rect 22388 21554 22416 24126
rect 22572 23322 22600 24550
rect 22664 24070 22692 24890
rect 22742 24712 22798 24721
rect 22742 24647 22798 24656
rect 22756 24614 22784 24647
rect 22744 24608 22796 24614
rect 22744 24550 22796 24556
rect 22742 24440 22798 24449
rect 22742 24375 22798 24384
rect 22756 24206 22784 24375
rect 22744 24200 22796 24206
rect 22744 24142 22796 24148
rect 22652 24064 22704 24070
rect 22652 24006 22704 24012
rect 22836 23724 22888 23730
rect 22836 23666 22888 23672
rect 22560 23316 22612 23322
rect 22560 23258 22612 23264
rect 22652 22636 22704 22642
rect 22652 22578 22704 22584
rect 22468 22228 22520 22234
rect 22468 22170 22520 22176
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22100 20460 22152 20466
rect 22100 20402 22152 20408
rect 22100 19984 22152 19990
rect 22100 19926 22152 19932
rect 21914 19816 21970 19825
rect 21914 19751 21916 19760
rect 21968 19751 21970 19760
rect 21916 19722 21968 19728
rect 21914 18864 21970 18873
rect 21914 18799 21970 18808
rect 21928 18766 21956 18799
rect 21916 18760 21968 18766
rect 21916 18702 21968 18708
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 22020 17785 22048 18226
rect 22006 17776 22062 17785
rect 22006 17711 22062 17720
rect 22112 17678 22140 19926
rect 22204 19786 22232 21490
rect 22284 20256 22336 20262
rect 22284 20198 22336 20204
rect 22296 20058 22324 20198
rect 22388 20058 22416 21490
rect 22480 20754 22508 22170
rect 22480 20726 22600 20754
rect 22284 20052 22336 20058
rect 22284 19994 22336 20000
rect 22376 20052 22428 20058
rect 22376 19994 22428 20000
rect 22388 19854 22416 19994
rect 22376 19848 22428 19854
rect 22376 19790 22428 19796
rect 22192 19780 22244 19786
rect 22192 19722 22244 19728
rect 22100 17672 22152 17678
rect 22100 17614 22152 17620
rect 22112 17490 22140 17614
rect 22204 17610 22232 19722
rect 22572 19378 22600 20726
rect 22664 20602 22692 22578
rect 22848 21729 22876 23666
rect 22940 22642 22968 28358
rect 23124 28082 23152 30110
rect 23296 30116 23348 30122
rect 23296 30058 23348 30064
rect 23308 29050 23336 30058
rect 23400 29850 23428 30631
rect 23388 29844 23440 29850
rect 23388 29786 23440 29792
rect 23388 29640 23440 29646
rect 23388 29582 23440 29588
rect 23400 29306 23428 29582
rect 23388 29300 23440 29306
rect 23388 29242 23440 29248
rect 23400 29170 23428 29242
rect 23388 29164 23440 29170
rect 23388 29106 23440 29112
rect 23204 29028 23256 29034
rect 23308 29022 23428 29050
rect 23204 28970 23256 28976
rect 23112 28076 23164 28082
rect 23112 28018 23164 28024
rect 23018 27160 23074 27169
rect 23018 27095 23074 27104
rect 23032 26382 23060 27095
rect 23124 26926 23152 28018
rect 23112 26920 23164 26926
rect 23112 26862 23164 26868
rect 23020 26376 23072 26382
rect 23020 26318 23072 26324
rect 23032 25974 23060 26318
rect 23020 25968 23072 25974
rect 23020 25910 23072 25916
rect 23020 25152 23072 25158
rect 23020 25094 23072 25100
rect 23032 24206 23060 25094
rect 23112 24744 23164 24750
rect 23112 24686 23164 24692
rect 23020 24200 23072 24206
rect 23020 24142 23072 24148
rect 22928 22636 22980 22642
rect 22928 22578 22980 22584
rect 23020 22094 23072 22098
rect 23124 22094 23152 24686
rect 23216 23610 23244 28970
rect 23296 28960 23348 28966
rect 23296 28902 23348 28908
rect 23308 28422 23336 28902
rect 23296 28416 23348 28422
rect 23296 28358 23348 28364
rect 23294 28112 23350 28121
rect 23294 28047 23350 28056
rect 23308 27674 23336 28047
rect 23296 27668 23348 27674
rect 23296 27610 23348 27616
rect 23400 27169 23428 29022
rect 23492 28762 23520 30670
rect 23584 30394 23612 30670
rect 23572 30388 23624 30394
rect 23572 30330 23624 30336
rect 23676 30326 23704 31282
rect 23768 30734 23796 31282
rect 23756 30728 23808 30734
rect 23756 30670 23808 30676
rect 23756 30592 23808 30598
rect 23756 30534 23808 30540
rect 23664 30320 23716 30326
rect 23664 30262 23716 30268
rect 23664 29640 23716 29646
rect 23664 29582 23716 29588
rect 23572 29300 23624 29306
rect 23572 29242 23624 29248
rect 23584 29170 23612 29242
rect 23572 29164 23624 29170
rect 23572 29106 23624 29112
rect 23480 28756 23532 28762
rect 23480 28698 23532 28704
rect 23480 27464 23532 27470
rect 23478 27432 23480 27441
rect 23532 27432 23534 27441
rect 23478 27367 23534 27376
rect 23386 27160 23442 27169
rect 23386 27095 23442 27104
rect 23388 27056 23440 27062
rect 23388 26998 23440 27004
rect 23480 27056 23532 27062
rect 23480 26998 23532 27004
rect 23296 26784 23348 26790
rect 23294 26752 23296 26761
rect 23348 26752 23350 26761
rect 23294 26687 23350 26696
rect 23400 26382 23428 26998
rect 23388 26376 23440 26382
rect 23388 26318 23440 26324
rect 23492 24818 23520 26998
rect 23584 25906 23612 29106
rect 23676 29102 23704 29582
rect 23768 29170 23796 30534
rect 23756 29164 23808 29170
rect 23756 29106 23808 29112
rect 23664 29096 23716 29102
rect 23664 29038 23716 29044
rect 23662 26344 23718 26353
rect 23662 26279 23718 26288
rect 23572 25900 23624 25906
rect 23572 25842 23624 25848
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23388 24404 23440 24410
rect 23388 24346 23440 24352
rect 23400 24206 23428 24346
rect 23296 24200 23348 24206
rect 23296 24142 23348 24148
rect 23388 24200 23440 24206
rect 23388 24142 23440 24148
rect 23308 23866 23336 24142
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 23388 23860 23440 23866
rect 23388 23802 23440 23808
rect 23308 23730 23336 23802
rect 23296 23724 23348 23730
rect 23296 23666 23348 23672
rect 23400 23610 23428 23802
rect 23216 23582 23428 23610
rect 23216 23186 23244 23582
rect 23294 23488 23350 23497
rect 23294 23423 23350 23432
rect 23204 23180 23256 23186
rect 23204 23122 23256 23128
rect 23308 23066 23336 23423
rect 23020 22092 23152 22094
rect 23072 22066 23152 22092
rect 23216 23038 23336 23066
rect 23020 22034 23072 22040
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 22834 21720 22890 21729
rect 22834 21655 22890 21664
rect 22652 20596 22704 20602
rect 22652 20538 22704 20544
rect 22744 19984 22796 19990
rect 22744 19926 22796 19932
rect 22376 19372 22428 19378
rect 22376 19314 22428 19320
rect 22560 19372 22612 19378
rect 22560 19314 22612 19320
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 22284 19236 22336 19242
rect 22284 19178 22336 19184
rect 22192 17604 22244 17610
rect 22192 17546 22244 17552
rect 22112 17462 22232 17490
rect 22008 16788 22060 16794
rect 22008 16730 22060 16736
rect 21824 16584 21876 16590
rect 21824 16526 21876 16532
rect 21640 16176 21692 16182
rect 21640 16118 21692 16124
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21468 14958 21496 15438
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 21456 14952 21508 14958
rect 21456 14894 21508 14900
rect 21640 14952 21692 14958
rect 21640 14894 21692 14900
rect 21454 14512 21510 14521
rect 21454 14447 21510 14456
rect 21468 14414 21496 14447
rect 21652 14414 21680 14894
rect 21928 14414 21956 14962
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21916 14408 21968 14414
rect 21916 14350 21968 14356
rect 21364 13796 21416 13802
rect 21364 13738 21416 13744
rect 21732 13388 21784 13394
rect 21732 13330 21784 13336
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21640 13320 21692 13326
rect 21640 13262 21692 13268
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 21100 12986 21128 13126
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 21364 12844 21416 12850
rect 21364 12786 21416 12792
rect 21192 12442 21220 12786
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 21180 12436 21232 12442
rect 21180 12378 21232 12384
rect 21376 12102 21404 12786
rect 21560 12782 21588 13262
rect 21548 12776 21600 12782
rect 21548 12718 21600 12724
rect 21456 12640 21508 12646
rect 21454 12608 21456 12617
rect 21508 12608 21510 12617
rect 21454 12543 21510 12552
rect 20812 12096 20864 12102
rect 20812 12038 20864 12044
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 20824 10674 20852 12038
rect 21468 11354 21496 12543
rect 21560 12374 21588 12718
rect 21548 12368 21600 12374
rect 21548 12310 21600 12316
rect 21652 12306 21680 13262
rect 21640 12300 21692 12306
rect 21640 12242 21692 12248
rect 21640 11824 21692 11830
rect 21640 11766 21692 11772
rect 21456 11348 21508 11354
rect 21456 11290 21508 11296
rect 21468 10742 21496 11290
rect 21652 11150 21680 11766
rect 21744 11626 21772 13330
rect 21916 13252 21968 13258
rect 21916 13194 21968 13200
rect 21928 12238 21956 13194
rect 21916 12232 21968 12238
rect 21916 12174 21968 12180
rect 21732 11620 21784 11626
rect 21732 11562 21784 11568
rect 21640 11144 21692 11150
rect 21640 11086 21692 11092
rect 21456 10736 21508 10742
rect 21456 10678 21508 10684
rect 20812 10668 20864 10674
rect 20812 10610 20864 10616
rect 20720 10464 20772 10470
rect 20720 10406 20772 10412
rect 20732 8498 20760 10406
rect 20824 10062 20852 10610
rect 21468 10062 21496 10678
rect 21744 10198 21772 11562
rect 21732 10192 21784 10198
rect 21732 10134 21784 10140
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 20812 9104 20864 9110
rect 20812 9046 20864 9052
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20260 7744 20312 7750
rect 20260 7686 20312 7692
rect 20272 7410 20300 7686
rect 20548 7546 20576 7822
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20640 7410 20668 7890
rect 20824 7818 20852 9046
rect 21100 8906 21128 9522
rect 21284 8906 21312 9522
rect 21928 9042 21956 12174
rect 22020 11762 22048 16730
rect 22100 16584 22152 16590
rect 22100 16526 22152 16532
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 22008 11008 22060 11014
rect 22008 10950 22060 10956
rect 22020 10674 22048 10950
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 22112 9994 22140 16526
rect 22204 15502 22232 17462
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 22204 14414 22232 15438
rect 22192 14408 22244 14414
rect 22192 14350 22244 14356
rect 22192 13184 22244 13190
rect 22192 13126 22244 13132
rect 22204 12850 22232 13126
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22296 12238 22324 19178
rect 22284 12232 22336 12238
rect 22284 12174 22336 12180
rect 22388 10826 22416 19314
rect 22468 18760 22520 18766
rect 22468 18702 22520 18708
rect 22480 18086 22508 18702
rect 22560 18624 22612 18630
rect 22560 18566 22612 18572
rect 22572 18465 22600 18566
rect 22558 18456 22614 18465
rect 22558 18391 22614 18400
rect 22560 18284 22612 18290
rect 22560 18226 22612 18232
rect 22468 18080 22520 18086
rect 22468 18022 22520 18028
rect 22468 17060 22520 17066
rect 22468 17002 22520 17008
rect 22480 16590 22508 17002
rect 22468 16584 22520 16590
rect 22468 16526 22520 16532
rect 22480 16182 22508 16526
rect 22468 16176 22520 16182
rect 22468 16118 22520 16124
rect 22572 16114 22600 18226
rect 22664 17921 22692 19314
rect 22650 17912 22706 17921
rect 22650 17847 22706 17856
rect 22652 17740 22704 17746
rect 22652 17682 22704 17688
rect 22664 16726 22692 17682
rect 22652 16720 22704 16726
rect 22652 16662 22704 16668
rect 22560 16108 22612 16114
rect 22560 16050 22612 16056
rect 22468 15496 22520 15502
rect 22468 15438 22520 15444
rect 22756 15450 22784 19926
rect 22848 19242 22876 21655
rect 22940 20602 22968 21966
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 22836 19236 22888 19242
rect 22836 19178 22888 19184
rect 22928 17264 22980 17270
rect 22928 17206 22980 17212
rect 22836 17128 22888 17134
rect 22836 17070 22888 17076
rect 22848 16794 22876 17070
rect 22836 16788 22888 16794
rect 22836 16730 22888 16736
rect 22848 15570 22876 16730
rect 22940 16590 22968 17206
rect 23032 17202 23060 22034
rect 23216 19854 23244 23038
rect 23492 22681 23520 24754
rect 23572 24744 23624 24750
rect 23572 24686 23624 24692
rect 23584 24342 23612 24686
rect 23572 24336 23624 24342
rect 23572 24278 23624 24284
rect 23676 23594 23704 26279
rect 23860 26042 23888 32846
rect 24044 32337 24072 33390
rect 24216 32768 24268 32774
rect 24216 32710 24268 32716
rect 24228 32434 24256 32710
rect 24124 32428 24176 32434
rect 24124 32370 24176 32376
rect 24216 32428 24268 32434
rect 24216 32370 24268 32376
rect 24030 32328 24086 32337
rect 24030 32263 24086 32272
rect 24044 29306 24072 32263
rect 24136 32026 24164 32370
rect 24124 32020 24176 32026
rect 24124 31962 24176 31968
rect 24228 30258 24256 32370
rect 24320 32314 24348 36654
rect 25688 36576 25740 36582
rect 25688 36518 25740 36524
rect 24860 36304 24912 36310
rect 24860 36246 24912 36252
rect 24676 36168 24728 36174
rect 24676 36110 24728 36116
rect 24688 35494 24716 36110
rect 24872 35630 24900 36246
rect 24952 36236 25004 36242
rect 24952 36178 25004 36184
rect 24964 35698 24992 36178
rect 24952 35692 25004 35698
rect 24952 35634 25004 35640
rect 24860 35624 24912 35630
rect 24860 35566 24912 35572
rect 24676 35488 24728 35494
rect 24676 35430 24728 35436
rect 24872 35290 24900 35566
rect 24860 35284 24912 35290
rect 24860 35226 24912 35232
rect 24676 34944 24728 34950
rect 24676 34886 24728 34892
rect 24688 34610 24716 34886
rect 24872 34762 24900 35226
rect 24964 35086 24992 35634
rect 25412 35624 25464 35630
rect 25412 35566 25464 35572
rect 24952 35080 25004 35086
rect 24952 35022 25004 35028
rect 25042 35048 25098 35057
rect 24780 34734 24900 34762
rect 24676 34604 24728 34610
rect 24676 34546 24728 34552
rect 24320 32286 24624 32314
rect 24596 31754 24624 32286
rect 24412 31726 24624 31754
rect 24308 31204 24360 31210
rect 24308 31146 24360 31152
rect 24216 30252 24268 30258
rect 24216 30194 24268 30200
rect 24320 30054 24348 31146
rect 24308 30048 24360 30054
rect 24308 29990 24360 29996
rect 24124 29708 24176 29714
rect 24124 29650 24176 29656
rect 24032 29300 24084 29306
rect 24032 29242 24084 29248
rect 24136 28490 24164 29650
rect 24320 29345 24348 29990
rect 24306 29336 24362 29345
rect 24306 29271 24362 29280
rect 24124 28484 24176 28490
rect 24124 28426 24176 28432
rect 24032 27940 24084 27946
rect 24136 27928 24164 28426
rect 24308 28144 24360 28150
rect 24308 28086 24360 28092
rect 24084 27900 24164 27928
rect 24032 27882 24084 27888
rect 24044 27062 24072 27882
rect 24124 27532 24176 27538
rect 24124 27474 24176 27480
rect 24032 27056 24084 27062
rect 24032 26998 24084 27004
rect 24032 26240 24084 26246
rect 24032 26182 24084 26188
rect 23848 26036 23900 26042
rect 23848 25978 23900 25984
rect 23940 24812 23992 24818
rect 23940 24754 23992 24760
rect 23754 24712 23810 24721
rect 23754 24647 23810 24656
rect 23768 23730 23796 24647
rect 23952 24410 23980 24754
rect 23940 24404 23992 24410
rect 23940 24346 23992 24352
rect 24044 24206 24072 26182
rect 24136 24886 24164 27474
rect 24320 26994 24348 28086
rect 24308 26988 24360 26994
rect 24308 26930 24360 26936
rect 24124 24880 24176 24886
rect 24124 24822 24176 24828
rect 24032 24200 24084 24206
rect 24032 24142 24084 24148
rect 24044 23798 24072 24142
rect 24032 23792 24084 23798
rect 24032 23734 24084 23740
rect 23756 23724 23808 23730
rect 23756 23666 23808 23672
rect 23664 23588 23716 23594
rect 23664 23530 23716 23536
rect 23478 22672 23534 22681
rect 23676 22642 23704 23530
rect 23478 22607 23534 22616
rect 23664 22636 23716 22642
rect 23388 22568 23440 22574
rect 23388 22510 23440 22516
rect 23400 22094 23428 22510
rect 23308 22066 23428 22094
rect 23204 19848 23256 19854
rect 23204 19790 23256 19796
rect 23204 18080 23256 18086
rect 23204 18022 23256 18028
rect 23112 17740 23164 17746
rect 23112 17682 23164 17688
rect 23124 17542 23152 17682
rect 23216 17678 23244 18022
rect 23204 17672 23256 17678
rect 23204 17614 23256 17620
rect 23112 17536 23164 17542
rect 23112 17478 23164 17484
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 23020 17196 23072 17202
rect 23020 17138 23072 17144
rect 23124 16998 23152 17274
rect 23216 17270 23244 17614
rect 23204 17264 23256 17270
rect 23204 17206 23256 17212
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 22928 16584 22980 16590
rect 22928 16526 22980 16532
rect 23112 16584 23164 16590
rect 23112 16526 23164 16532
rect 22940 16454 22968 16526
rect 22928 16448 22980 16454
rect 22928 16390 22980 16396
rect 22940 15910 22968 16390
rect 23020 16176 23072 16182
rect 23020 16118 23072 16124
rect 22928 15904 22980 15910
rect 22928 15846 22980 15852
rect 22836 15564 22888 15570
rect 22836 15506 22888 15512
rect 23032 15502 23060 16118
rect 23020 15496 23072 15502
rect 22480 15026 22508 15438
rect 22756 15422 22968 15450
rect 23020 15438 23072 15444
rect 22468 15020 22520 15026
rect 22468 14962 22520 14968
rect 22560 15020 22612 15026
rect 22560 14962 22612 14968
rect 22572 14278 22600 14962
rect 22744 14476 22796 14482
rect 22744 14418 22796 14424
rect 22560 14272 22612 14278
rect 22560 14214 22612 14220
rect 22756 14074 22784 14418
rect 22744 14068 22796 14074
rect 22744 14010 22796 14016
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 22756 13258 22784 13806
rect 22836 13728 22888 13734
rect 22836 13670 22888 13676
rect 22744 13252 22796 13258
rect 22744 13194 22796 13200
rect 22468 13184 22520 13190
rect 22468 13126 22520 13132
rect 22480 12782 22508 13126
rect 22468 12776 22520 12782
rect 22468 12718 22520 12724
rect 22468 11212 22520 11218
rect 22468 11154 22520 11160
rect 22296 10798 22416 10826
rect 22192 10668 22244 10674
rect 22192 10610 22244 10616
rect 22204 10266 22232 10610
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 22100 9988 22152 9994
rect 22100 9930 22152 9936
rect 22296 9586 22324 10798
rect 22376 10668 22428 10674
rect 22376 10610 22428 10616
rect 22388 10198 22416 10610
rect 22376 10192 22428 10198
rect 22376 10134 22428 10140
rect 22480 10062 22508 11154
rect 22652 10464 22704 10470
rect 22652 10406 22704 10412
rect 22664 10062 22692 10406
rect 22468 10056 22520 10062
rect 22468 9998 22520 10004
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22284 9580 22336 9586
rect 22284 9522 22336 9528
rect 22480 9518 22508 9998
rect 22468 9512 22520 9518
rect 22468 9454 22520 9460
rect 22560 9444 22612 9450
rect 22560 9386 22612 9392
rect 21916 9036 21968 9042
rect 21916 8978 21968 8984
rect 21088 8900 21140 8906
rect 21088 8842 21140 8848
rect 21272 8900 21324 8906
rect 21272 8842 21324 8848
rect 20904 8424 20956 8430
rect 20904 8366 20956 8372
rect 20916 8090 20944 8366
rect 20904 8084 20956 8090
rect 20904 8026 20956 8032
rect 20812 7812 20864 7818
rect 20812 7754 20864 7760
rect 20824 7478 20852 7754
rect 20812 7472 20864 7478
rect 20812 7414 20864 7420
rect 20916 7410 20944 8026
rect 22468 7880 22520 7886
rect 22468 7822 22520 7828
rect 21732 7812 21784 7818
rect 21732 7754 21784 7760
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 20088 6798 20116 7142
rect 21744 7002 21772 7754
rect 21732 6996 21784 7002
rect 21732 6938 21784 6944
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 19984 6792 20036 6798
rect 19984 6734 20036 6740
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19996 6390 20024 6734
rect 20456 6458 20484 6802
rect 22480 6798 22508 7822
rect 22572 7546 22600 9386
rect 22560 7540 22612 7546
rect 22560 7482 22612 7488
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 22468 6792 22520 6798
rect 22468 6734 22520 6740
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 19984 6384 20036 6390
rect 19984 6326 20036 6332
rect 20548 6118 20576 6734
rect 21364 6656 21416 6662
rect 21364 6598 21416 6604
rect 21376 6322 21404 6598
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 20536 6112 20588 6118
rect 20536 6054 20588 6060
rect 21180 6112 21232 6118
rect 21180 6054 21232 6060
rect 21192 5710 21220 6054
rect 22100 5772 22152 5778
rect 22100 5714 22152 5720
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 22112 5234 22140 5714
rect 22848 5370 22876 13670
rect 22940 11218 22968 15422
rect 22928 11212 22980 11218
rect 22928 11154 22980 11160
rect 23032 8090 23060 15438
rect 23124 14346 23152 16526
rect 23112 14340 23164 14346
rect 23112 14282 23164 14288
rect 23204 14340 23256 14346
rect 23204 14282 23256 14288
rect 23216 13938 23244 14282
rect 23204 13932 23256 13938
rect 23204 13874 23256 13880
rect 23308 13462 23336 22066
rect 23388 20596 23440 20602
rect 23388 20538 23440 20544
rect 23400 19378 23428 20538
rect 23492 19446 23520 22607
rect 23664 22578 23716 22584
rect 24136 22030 24164 24822
rect 24320 22166 24348 26930
rect 24412 22710 24440 31726
rect 24688 30054 24716 34546
rect 24780 33998 24808 34734
rect 24964 34626 24992 35022
rect 25042 34983 25098 34992
rect 25136 35012 25188 35018
rect 24872 34598 24992 34626
rect 24768 33992 24820 33998
rect 24768 33934 24820 33940
rect 24780 33522 24808 33934
rect 24768 33516 24820 33522
rect 24768 33458 24820 33464
rect 24780 32774 24808 33458
rect 24872 33386 24900 34598
rect 25056 33998 25084 34983
rect 25136 34954 25188 34960
rect 25148 34406 25176 34954
rect 25136 34400 25188 34406
rect 25136 34342 25188 34348
rect 25044 33992 25096 33998
rect 25044 33934 25096 33940
rect 24860 33380 24912 33386
rect 24860 33322 24912 33328
rect 24768 32768 24820 32774
rect 24768 32710 24820 32716
rect 24872 31822 24900 33322
rect 24952 32972 25004 32978
rect 24952 32914 25004 32920
rect 24860 31816 24912 31822
rect 24860 31758 24912 31764
rect 24858 30832 24914 30841
rect 24858 30767 24914 30776
rect 24872 30734 24900 30767
rect 24860 30728 24912 30734
rect 24860 30670 24912 30676
rect 24768 30320 24820 30326
rect 24768 30262 24820 30268
rect 24676 30048 24728 30054
rect 24676 29990 24728 29996
rect 24780 29510 24808 30262
rect 24860 30252 24912 30258
rect 24860 30194 24912 30200
rect 24676 29504 24728 29510
rect 24676 29446 24728 29452
rect 24768 29504 24820 29510
rect 24768 29446 24820 29452
rect 24688 28558 24716 29446
rect 24780 29170 24808 29446
rect 24768 29164 24820 29170
rect 24768 29106 24820 29112
rect 24872 28762 24900 30194
rect 24964 29306 24992 32914
rect 25056 32434 25084 33934
rect 25148 33590 25176 34342
rect 25424 34202 25452 35566
rect 25700 34610 25728 36518
rect 26252 35630 26280 37198
rect 26424 36780 26476 36786
rect 26424 36722 26476 36728
rect 26332 36168 26384 36174
rect 26332 36110 26384 36116
rect 26240 35624 26292 35630
rect 26240 35566 26292 35572
rect 26344 35562 26372 36110
rect 26436 35766 26464 36722
rect 26424 35760 26476 35766
rect 26424 35702 26476 35708
rect 26528 35698 26556 37266
rect 27436 37256 27488 37262
rect 27436 37198 27488 37204
rect 27068 36712 27120 36718
rect 27068 36654 27120 36660
rect 27080 36310 27108 36654
rect 27448 36378 27476 37198
rect 27620 36848 27672 36854
rect 27620 36790 27672 36796
rect 27436 36372 27488 36378
rect 27436 36314 27488 36320
rect 27068 36304 27120 36310
rect 27068 36246 27120 36252
rect 27632 36242 27660 36790
rect 27620 36236 27672 36242
rect 27620 36178 27672 36184
rect 27528 36100 27580 36106
rect 27528 36042 27580 36048
rect 26792 36032 26844 36038
rect 26792 35974 26844 35980
rect 26516 35692 26568 35698
rect 26516 35634 26568 35640
rect 26332 35556 26384 35562
rect 26332 35498 26384 35504
rect 26424 35488 26476 35494
rect 26424 35430 26476 35436
rect 25688 34604 25740 34610
rect 25688 34546 25740 34552
rect 25412 34196 25464 34202
rect 25412 34138 25464 34144
rect 25596 33924 25648 33930
rect 25596 33866 25648 33872
rect 25136 33584 25188 33590
rect 25136 33526 25188 33532
rect 25228 33108 25280 33114
rect 25228 33050 25280 33056
rect 25240 32473 25268 33050
rect 25226 32464 25282 32473
rect 25044 32428 25096 32434
rect 25226 32399 25282 32408
rect 25044 32370 25096 32376
rect 25320 32020 25372 32026
rect 25320 31962 25372 31968
rect 25044 31680 25096 31686
rect 25044 31622 25096 31628
rect 25056 30938 25084 31622
rect 25228 31272 25280 31278
rect 25228 31214 25280 31220
rect 25044 30932 25096 30938
rect 25044 30874 25096 30880
rect 25056 29646 25084 30874
rect 25136 30728 25188 30734
rect 25136 30670 25188 30676
rect 25044 29640 25096 29646
rect 25044 29582 25096 29588
rect 24952 29300 25004 29306
rect 24952 29242 25004 29248
rect 25148 29209 25176 30670
rect 25240 30190 25268 31214
rect 25228 30184 25280 30190
rect 25228 30126 25280 30132
rect 25226 29336 25282 29345
rect 25226 29271 25282 29280
rect 25240 29238 25268 29271
rect 25228 29232 25280 29238
rect 25134 29200 25190 29209
rect 25228 29174 25280 29180
rect 25134 29135 25190 29144
rect 25332 29152 25360 31962
rect 25504 31884 25556 31890
rect 25504 31826 25556 31832
rect 25412 31748 25464 31754
rect 25412 31690 25464 31696
rect 25424 31346 25452 31690
rect 25412 31340 25464 31346
rect 25412 31282 25464 31288
rect 25412 31136 25464 31142
rect 25412 31078 25464 31084
rect 25424 30870 25452 31078
rect 25412 30864 25464 30870
rect 25412 30806 25464 30812
rect 25516 30734 25544 31826
rect 25608 31822 25636 33866
rect 25700 33862 25728 34546
rect 25872 34536 25924 34542
rect 25872 34478 25924 34484
rect 25780 34196 25832 34202
rect 25780 34138 25832 34144
rect 25688 33856 25740 33862
rect 25688 33798 25740 33804
rect 25700 32842 25728 33798
rect 25792 33318 25820 34138
rect 25884 34066 25912 34478
rect 25872 34060 25924 34066
rect 25872 34002 25924 34008
rect 25780 33312 25832 33318
rect 25780 33254 25832 33260
rect 25688 32836 25740 32842
rect 25688 32778 25740 32784
rect 25700 32434 25728 32778
rect 25688 32428 25740 32434
rect 25688 32370 25740 32376
rect 25688 32224 25740 32230
rect 25688 32166 25740 32172
rect 25596 31816 25648 31822
rect 25700 31793 25728 32166
rect 25792 31822 25820 33254
rect 25780 31816 25832 31822
rect 25596 31758 25648 31764
rect 25686 31784 25742 31793
rect 25780 31758 25832 31764
rect 25686 31719 25742 31728
rect 25596 31476 25648 31482
rect 25596 31418 25648 31424
rect 25608 31346 25636 31418
rect 25596 31340 25648 31346
rect 25596 31282 25648 31288
rect 25504 30728 25556 30734
rect 25504 30670 25556 30676
rect 25504 30048 25556 30054
rect 25504 29990 25556 29996
rect 25516 29889 25544 29990
rect 25502 29880 25558 29889
rect 25502 29815 25558 29824
rect 25504 29640 25556 29646
rect 25504 29582 25556 29588
rect 25412 29164 25464 29170
rect 25332 29124 25412 29152
rect 25228 29096 25280 29102
rect 25228 29038 25280 29044
rect 24860 28756 24912 28762
rect 24860 28698 24912 28704
rect 24676 28552 24728 28558
rect 24676 28494 24728 28500
rect 24688 28082 24716 28494
rect 24952 28416 25004 28422
rect 24952 28358 25004 28364
rect 24860 28144 24912 28150
rect 24860 28086 24912 28092
rect 24676 28076 24728 28082
rect 24676 28018 24728 28024
rect 24676 27940 24728 27946
rect 24676 27882 24728 27888
rect 24492 27396 24544 27402
rect 24492 27338 24544 27344
rect 24504 26024 24532 27338
rect 24688 27130 24716 27882
rect 24872 27656 24900 28086
rect 24780 27628 24900 27656
rect 24676 27124 24728 27130
rect 24676 27066 24728 27072
rect 24584 26784 24636 26790
rect 24584 26726 24636 26732
rect 24596 26382 24624 26726
rect 24676 26444 24728 26450
rect 24676 26386 24728 26392
rect 24584 26376 24636 26382
rect 24584 26318 24636 26324
rect 24584 26036 24636 26042
rect 24504 25996 24584 26024
rect 24584 25978 24636 25984
rect 24490 25936 24546 25945
rect 24490 25871 24492 25880
rect 24544 25871 24546 25880
rect 24492 25842 24544 25848
rect 24584 25764 24636 25770
rect 24584 25706 24636 25712
rect 24596 25158 24624 25706
rect 24688 25537 24716 26386
rect 24674 25528 24730 25537
rect 24674 25463 24730 25472
rect 24780 25430 24808 27628
rect 24964 27441 24992 28358
rect 25240 28150 25268 29038
rect 25332 28966 25360 29124
rect 25412 29106 25464 29112
rect 25320 28960 25372 28966
rect 25320 28902 25372 28908
rect 25228 28144 25280 28150
rect 25228 28086 25280 28092
rect 24950 27432 25006 27441
rect 24950 27367 25006 27376
rect 24964 26382 24992 27367
rect 25134 26888 25190 26897
rect 25134 26823 25190 26832
rect 25148 26382 25176 26823
rect 24952 26376 25004 26382
rect 24952 26318 25004 26324
rect 25136 26376 25188 26382
rect 25332 26330 25360 28902
rect 25516 28082 25544 29582
rect 25504 28076 25556 28082
rect 25504 28018 25556 28024
rect 25516 27470 25544 28018
rect 25608 27538 25636 31282
rect 25700 30666 25728 31719
rect 25688 30660 25740 30666
rect 25688 30602 25740 30608
rect 25596 27532 25648 27538
rect 25596 27474 25648 27480
rect 25504 27464 25556 27470
rect 25700 27452 25728 30602
rect 25792 30410 25820 31758
rect 25884 31686 25912 34002
rect 26436 33522 26464 35430
rect 26700 34128 26752 34134
rect 26700 34070 26752 34076
rect 26516 33856 26568 33862
rect 26516 33798 26568 33804
rect 26240 33516 26292 33522
rect 26240 33458 26292 33464
rect 26424 33516 26476 33522
rect 26424 33458 26476 33464
rect 26252 33046 26280 33458
rect 26240 33040 26292 33046
rect 26240 32982 26292 32988
rect 25964 32904 26016 32910
rect 25964 32846 26016 32852
rect 26240 32904 26292 32910
rect 26240 32846 26292 32852
rect 25976 32586 26004 32846
rect 25976 32570 26188 32586
rect 25964 32564 26188 32570
rect 26016 32558 26188 32564
rect 25964 32506 26016 32512
rect 26160 32502 26188 32558
rect 26148 32496 26200 32502
rect 26148 32438 26200 32444
rect 26252 32434 26280 32846
rect 26240 32428 26292 32434
rect 26240 32370 26292 32376
rect 26252 32337 26280 32370
rect 26238 32328 26294 32337
rect 26238 32263 26294 32272
rect 26436 31754 26464 33458
rect 26240 31748 26292 31754
rect 26240 31690 26292 31696
rect 26424 31748 26476 31754
rect 26424 31690 26476 31696
rect 25872 31680 25924 31686
rect 25872 31622 25924 31628
rect 26056 31680 26108 31686
rect 26056 31622 26108 31628
rect 25872 31340 25924 31346
rect 25872 31282 25924 31288
rect 25884 30870 25912 31282
rect 25964 31204 26016 31210
rect 25964 31146 26016 31152
rect 25872 30864 25924 30870
rect 25872 30806 25924 30812
rect 25976 30734 26004 31146
rect 26068 31142 26096 31622
rect 26056 31136 26108 31142
rect 26056 31078 26108 31084
rect 25964 30728 26016 30734
rect 25964 30670 26016 30676
rect 26252 30546 26280 31690
rect 26424 31204 26476 31210
rect 26424 31146 26476 31152
rect 26436 30841 26464 31146
rect 26422 30832 26478 30841
rect 26422 30767 26478 30776
rect 26528 30682 26556 33798
rect 26436 30654 26556 30682
rect 26252 30518 26372 30546
rect 25792 30382 25912 30410
rect 25780 30252 25832 30258
rect 25780 30194 25832 30200
rect 25792 28218 25820 30194
rect 25884 29102 25912 30382
rect 26240 30388 26292 30394
rect 26240 30330 26292 30336
rect 26252 30258 26280 30330
rect 26240 30252 26292 30258
rect 26240 30194 26292 30200
rect 26056 29844 26108 29850
rect 26056 29786 26108 29792
rect 25964 29504 26016 29510
rect 25964 29446 26016 29452
rect 25976 29306 26004 29446
rect 25964 29300 26016 29306
rect 25964 29242 26016 29248
rect 25964 29164 26016 29170
rect 25964 29106 26016 29112
rect 25872 29096 25924 29102
rect 25872 29038 25924 29044
rect 25884 28626 25912 29038
rect 25976 28762 26004 29106
rect 25964 28756 26016 28762
rect 25964 28698 26016 28704
rect 25872 28620 25924 28626
rect 25872 28562 25924 28568
rect 25780 28212 25832 28218
rect 25780 28154 25832 28160
rect 25964 27940 26016 27946
rect 25964 27882 26016 27888
rect 25872 27600 25924 27606
rect 25872 27542 25924 27548
rect 25884 27452 25912 27542
rect 25700 27424 25912 27452
rect 25504 27406 25556 27412
rect 25780 27328 25832 27334
rect 25780 27270 25832 27276
rect 25596 27124 25648 27130
rect 25596 27066 25648 27072
rect 25412 26988 25464 26994
rect 25412 26930 25464 26936
rect 25136 26318 25188 26324
rect 24858 25800 24914 25809
rect 24858 25735 24860 25744
rect 24912 25735 24914 25744
rect 24860 25706 24912 25712
rect 24768 25424 24820 25430
rect 24768 25366 24820 25372
rect 24860 25424 24912 25430
rect 24860 25366 24912 25372
rect 24872 25276 24900 25366
rect 24964 25294 24992 26318
rect 25240 26302 25360 26330
rect 25044 25968 25096 25974
rect 25044 25910 25096 25916
rect 24780 25248 24900 25276
rect 24952 25288 25004 25294
rect 24584 25152 24636 25158
rect 24584 25094 24636 25100
rect 24584 24404 24636 24410
rect 24584 24346 24636 24352
rect 24492 22976 24544 22982
rect 24492 22918 24544 22924
rect 24400 22704 24452 22710
rect 24400 22646 24452 22652
rect 24504 22642 24532 22918
rect 24492 22636 24544 22642
rect 24492 22578 24544 22584
rect 24308 22160 24360 22166
rect 24308 22102 24360 22108
rect 24124 22024 24176 22030
rect 24124 21966 24176 21972
rect 24136 21010 24164 21966
rect 24596 21690 24624 24346
rect 24780 24206 24808 25248
rect 24952 25230 25004 25236
rect 24768 24200 24820 24206
rect 24768 24142 24820 24148
rect 24780 23118 24808 24142
rect 24952 24132 25004 24138
rect 24952 24074 25004 24080
rect 24964 23730 24992 24074
rect 24952 23724 25004 23730
rect 24952 23666 25004 23672
rect 24768 23112 24820 23118
rect 24768 23054 24820 23060
rect 24964 22030 24992 23666
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 24676 21888 24728 21894
rect 24676 21830 24728 21836
rect 24952 21888 25004 21894
rect 24952 21830 25004 21836
rect 24584 21684 24636 21690
rect 24584 21626 24636 21632
rect 24596 21536 24624 21626
rect 24688 21554 24716 21830
rect 24504 21508 24624 21536
rect 24676 21548 24728 21554
rect 24124 21004 24176 21010
rect 24124 20946 24176 20952
rect 24504 20942 24532 21508
rect 24676 21490 24728 21496
rect 24584 21412 24636 21418
rect 24584 21354 24636 21360
rect 24492 20936 24544 20942
rect 24492 20878 24544 20884
rect 24032 20460 24084 20466
rect 24032 20402 24084 20408
rect 23848 20392 23900 20398
rect 24044 20369 24072 20402
rect 23848 20334 23900 20340
rect 24030 20360 24086 20369
rect 23480 19440 23532 19446
rect 23480 19382 23532 19388
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 23388 19236 23440 19242
rect 23388 19178 23440 19184
rect 23400 18426 23428 19178
rect 23480 18828 23532 18834
rect 23480 18770 23532 18776
rect 23388 18420 23440 18426
rect 23388 18362 23440 18368
rect 23400 13734 23428 18362
rect 23492 18290 23520 18770
rect 23860 18766 23888 20334
rect 24030 20295 24086 20304
rect 23940 19984 23992 19990
rect 23940 19926 23992 19932
rect 23952 19825 23980 19926
rect 23938 19816 23994 19825
rect 23938 19751 23994 19760
rect 24596 19718 24624 21354
rect 24584 19712 24636 19718
rect 24584 19654 24636 19660
rect 24306 19408 24362 19417
rect 24306 19343 24308 19352
rect 24360 19343 24362 19352
rect 24308 19314 24360 19320
rect 24492 19168 24544 19174
rect 24492 19110 24544 19116
rect 24504 18970 24532 19110
rect 24032 18964 24084 18970
rect 24032 18906 24084 18912
rect 24492 18964 24544 18970
rect 24492 18906 24544 18912
rect 23940 18828 23992 18834
rect 23940 18770 23992 18776
rect 23848 18760 23900 18766
rect 23848 18702 23900 18708
rect 23480 18284 23532 18290
rect 23480 18226 23532 18232
rect 23572 18216 23624 18222
rect 23572 18158 23624 18164
rect 23584 17678 23612 18158
rect 23756 18148 23808 18154
rect 23756 18090 23808 18096
rect 23664 18080 23716 18086
rect 23664 18022 23716 18028
rect 23572 17672 23624 17678
rect 23572 17614 23624 17620
rect 23676 15026 23704 18022
rect 23768 17610 23796 18090
rect 23756 17604 23808 17610
rect 23756 17546 23808 17552
rect 23860 17338 23888 18702
rect 23952 18358 23980 18770
rect 23940 18352 23992 18358
rect 23940 18294 23992 18300
rect 23952 17678 23980 18294
rect 24044 18290 24072 18906
rect 24688 18358 24716 21490
rect 24768 21004 24820 21010
rect 24768 20946 24820 20952
rect 24780 20806 24808 20946
rect 24768 20800 24820 20806
rect 24964 20754 24992 21830
rect 25056 21146 25084 25910
rect 25240 25294 25268 26302
rect 25320 26240 25372 26246
rect 25320 26182 25372 26188
rect 25228 25288 25280 25294
rect 25228 25230 25280 25236
rect 25240 24818 25268 25230
rect 25332 24954 25360 26182
rect 25424 25838 25452 26930
rect 25412 25832 25464 25838
rect 25412 25774 25464 25780
rect 25412 25356 25464 25362
rect 25412 25298 25464 25304
rect 25320 24948 25372 24954
rect 25320 24890 25372 24896
rect 25228 24812 25280 24818
rect 25228 24754 25280 24760
rect 25424 23186 25452 25298
rect 25504 25220 25556 25226
rect 25504 25162 25556 25168
rect 25516 24818 25544 25162
rect 25608 24886 25636 27066
rect 25792 27062 25820 27270
rect 25780 27056 25832 27062
rect 25700 27016 25780 27044
rect 25700 25362 25728 27016
rect 25780 26998 25832 27004
rect 25778 26480 25834 26489
rect 25884 26466 25912 27424
rect 25976 26926 26004 27882
rect 25964 26920 26016 26926
rect 25964 26862 26016 26868
rect 25834 26438 25912 26466
rect 25778 26415 25834 26424
rect 25792 26314 25820 26415
rect 25780 26308 25832 26314
rect 25780 26250 25832 26256
rect 25964 26308 26016 26314
rect 25964 26250 26016 26256
rect 25976 25945 26004 26250
rect 25962 25936 26018 25945
rect 25962 25871 26018 25880
rect 25688 25356 25740 25362
rect 25688 25298 25740 25304
rect 25872 25356 25924 25362
rect 25872 25298 25924 25304
rect 25596 24880 25648 24886
rect 25596 24822 25648 24828
rect 25504 24812 25556 24818
rect 25504 24754 25556 24760
rect 25688 24744 25740 24750
rect 25688 24686 25740 24692
rect 25700 24449 25728 24686
rect 25686 24440 25742 24449
rect 25686 24375 25742 24384
rect 25504 24064 25556 24070
rect 25504 24006 25556 24012
rect 25412 23180 25464 23186
rect 25412 23122 25464 23128
rect 25320 22704 25372 22710
rect 25320 22646 25372 22652
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 25228 22024 25280 22030
rect 25228 21966 25280 21972
rect 25148 21350 25176 21966
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 25044 21140 25096 21146
rect 25044 21082 25096 21088
rect 25148 20754 25176 21286
rect 25240 20806 25268 21966
rect 25332 21146 25360 22646
rect 25320 21140 25372 21146
rect 25320 21082 25372 21088
rect 25320 20936 25372 20942
rect 25320 20878 25372 20884
rect 25412 20936 25464 20942
rect 25412 20878 25464 20884
rect 24768 20742 24820 20748
rect 24872 20726 24992 20754
rect 25056 20726 25176 20754
rect 25228 20800 25280 20806
rect 25228 20742 25280 20748
rect 24768 20324 24820 20330
rect 24768 20266 24820 20272
rect 24780 19854 24808 20266
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24676 18352 24728 18358
rect 24676 18294 24728 18300
rect 24032 18284 24084 18290
rect 24032 18226 24084 18232
rect 24044 17882 24072 18226
rect 24124 18216 24176 18222
rect 24124 18158 24176 18164
rect 24032 17876 24084 17882
rect 24032 17818 24084 17824
rect 23940 17672 23992 17678
rect 23940 17614 23992 17620
rect 23848 17332 23900 17338
rect 23848 17274 23900 17280
rect 23952 17066 23980 17614
rect 24044 17134 24072 17818
rect 24136 17746 24164 18158
rect 24124 17740 24176 17746
rect 24124 17682 24176 17688
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24136 17542 24164 17682
rect 24124 17536 24176 17542
rect 24124 17478 24176 17484
rect 24584 17536 24636 17542
rect 24688 17513 24716 17682
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24584 17478 24636 17484
rect 24674 17504 24730 17513
rect 24596 17202 24624 17478
rect 24674 17439 24730 17448
rect 24584 17196 24636 17202
rect 24584 17138 24636 17144
rect 24780 17134 24808 17614
rect 24032 17128 24084 17134
rect 24032 17070 24084 17076
rect 24768 17128 24820 17134
rect 24768 17070 24820 17076
rect 23940 17060 23992 17066
rect 23940 17002 23992 17008
rect 23940 16788 23992 16794
rect 23940 16730 23992 16736
rect 23664 15020 23716 15026
rect 23664 14962 23716 14968
rect 23572 14408 23624 14414
rect 23572 14350 23624 14356
rect 23480 13864 23532 13870
rect 23480 13806 23532 13812
rect 23388 13728 23440 13734
rect 23388 13670 23440 13676
rect 23296 13456 23348 13462
rect 23296 13398 23348 13404
rect 23492 13326 23520 13806
rect 23584 13530 23612 14350
rect 23572 13524 23624 13530
rect 23572 13466 23624 13472
rect 23480 13320 23532 13326
rect 23480 13262 23532 13268
rect 23480 11824 23532 11830
rect 23480 11766 23532 11772
rect 23492 10606 23520 11766
rect 23480 10600 23532 10606
rect 23480 10542 23532 10548
rect 23492 9654 23520 10542
rect 23480 9648 23532 9654
rect 23480 9590 23532 9596
rect 23492 8498 23520 9590
rect 23480 8492 23532 8498
rect 23480 8434 23532 8440
rect 23020 8084 23072 8090
rect 23020 8026 23072 8032
rect 23204 6792 23256 6798
rect 23204 6734 23256 6740
rect 22836 5364 22888 5370
rect 22836 5306 22888 5312
rect 23216 5302 23244 6734
rect 23296 6724 23348 6730
rect 23296 6666 23348 6672
rect 23308 6458 23336 6666
rect 23296 6452 23348 6458
rect 23296 6394 23348 6400
rect 23480 5364 23532 5370
rect 23480 5306 23532 5312
rect 23204 5296 23256 5302
rect 23204 5238 23256 5244
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 23020 5228 23072 5234
rect 23020 5170 23072 5176
rect 23032 4826 23060 5170
rect 23216 5166 23244 5238
rect 23204 5160 23256 5166
rect 23204 5102 23256 5108
rect 23020 4820 23072 4826
rect 23020 4762 23072 4768
rect 23492 4622 23520 5306
rect 23676 4758 23704 14962
rect 23952 14890 23980 16730
rect 24216 15564 24268 15570
rect 24216 15506 24268 15512
rect 24228 15026 24256 15506
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 23940 14884 23992 14890
rect 23940 14826 23992 14832
rect 23952 14482 23980 14826
rect 24412 14822 24440 15438
rect 24584 15020 24636 15026
rect 24584 14962 24636 14968
rect 24124 14816 24176 14822
rect 24124 14758 24176 14764
rect 24400 14816 24452 14822
rect 24400 14758 24452 14764
rect 24136 14482 24164 14758
rect 24412 14550 24440 14758
rect 24400 14544 24452 14550
rect 24400 14486 24452 14492
rect 23940 14476 23992 14482
rect 23940 14418 23992 14424
rect 24124 14476 24176 14482
rect 24124 14418 24176 14424
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23860 6390 23888 14214
rect 23940 14000 23992 14006
rect 23940 13942 23992 13948
rect 23952 13326 23980 13942
rect 24136 13870 24164 14418
rect 24596 14414 24624 14962
rect 24584 14408 24636 14414
rect 24584 14350 24636 14356
rect 24216 14272 24268 14278
rect 24216 14214 24268 14220
rect 24228 13938 24256 14214
rect 24596 13938 24624 14350
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 24124 13864 24176 13870
rect 24124 13806 24176 13812
rect 23940 13320 23992 13326
rect 23940 13262 23992 13268
rect 24228 13258 24256 13874
rect 24216 13252 24268 13258
rect 24216 13194 24268 13200
rect 24872 12434 24900 20726
rect 25056 20466 25084 20726
rect 25044 20460 25096 20466
rect 25044 20402 25096 20408
rect 25136 20460 25188 20466
rect 25136 20402 25188 20408
rect 24952 19372 25004 19378
rect 24952 19314 25004 19320
rect 24964 18970 24992 19314
rect 25056 19310 25084 20402
rect 25148 19854 25176 20402
rect 25240 20262 25268 20742
rect 25228 20256 25280 20262
rect 25228 20198 25280 20204
rect 25226 20088 25282 20097
rect 25332 20058 25360 20878
rect 25424 20602 25452 20878
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25412 20324 25464 20330
rect 25412 20266 25464 20272
rect 25226 20023 25282 20032
rect 25320 20052 25372 20058
rect 25136 19848 25188 19854
rect 25136 19790 25188 19796
rect 25044 19304 25096 19310
rect 25044 19246 25096 19252
rect 24952 18964 25004 18970
rect 24952 18906 25004 18912
rect 25148 18426 25176 19790
rect 25136 18420 25188 18426
rect 25136 18362 25188 18368
rect 25240 17218 25268 20023
rect 25320 19994 25372 20000
rect 25424 19378 25452 20266
rect 25412 19372 25464 19378
rect 25412 19314 25464 19320
rect 25320 17672 25372 17678
rect 25320 17614 25372 17620
rect 25332 17338 25360 17614
rect 25320 17332 25372 17338
rect 25320 17274 25372 17280
rect 25240 17190 25360 17218
rect 25332 16250 25360 17190
rect 25320 16244 25372 16250
rect 25320 16186 25372 16192
rect 24952 15972 25004 15978
rect 24952 15914 25004 15920
rect 24964 15706 24992 15914
rect 25228 15904 25280 15910
rect 25228 15846 25280 15852
rect 24952 15700 25004 15706
rect 24952 15642 25004 15648
rect 24964 15026 24992 15642
rect 25136 15360 25188 15366
rect 25136 15302 25188 15308
rect 25148 15094 25176 15302
rect 25136 15088 25188 15094
rect 25136 15030 25188 15036
rect 24952 15020 25004 15026
rect 24952 14962 25004 14968
rect 25044 14884 25096 14890
rect 25044 14826 25096 14832
rect 25056 14618 25084 14826
rect 25044 14612 25096 14618
rect 25044 14554 25096 14560
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 25056 14278 25084 14350
rect 25044 14272 25096 14278
rect 25044 14214 25096 14220
rect 25056 13938 25084 14214
rect 25044 13932 25096 13938
rect 25044 13874 25096 13880
rect 25056 13734 25084 13874
rect 25044 13728 25096 13734
rect 25044 13670 25096 13676
rect 25056 13258 25084 13670
rect 25044 13252 25096 13258
rect 25044 13194 25096 13200
rect 25136 12912 25188 12918
rect 25136 12854 25188 12860
rect 24872 12406 24992 12434
rect 24860 12232 24912 12238
rect 24860 12174 24912 12180
rect 24768 12096 24820 12102
rect 24768 12038 24820 12044
rect 24780 11626 24808 12038
rect 24768 11620 24820 11626
rect 24768 11562 24820 11568
rect 24872 11098 24900 12174
rect 24780 11070 24900 11098
rect 24780 10554 24808 11070
rect 24860 11008 24912 11014
rect 24860 10950 24912 10956
rect 24872 10674 24900 10950
rect 24964 10810 24992 12406
rect 24952 10804 25004 10810
rect 24952 10746 25004 10752
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 24780 10526 24900 10554
rect 24872 10266 24900 10526
rect 24860 10260 24912 10266
rect 24860 10202 24912 10208
rect 24768 10056 24820 10062
rect 24768 9998 24820 10004
rect 24780 9654 24808 9998
rect 24872 9722 24900 10202
rect 24860 9716 24912 9722
rect 24860 9658 24912 9664
rect 24768 9648 24820 9654
rect 24768 9590 24820 9596
rect 24216 8968 24268 8974
rect 24216 8910 24268 8916
rect 24032 7472 24084 7478
rect 24032 7414 24084 7420
rect 24044 7002 24072 7414
rect 24228 7206 24256 8910
rect 25044 8832 25096 8838
rect 25044 8774 25096 8780
rect 25056 8566 25084 8774
rect 25044 8560 25096 8566
rect 25044 8502 25096 8508
rect 24216 7200 24268 7206
rect 24216 7142 24268 7148
rect 24400 7200 24452 7206
rect 24400 7142 24452 7148
rect 24032 6996 24084 7002
rect 24032 6938 24084 6944
rect 24044 6458 24072 6938
rect 24032 6452 24084 6458
rect 24032 6394 24084 6400
rect 24412 6390 24440 7142
rect 25148 7002 25176 12854
rect 25240 11898 25268 15846
rect 25332 15434 25360 16186
rect 25516 15502 25544 24006
rect 25700 23866 25728 24375
rect 25688 23860 25740 23866
rect 25688 23802 25740 23808
rect 25596 22636 25648 22642
rect 25596 22578 25648 22584
rect 25608 17882 25636 22578
rect 25780 22568 25832 22574
rect 25780 22510 25832 22516
rect 25792 22098 25820 22510
rect 25780 22092 25832 22098
rect 25780 22034 25832 22040
rect 25780 21888 25832 21894
rect 25780 21830 25832 21836
rect 25688 21140 25740 21146
rect 25688 21082 25740 21088
rect 25700 20097 25728 21082
rect 25792 20466 25820 21830
rect 25884 20602 25912 25298
rect 26068 25226 26096 29786
rect 26252 28966 26280 30194
rect 26240 28960 26292 28966
rect 26240 28902 26292 28908
rect 26252 28694 26280 28902
rect 26240 28688 26292 28694
rect 26240 28630 26292 28636
rect 26148 27872 26200 27878
rect 26148 27814 26200 27820
rect 26160 26926 26188 27814
rect 26148 26920 26200 26926
rect 26148 26862 26200 26868
rect 26344 26382 26372 30518
rect 26436 29850 26464 30654
rect 26516 30592 26568 30598
rect 26516 30534 26568 30540
rect 26528 30258 26556 30534
rect 26516 30252 26568 30258
rect 26516 30194 26568 30200
rect 26514 29880 26570 29889
rect 26424 29844 26476 29850
rect 26514 29815 26516 29824
rect 26424 29786 26476 29792
rect 26568 29815 26570 29824
rect 26516 29786 26568 29792
rect 26608 29504 26660 29510
rect 26608 29446 26660 29452
rect 26516 28212 26568 28218
rect 26516 28154 26568 28160
rect 26424 27464 26476 27470
rect 26424 27406 26476 27412
rect 26332 26376 26384 26382
rect 26332 26318 26384 26324
rect 26148 26240 26200 26246
rect 26148 26182 26200 26188
rect 26160 25906 26188 26182
rect 26148 25900 26200 25906
rect 26148 25842 26200 25848
rect 26240 25764 26292 25770
rect 26240 25706 26292 25712
rect 26252 25498 26280 25706
rect 26240 25492 26292 25498
rect 26240 25434 26292 25440
rect 26148 25288 26200 25294
rect 26148 25230 26200 25236
rect 26056 25220 26108 25226
rect 26056 25162 26108 25168
rect 26160 24426 26188 25230
rect 26252 25140 26280 25434
rect 26344 25294 26372 26318
rect 26436 26314 26464 27406
rect 26424 26308 26476 26314
rect 26424 26250 26476 26256
rect 26332 25288 26384 25294
rect 26332 25230 26384 25236
rect 26252 25112 26372 25140
rect 26160 24398 26280 24426
rect 26148 24336 26200 24342
rect 26148 24278 26200 24284
rect 25964 24200 26016 24206
rect 26160 24188 26188 24278
rect 26016 24160 26188 24188
rect 25964 24142 26016 24148
rect 26252 24120 26280 24398
rect 26344 24206 26372 25112
rect 26424 24948 26476 24954
rect 26424 24890 26476 24896
rect 26332 24200 26384 24206
rect 26332 24142 26384 24148
rect 26068 24092 26280 24120
rect 26068 22166 26096 24092
rect 26344 23848 26372 24142
rect 26436 24138 26464 24890
rect 26528 24410 26556 28154
rect 26620 27436 26648 29446
rect 26712 28082 26740 34070
rect 26804 33930 26832 35974
rect 27252 35692 27304 35698
rect 27252 35634 27304 35640
rect 27160 35080 27212 35086
rect 27160 35022 27212 35028
rect 27172 34610 27200 35022
rect 27160 34604 27212 34610
rect 27160 34546 27212 34552
rect 27264 34202 27292 35634
rect 27540 35630 27568 36042
rect 27528 35624 27580 35630
rect 27528 35566 27580 35572
rect 27804 35624 27856 35630
rect 27804 35566 27856 35572
rect 27436 35080 27488 35086
rect 27436 35022 27488 35028
rect 27448 34678 27476 35022
rect 27712 34944 27764 34950
rect 27712 34886 27764 34892
rect 27436 34672 27488 34678
rect 27436 34614 27488 34620
rect 27252 34196 27304 34202
rect 27252 34138 27304 34144
rect 27344 33992 27396 33998
rect 27344 33934 27396 33940
rect 26792 33924 26844 33930
rect 26792 33866 26844 33872
rect 27356 33658 27384 33934
rect 27344 33652 27396 33658
rect 27344 33594 27396 33600
rect 26884 33448 26936 33454
rect 26884 33390 26936 33396
rect 26896 32026 26924 33390
rect 26976 32768 27028 32774
rect 26976 32710 27028 32716
rect 26884 32020 26936 32026
rect 26884 31962 26936 31968
rect 26896 31822 26924 31962
rect 26884 31816 26936 31822
rect 26884 31758 26936 31764
rect 26792 31748 26844 31754
rect 26792 31690 26844 31696
rect 26700 28076 26752 28082
rect 26700 28018 26752 28024
rect 26804 27674 26832 31690
rect 26884 31272 26936 31278
rect 26884 31214 26936 31220
rect 26896 29646 26924 31214
rect 26884 29640 26936 29646
rect 26884 29582 26936 29588
rect 26896 29238 26924 29582
rect 26884 29232 26936 29238
rect 26884 29174 26936 29180
rect 26792 27668 26844 27674
rect 26792 27610 26844 27616
rect 26700 27464 26752 27470
rect 26608 27430 26660 27436
rect 26700 27406 26752 27412
rect 26884 27464 26936 27470
rect 26884 27406 26936 27412
rect 26608 27372 26660 27378
rect 26712 26994 26740 27406
rect 26700 26988 26752 26994
rect 26700 26930 26752 26936
rect 26896 26790 26924 27406
rect 26884 26784 26936 26790
rect 26884 26726 26936 26732
rect 26700 25832 26752 25838
rect 26700 25774 26752 25780
rect 26516 24404 26568 24410
rect 26516 24346 26568 24352
rect 26516 24268 26568 24274
rect 26516 24210 26568 24216
rect 26528 24177 26556 24210
rect 26712 24206 26740 25774
rect 26884 25288 26936 25294
rect 26884 25230 26936 25236
rect 26792 24744 26844 24750
rect 26792 24686 26844 24692
rect 26700 24200 26752 24206
rect 26514 24168 26570 24177
rect 26424 24132 26476 24138
rect 26700 24142 26752 24148
rect 26514 24103 26570 24112
rect 26424 24074 26476 24080
rect 26160 23820 26372 23848
rect 26160 22574 26188 23820
rect 26332 23724 26384 23730
rect 26332 23666 26384 23672
rect 26240 23520 26292 23526
rect 26240 23462 26292 23468
rect 26252 23118 26280 23462
rect 26240 23112 26292 23118
rect 26240 23054 26292 23060
rect 26148 22568 26200 22574
rect 26148 22510 26200 22516
rect 26056 22160 26108 22166
rect 26056 22102 26108 22108
rect 26068 20942 26096 22102
rect 26056 20936 26108 20942
rect 26056 20878 26108 20884
rect 26148 20868 26200 20874
rect 26148 20810 26200 20816
rect 26054 20632 26110 20641
rect 25872 20596 25924 20602
rect 26054 20567 26110 20576
rect 25872 20538 25924 20544
rect 25780 20460 25832 20466
rect 25780 20402 25832 20408
rect 25686 20088 25742 20097
rect 25686 20023 25742 20032
rect 25792 19446 25820 20402
rect 25780 19440 25832 19446
rect 25780 19382 25832 19388
rect 25884 18834 25912 20538
rect 25964 19984 26016 19990
rect 25964 19926 26016 19932
rect 25872 18828 25924 18834
rect 25872 18770 25924 18776
rect 25780 18216 25832 18222
rect 25780 18158 25832 18164
rect 25596 17876 25648 17882
rect 25596 17818 25648 17824
rect 25688 17536 25740 17542
rect 25688 17478 25740 17484
rect 25504 15496 25556 15502
rect 25504 15438 25556 15444
rect 25320 15428 25372 15434
rect 25320 15370 25372 15376
rect 25412 15020 25464 15026
rect 25412 14962 25464 14968
rect 25424 14618 25452 14962
rect 25412 14612 25464 14618
rect 25412 14554 25464 14560
rect 25596 13456 25648 13462
rect 25596 13398 25648 13404
rect 25410 12880 25466 12889
rect 25608 12850 25636 13398
rect 25410 12815 25412 12824
rect 25464 12815 25466 12824
rect 25596 12844 25648 12850
rect 25412 12786 25464 12792
rect 25596 12786 25648 12792
rect 25228 11892 25280 11898
rect 25228 11834 25280 11840
rect 25240 11218 25268 11834
rect 25228 11212 25280 11218
rect 25228 11154 25280 11160
rect 25240 9654 25268 11154
rect 25700 10470 25728 17478
rect 25792 17134 25820 18158
rect 25780 17128 25832 17134
rect 25780 17070 25832 17076
rect 25792 16046 25820 17070
rect 25780 16040 25832 16046
rect 25780 15982 25832 15988
rect 25792 15026 25820 15982
rect 25872 15632 25924 15638
rect 25872 15574 25924 15580
rect 25780 15020 25832 15026
rect 25780 14962 25832 14968
rect 25792 14414 25820 14962
rect 25780 14408 25832 14414
rect 25780 14350 25832 14356
rect 25884 13938 25912 15574
rect 25872 13932 25924 13938
rect 25872 13874 25924 13880
rect 25870 13696 25926 13705
rect 25870 13631 25926 13640
rect 25884 13326 25912 13631
rect 25872 13320 25924 13326
rect 25872 13262 25924 13268
rect 25976 12306 26004 19926
rect 26068 19378 26096 20567
rect 26056 19372 26108 19378
rect 26056 19314 26108 19320
rect 26056 17196 26108 17202
rect 26056 17138 26108 17144
rect 26068 16522 26096 17138
rect 26056 16516 26108 16522
rect 26056 16458 26108 16464
rect 26056 16040 26108 16046
rect 26056 15982 26108 15988
rect 26068 15638 26096 15982
rect 26056 15632 26108 15638
rect 26056 15574 26108 15580
rect 26160 12434 26188 20810
rect 26252 19417 26280 23054
rect 26344 21554 26372 23666
rect 26436 22710 26464 24074
rect 26608 23860 26660 23866
rect 26608 23802 26660 23808
rect 26424 22704 26476 22710
rect 26424 22646 26476 22652
rect 26620 21554 26648 23802
rect 26804 23798 26832 24686
rect 26792 23792 26844 23798
rect 26792 23734 26844 23740
rect 26790 23216 26846 23225
rect 26790 23151 26846 23160
rect 26804 23118 26832 23151
rect 26792 23112 26844 23118
rect 26896 23100 26924 25230
rect 26988 23730 27016 32710
rect 27160 32224 27212 32230
rect 27160 32166 27212 32172
rect 27068 29028 27120 29034
rect 27068 28970 27120 28976
rect 26976 23724 27028 23730
rect 26976 23666 27028 23672
rect 27080 23662 27108 28970
rect 27172 28150 27200 32166
rect 27356 31906 27384 33594
rect 27448 33538 27476 34614
rect 27724 33998 27752 34886
rect 27712 33992 27764 33998
rect 27712 33934 27764 33940
rect 27448 33522 27660 33538
rect 27448 33516 27672 33522
rect 27448 33510 27620 33516
rect 27620 33458 27672 33464
rect 27436 33380 27488 33386
rect 27436 33322 27488 33328
rect 27264 31878 27384 31906
rect 27264 31346 27292 31878
rect 27448 31668 27476 33322
rect 27528 32496 27580 32502
rect 27528 32438 27580 32444
rect 27540 31890 27568 32438
rect 27528 31884 27580 31890
rect 27528 31826 27580 31832
rect 27712 31816 27764 31822
rect 27356 31640 27476 31668
rect 27632 31776 27712 31804
rect 27252 31340 27304 31346
rect 27252 31282 27304 31288
rect 27264 30870 27292 31282
rect 27252 30864 27304 30870
rect 27252 30806 27304 30812
rect 27252 28756 27304 28762
rect 27252 28698 27304 28704
rect 27264 28422 27292 28698
rect 27252 28416 27304 28422
rect 27252 28358 27304 28364
rect 27160 28144 27212 28150
rect 27160 28086 27212 28092
rect 27172 27674 27200 28086
rect 27160 27668 27212 27674
rect 27160 27610 27212 27616
rect 27264 27554 27292 28358
rect 27356 27946 27384 31640
rect 27436 31476 27488 31482
rect 27436 31418 27488 31424
rect 27448 31346 27476 31418
rect 27436 31340 27488 31346
rect 27436 31282 27488 31288
rect 27448 30802 27476 31282
rect 27632 31278 27660 31776
rect 27712 31758 27764 31764
rect 27620 31272 27672 31278
rect 27620 31214 27672 31220
rect 27436 30796 27488 30802
rect 27436 30738 27488 30744
rect 27436 30592 27488 30598
rect 27436 30534 27488 30540
rect 27344 27940 27396 27946
rect 27344 27882 27396 27888
rect 27448 27878 27476 30534
rect 27528 29640 27580 29646
rect 27528 29582 27580 29588
rect 27540 29034 27568 29582
rect 27632 29170 27660 31214
rect 27712 30728 27764 30734
rect 27710 30696 27712 30705
rect 27764 30696 27766 30705
rect 27710 30631 27766 30640
rect 27710 30288 27766 30297
rect 27710 30223 27766 30232
rect 27724 30190 27752 30223
rect 27712 30184 27764 30190
rect 27712 30126 27764 30132
rect 27712 29708 27764 29714
rect 27712 29650 27764 29656
rect 27724 29238 27752 29650
rect 27712 29232 27764 29238
rect 27712 29174 27764 29180
rect 27620 29164 27672 29170
rect 27620 29106 27672 29112
rect 27632 29073 27660 29106
rect 27618 29064 27674 29073
rect 27528 29028 27580 29034
rect 27618 28999 27674 29008
rect 27816 28994 27844 35566
rect 27896 33924 27948 33930
rect 27896 33866 27948 33872
rect 27908 31482 27936 33866
rect 27988 33448 28040 33454
rect 27988 33390 28040 33396
rect 28000 32910 28028 33390
rect 27988 32904 28040 32910
rect 27988 32846 28040 32852
rect 27896 31476 27948 31482
rect 27896 31418 27948 31424
rect 27908 31278 27936 31418
rect 27896 31272 27948 31278
rect 27896 31214 27948 31220
rect 27896 30796 27948 30802
rect 27896 30738 27948 30744
rect 27908 29578 27936 30738
rect 27988 30660 28040 30666
rect 27988 30602 28040 30608
rect 27896 29572 27948 29578
rect 27896 29514 27948 29520
rect 27528 28970 27580 28976
rect 27724 28966 27844 28994
rect 27620 28416 27672 28422
rect 27620 28358 27672 28364
rect 27528 27940 27580 27946
rect 27528 27882 27580 27888
rect 27436 27872 27488 27878
rect 27436 27814 27488 27820
rect 27540 27690 27568 27882
rect 27632 27713 27660 28358
rect 27172 27526 27292 27554
rect 27448 27662 27568 27690
rect 27618 27704 27674 27713
rect 27172 25838 27200 27526
rect 27252 27328 27304 27334
rect 27252 27270 27304 27276
rect 27160 25832 27212 25838
rect 27160 25774 27212 25780
rect 27160 24200 27212 24206
rect 27160 24142 27212 24148
rect 27172 23798 27200 24142
rect 27160 23792 27212 23798
rect 27160 23734 27212 23740
rect 27068 23656 27120 23662
rect 27068 23598 27120 23604
rect 26896 23072 27016 23100
rect 26792 23054 26844 23060
rect 26804 22094 26832 23054
rect 26988 22953 27016 23072
rect 26974 22944 27030 22953
rect 26974 22879 27030 22888
rect 26804 22066 26924 22094
rect 26792 22024 26844 22030
rect 26790 21992 26792 22001
rect 26844 21992 26846 22001
rect 26700 21956 26752 21962
rect 26790 21927 26846 21936
rect 26700 21898 26752 21904
rect 26712 21554 26740 21898
rect 26896 21690 26924 22066
rect 26884 21684 26936 21690
rect 26884 21626 26936 21632
rect 26332 21548 26384 21554
rect 26332 21490 26384 21496
rect 26608 21548 26660 21554
rect 26608 21490 26660 21496
rect 26700 21548 26752 21554
rect 26700 21490 26752 21496
rect 26344 21146 26372 21490
rect 26332 21140 26384 21146
rect 26332 21082 26384 21088
rect 26344 20262 26372 21082
rect 26620 20466 26648 21490
rect 26700 20528 26752 20534
rect 26700 20470 26752 20476
rect 26608 20460 26660 20466
rect 26608 20402 26660 20408
rect 26424 20392 26476 20398
rect 26424 20334 26476 20340
rect 26332 20256 26384 20262
rect 26332 20198 26384 20204
rect 26332 19984 26384 19990
rect 26332 19926 26384 19932
rect 26238 19408 26294 19417
rect 26344 19378 26372 19926
rect 26436 19378 26464 20334
rect 26238 19343 26294 19352
rect 26332 19372 26384 19378
rect 26332 19314 26384 19320
rect 26424 19372 26476 19378
rect 26424 19314 26476 19320
rect 26344 17762 26372 19314
rect 26252 17734 26372 17762
rect 26252 16590 26280 17734
rect 26332 17672 26384 17678
rect 26332 17614 26384 17620
rect 26344 17202 26372 17614
rect 26436 17202 26464 19314
rect 26608 19168 26660 19174
rect 26608 19110 26660 19116
rect 26620 17678 26648 19110
rect 26608 17672 26660 17678
rect 26608 17614 26660 17620
rect 26712 17610 26740 20470
rect 26884 20256 26936 20262
rect 26884 20198 26936 20204
rect 26896 19854 26924 20198
rect 26884 19848 26936 19854
rect 26884 19790 26936 19796
rect 26896 19514 26924 19790
rect 26884 19508 26936 19514
rect 26884 19450 26936 19456
rect 26896 19378 26924 19450
rect 26884 19372 26936 19378
rect 26884 19314 26936 19320
rect 26792 18624 26844 18630
rect 26792 18566 26844 18572
rect 26700 17604 26752 17610
rect 26700 17546 26752 17552
rect 26332 17196 26384 17202
rect 26332 17138 26384 17144
rect 26424 17196 26476 17202
rect 26424 17138 26476 17144
rect 26344 16726 26372 17138
rect 26332 16720 26384 16726
rect 26332 16662 26384 16668
rect 26436 16658 26464 17138
rect 26424 16652 26476 16658
rect 26424 16594 26476 16600
rect 26712 16590 26740 17546
rect 26240 16584 26292 16590
rect 26240 16526 26292 16532
rect 26516 16584 26568 16590
rect 26516 16526 26568 16532
rect 26700 16584 26752 16590
rect 26700 16526 26752 16532
rect 26528 16425 26556 16526
rect 26804 16522 26832 18566
rect 26988 18290 27016 22879
rect 27264 22094 27292 27270
rect 27448 26874 27476 27662
rect 27618 27639 27674 27648
rect 27620 27464 27672 27470
rect 27620 27406 27672 27412
rect 27356 26846 27476 26874
rect 27526 26888 27582 26897
rect 27356 24052 27384 26846
rect 27526 26823 27582 26832
rect 27540 25906 27568 26823
rect 27632 26450 27660 27406
rect 27724 26926 27752 28966
rect 27804 27872 27856 27878
rect 27804 27814 27856 27820
rect 27816 27130 27844 27814
rect 27804 27124 27856 27130
rect 27804 27066 27856 27072
rect 27712 26920 27764 26926
rect 27712 26862 27764 26868
rect 27620 26444 27672 26450
rect 27620 26386 27672 26392
rect 27618 26208 27674 26217
rect 27618 26143 27674 26152
rect 27528 25900 27580 25906
rect 27528 25842 27580 25848
rect 27434 24848 27490 24857
rect 27434 24783 27490 24792
rect 27448 24206 27476 24783
rect 27436 24200 27488 24206
rect 27436 24142 27488 24148
rect 27528 24132 27580 24138
rect 27528 24074 27580 24080
rect 27356 24024 27476 24052
rect 27344 23724 27396 23730
rect 27344 23666 27396 23672
rect 27356 23633 27384 23666
rect 27342 23624 27398 23633
rect 27342 23559 27398 23568
rect 27344 23180 27396 23186
rect 27344 23122 27396 23128
rect 27356 22710 27384 23122
rect 27344 22704 27396 22710
rect 27344 22646 27396 22652
rect 27172 22066 27292 22094
rect 27068 21956 27120 21962
rect 27068 21898 27120 21904
rect 27080 21622 27108 21898
rect 27068 21616 27120 21622
rect 27068 21558 27120 21564
rect 27068 20800 27120 20806
rect 27066 20768 27068 20777
rect 27120 20768 27122 20777
rect 27066 20703 27122 20712
rect 27068 19780 27120 19786
rect 27068 19722 27120 19728
rect 27080 19417 27108 19722
rect 27066 19408 27122 19417
rect 27066 19343 27122 19352
rect 27080 19310 27108 19343
rect 27068 19304 27120 19310
rect 27068 19246 27120 19252
rect 26976 18284 27028 18290
rect 26976 18226 27028 18232
rect 27172 18222 27200 22066
rect 27252 21888 27304 21894
rect 27252 21830 27304 21836
rect 27264 21690 27292 21830
rect 27252 21684 27304 21690
rect 27252 21626 27304 21632
rect 27252 21480 27304 21486
rect 27252 21422 27304 21428
rect 27264 20942 27292 21422
rect 27252 20936 27304 20942
rect 27252 20878 27304 20884
rect 27264 20346 27292 20878
rect 27356 20534 27384 22646
rect 27448 21622 27476 24024
rect 27540 22114 27568 24074
rect 27632 22778 27660 26143
rect 27712 25220 27764 25226
rect 27712 25162 27764 25168
rect 27724 23866 27752 25162
rect 27908 24936 27936 29514
rect 28000 29102 28028 30602
rect 27988 29096 28040 29102
rect 27988 29038 28040 29044
rect 28000 28762 28028 29038
rect 27988 28756 28040 28762
rect 27988 28698 28040 28704
rect 28000 28150 28028 28698
rect 27988 28144 28040 28150
rect 27988 28086 28040 28092
rect 28092 26518 28120 37266
rect 28276 37262 28304 39200
rect 30472 37324 30524 37330
rect 30472 37266 30524 37272
rect 28264 37256 28316 37262
rect 28264 37198 28316 37204
rect 28448 37120 28500 37126
rect 28448 37062 28500 37068
rect 28356 36916 28408 36922
rect 28356 36858 28408 36864
rect 28172 36780 28224 36786
rect 28172 36722 28224 36728
rect 28184 36378 28212 36722
rect 28264 36576 28316 36582
rect 28368 36530 28396 36858
rect 28316 36524 28396 36530
rect 28264 36518 28396 36524
rect 28276 36502 28396 36518
rect 28172 36372 28224 36378
rect 28172 36314 28224 36320
rect 28368 36174 28396 36502
rect 28356 36168 28408 36174
rect 28356 36110 28408 36116
rect 28172 32904 28224 32910
rect 28172 32846 28224 32852
rect 28184 32298 28212 32846
rect 28460 32586 28488 37062
rect 30484 36786 30512 37266
rect 31588 37210 31616 39200
rect 34900 37754 34928 39200
rect 36818 38312 36874 38321
rect 36818 38247 36874 38256
rect 34808 37726 34928 37754
rect 32680 37324 32732 37330
rect 32680 37266 32732 37272
rect 31760 37256 31812 37262
rect 31588 37204 31760 37210
rect 31588 37198 31812 37204
rect 31588 37182 31800 37198
rect 31024 37120 31076 37126
rect 31024 37062 31076 37068
rect 28632 36780 28684 36786
rect 28632 36722 28684 36728
rect 30472 36780 30524 36786
rect 30472 36722 30524 36728
rect 28644 35698 28672 36722
rect 29276 36576 29328 36582
rect 29276 36518 29328 36524
rect 30104 36576 30156 36582
rect 30104 36518 30156 36524
rect 29288 36106 29316 36518
rect 30116 36378 30144 36518
rect 30104 36372 30156 36378
rect 30104 36314 30156 36320
rect 30484 36242 30512 36722
rect 30472 36236 30524 36242
rect 30472 36178 30524 36184
rect 30012 36168 30064 36174
rect 30012 36110 30064 36116
rect 29276 36100 29328 36106
rect 29276 36042 29328 36048
rect 29092 36032 29144 36038
rect 29092 35974 29144 35980
rect 28632 35692 28684 35698
rect 28632 35634 28684 35640
rect 28908 35692 28960 35698
rect 28908 35634 28960 35640
rect 28540 35488 28592 35494
rect 28540 35430 28592 35436
rect 28552 34610 28580 35430
rect 28920 35290 28948 35634
rect 28908 35284 28960 35290
rect 28908 35226 28960 35232
rect 29104 35154 29132 35974
rect 29092 35148 29144 35154
rect 29092 35090 29144 35096
rect 28908 35080 28960 35086
rect 28908 35022 28960 35028
rect 28920 34649 28948 35022
rect 29184 35012 29236 35018
rect 29184 34954 29236 34960
rect 28906 34640 28962 34649
rect 28540 34604 28592 34610
rect 28906 34575 28962 34584
rect 29092 34604 29144 34610
rect 28540 34546 28592 34552
rect 29092 34546 29144 34552
rect 28368 32558 28488 32586
rect 28264 32360 28316 32366
rect 28264 32302 28316 32308
rect 28172 32292 28224 32298
rect 28172 32234 28224 32240
rect 28184 30598 28212 32234
rect 28276 31890 28304 32302
rect 28368 31906 28396 32558
rect 28448 32428 28500 32434
rect 28448 32370 28500 32376
rect 28460 32026 28488 32370
rect 28448 32020 28500 32026
rect 28448 31962 28500 31968
rect 28264 31884 28316 31890
rect 28368 31878 28488 31906
rect 28264 31826 28316 31832
rect 28276 31482 28304 31826
rect 28264 31476 28316 31482
rect 28264 31418 28316 31424
rect 28172 30592 28224 30598
rect 28172 30534 28224 30540
rect 28172 30320 28224 30326
rect 28172 30262 28224 30268
rect 28184 29170 28212 30262
rect 28356 30252 28408 30258
rect 28356 30194 28408 30200
rect 28368 29782 28396 30194
rect 28356 29776 28408 29782
rect 28356 29718 28408 29724
rect 28172 29164 28224 29170
rect 28172 29106 28224 29112
rect 28356 29028 28408 29034
rect 28356 28970 28408 28976
rect 28368 28558 28396 28970
rect 28460 28694 28488 31878
rect 28448 28688 28500 28694
rect 28448 28630 28500 28636
rect 28356 28552 28408 28558
rect 28356 28494 28408 28500
rect 28264 28484 28316 28490
rect 28264 28426 28316 28432
rect 28080 26512 28132 26518
rect 28080 26454 28132 26460
rect 28080 26376 28132 26382
rect 28080 26318 28132 26324
rect 27986 26072 28042 26081
rect 27986 26007 28042 26016
rect 28000 25838 28028 26007
rect 27988 25832 28040 25838
rect 27988 25774 28040 25780
rect 28092 25498 28120 26318
rect 28276 26217 28304 28426
rect 28262 26208 28318 26217
rect 28262 26143 28318 26152
rect 28368 25838 28396 28494
rect 28448 28144 28500 28150
rect 28448 28086 28500 28092
rect 28460 27470 28488 28086
rect 28448 27464 28500 27470
rect 28448 27406 28500 27412
rect 28448 27328 28500 27334
rect 28448 27270 28500 27276
rect 28460 27062 28488 27270
rect 28448 27056 28500 27062
rect 28448 26998 28500 27004
rect 28552 26450 28580 34546
rect 29000 34400 29052 34406
rect 29000 34342 29052 34348
rect 29012 34066 29040 34342
rect 29000 34060 29052 34066
rect 29000 34002 29052 34008
rect 28724 33856 28776 33862
rect 28724 33798 28776 33804
rect 28736 33658 28764 33798
rect 28724 33652 28776 33658
rect 28724 33594 28776 33600
rect 29104 33386 29132 34546
rect 29196 34542 29224 34954
rect 29184 34536 29236 34542
rect 29184 34478 29236 34484
rect 29196 33998 29224 34478
rect 29288 34066 29316 36042
rect 30024 35494 30052 36110
rect 30012 35488 30064 35494
rect 30012 35430 30064 35436
rect 31036 35086 31064 37062
rect 32404 36780 32456 36786
rect 32404 36722 32456 36728
rect 32416 36378 32444 36722
rect 32692 36378 32720 37266
rect 33784 37256 33836 37262
rect 33784 37198 33836 37204
rect 32772 36848 32824 36854
rect 32772 36790 32824 36796
rect 32404 36372 32456 36378
rect 32404 36314 32456 36320
rect 32680 36372 32732 36378
rect 32680 36314 32732 36320
rect 32312 36304 32364 36310
rect 32312 36246 32364 36252
rect 31208 36236 31260 36242
rect 31208 36178 31260 36184
rect 31220 35290 31248 36178
rect 32036 35760 32088 35766
rect 32036 35702 32088 35708
rect 31208 35284 31260 35290
rect 31208 35226 31260 35232
rect 31668 35216 31720 35222
rect 31668 35158 31720 35164
rect 31680 35086 31708 35158
rect 30656 35080 30708 35086
rect 30748 35080 30800 35086
rect 30656 35022 30708 35028
rect 30746 35048 30748 35057
rect 31024 35080 31076 35086
rect 30800 35048 30802 35057
rect 29276 34060 29328 34066
rect 29276 34002 29328 34008
rect 29184 33992 29236 33998
rect 29184 33934 29236 33940
rect 29092 33380 29144 33386
rect 29092 33322 29144 33328
rect 28724 32972 28776 32978
rect 28724 32914 28776 32920
rect 28736 32298 28764 32914
rect 28908 32904 28960 32910
rect 28908 32846 28960 32852
rect 28816 32428 28868 32434
rect 28816 32370 28868 32376
rect 28724 32292 28776 32298
rect 28724 32234 28776 32240
rect 28632 31680 28684 31686
rect 28632 31622 28684 31628
rect 28644 31346 28672 31622
rect 28632 31340 28684 31346
rect 28632 31282 28684 31288
rect 28632 30592 28684 30598
rect 28632 30534 28684 30540
rect 28644 30054 28672 30534
rect 28736 30190 28764 32234
rect 28828 31958 28856 32370
rect 28920 32042 28948 32846
rect 28920 32014 29040 32042
rect 29012 31958 29040 32014
rect 28816 31952 28868 31958
rect 28816 31894 28868 31900
rect 29000 31952 29052 31958
rect 29000 31894 29052 31900
rect 29092 31816 29144 31822
rect 28906 31784 28962 31793
rect 28906 31719 28908 31728
rect 28960 31719 28962 31728
rect 29012 31776 29092 31804
rect 28908 31690 28960 31696
rect 29012 31414 29040 31776
rect 29092 31758 29144 31764
rect 29000 31408 29052 31414
rect 29000 31350 29052 31356
rect 29184 31340 29236 31346
rect 29184 31282 29236 31288
rect 28908 31272 28960 31278
rect 28908 31214 28960 31220
rect 28920 30954 28948 31214
rect 28920 30926 29040 30954
rect 28908 30864 28960 30870
rect 28908 30806 28960 30812
rect 28920 30258 28948 30806
rect 29012 30734 29040 30926
rect 29000 30728 29052 30734
rect 29000 30670 29052 30676
rect 28908 30252 28960 30258
rect 28908 30194 28960 30200
rect 28724 30184 28776 30190
rect 28724 30126 28776 30132
rect 28632 30048 28684 30054
rect 28632 29990 28684 29996
rect 28644 27062 28672 29990
rect 28724 29028 28776 29034
rect 28724 28970 28776 28976
rect 28736 27849 28764 28970
rect 28908 28688 28960 28694
rect 28908 28630 28960 28636
rect 28816 28552 28868 28558
rect 28816 28494 28868 28500
rect 28828 28082 28856 28494
rect 28920 28218 28948 28630
rect 28908 28212 28960 28218
rect 28908 28154 28960 28160
rect 28816 28076 28868 28082
rect 28816 28018 28868 28024
rect 28920 27878 28948 28154
rect 28816 27872 28868 27878
rect 28722 27840 28778 27849
rect 28816 27814 28868 27820
rect 28908 27872 28960 27878
rect 28908 27814 28960 27820
rect 28722 27775 28778 27784
rect 28828 27713 28856 27814
rect 28814 27704 28870 27713
rect 28814 27639 28870 27648
rect 28908 27464 28960 27470
rect 28908 27406 28960 27412
rect 28632 27056 28684 27062
rect 28632 26998 28684 27004
rect 28920 26586 28948 27406
rect 29092 27396 29144 27402
rect 29092 27338 29144 27344
rect 29104 27130 29132 27338
rect 29092 27124 29144 27130
rect 29092 27066 29144 27072
rect 29000 26988 29052 26994
rect 29000 26930 29052 26936
rect 28908 26580 28960 26586
rect 28908 26522 28960 26528
rect 28632 26512 28684 26518
rect 28632 26454 28684 26460
rect 28540 26444 28592 26450
rect 28540 26386 28592 26392
rect 28448 26240 28500 26246
rect 28448 26182 28500 26188
rect 28460 25906 28488 26182
rect 28448 25900 28500 25906
rect 28448 25842 28500 25848
rect 28356 25832 28408 25838
rect 28356 25774 28408 25780
rect 28172 25696 28224 25702
rect 28172 25638 28224 25644
rect 28080 25492 28132 25498
rect 28080 25434 28132 25440
rect 27816 24908 27936 24936
rect 27816 24206 27844 24908
rect 27988 24880 28040 24886
rect 27988 24822 28040 24828
rect 27896 24812 27948 24818
rect 27896 24754 27948 24760
rect 27908 24410 27936 24754
rect 27896 24404 27948 24410
rect 27896 24346 27948 24352
rect 27804 24200 27856 24206
rect 27804 24142 27856 24148
rect 27896 24200 27948 24206
rect 27896 24142 27948 24148
rect 27712 23860 27764 23866
rect 27712 23802 27764 23808
rect 27712 23112 27764 23118
rect 27710 23080 27712 23089
rect 27764 23080 27766 23089
rect 27710 23015 27766 23024
rect 27620 22772 27672 22778
rect 27620 22714 27672 22720
rect 27620 22636 27672 22642
rect 27620 22578 27672 22584
rect 27712 22636 27764 22642
rect 27712 22578 27764 22584
rect 27632 22234 27660 22578
rect 27620 22228 27672 22234
rect 27620 22170 27672 22176
rect 27724 22166 27752 22578
rect 27712 22160 27764 22166
rect 27540 22086 27660 22114
rect 27712 22102 27764 22108
rect 27528 21888 27580 21894
rect 27528 21830 27580 21836
rect 27436 21616 27488 21622
rect 27436 21558 27488 21564
rect 27436 21344 27488 21350
rect 27436 21286 27488 21292
rect 27344 20528 27396 20534
rect 27344 20470 27396 20476
rect 27264 20318 27384 20346
rect 27160 18216 27212 18222
rect 27160 18158 27212 18164
rect 27158 17776 27214 17785
rect 27356 17746 27384 20318
rect 27448 18714 27476 21286
rect 27540 20942 27568 21830
rect 27632 21622 27660 22086
rect 27712 22024 27764 22030
rect 27816 22012 27844 24142
rect 27908 23798 27936 24142
rect 27896 23792 27948 23798
rect 27896 23734 27948 23740
rect 27896 23588 27948 23594
rect 27896 23530 27948 23536
rect 27908 23186 27936 23530
rect 27896 23180 27948 23186
rect 27896 23122 27948 23128
rect 27908 22642 27936 23122
rect 28000 23118 28028 24822
rect 28080 24132 28132 24138
rect 28080 24074 28132 24080
rect 27988 23112 28040 23118
rect 27988 23054 28040 23060
rect 27896 22636 27948 22642
rect 27896 22578 27948 22584
rect 28000 22030 28028 23054
rect 27764 21984 27844 22012
rect 27712 21966 27764 21972
rect 27620 21616 27672 21622
rect 27620 21558 27672 21564
rect 27816 21350 27844 21984
rect 27896 22024 27948 22030
rect 27896 21966 27948 21972
rect 27988 22024 28040 22030
rect 27988 21966 28040 21972
rect 27804 21344 27856 21350
rect 27804 21286 27856 21292
rect 27528 20936 27580 20942
rect 27528 20878 27580 20884
rect 27620 20936 27672 20942
rect 27620 20878 27672 20884
rect 27632 20602 27660 20878
rect 27620 20596 27672 20602
rect 27620 20538 27672 20544
rect 27528 20528 27580 20534
rect 27528 20470 27580 20476
rect 27540 19514 27568 20470
rect 27816 20398 27844 21286
rect 27908 20942 27936 21966
rect 27988 21888 28040 21894
rect 27988 21830 28040 21836
rect 27896 20936 27948 20942
rect 27896 20878 27948 20884
rect 28000 20788 28028 21830
rect 27908 20760 28028 20788
rect 27804 20392 27856 20398
rect 27804 20334 27856 20340
rect 27528 19508 27580 19514
rect 27528 19450 27580 19456
rect 27908 18834 27936 20760
rect 28092 20602 28120 24074
rect 28080 20596 28132 20602
rect 28080 20538 28132 20544
rect 27988 20392 28040 20398
rect 27988 20334 28040 20340
rect 28000 19854 28028 20334
rect 28092 19922 28120 20538
rect 28080 19916 28132 19922
rect 28080 19858 28132 19864
rect 27988 19848 28040 19854
rect 27988 19790 28040 19796
rect 27896 18828 27948 18834
rect 27896 18770 27948 18776
rect 27448 18686 27568 18714
rect 27158 17711 27214 17720
rect 27344 17740 27396 17746
rect 27172 17678 27200 17711
rect 27344 17682 27396 17688
rect 27160 17672 27212 17678
rect 27212 17632 27292 17660
rect 27160 17614 27212 17620
rect 26792 16516 26844 16522
rect 26792 16458 26844 16464
rect 26514 16416 26570 16425
rect 26514 16351 26570 16360
rect 26528 16114 26556 16351
rect 26516 16108 26568 16114
rect 26516 16050 26568 16056
rect 26528 15570 26556 16050
rect 26804 15706 26832 16458
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 26976 15972 27028 15978
rect 26976 15914 27028 15920
rect 26792 15700 26844 15706
rect 26792 15642 26844 15648
rect 26516 15564 26568 15570
rect 26516 15506 26568 15512
rect 26988 15502 27016 15914
rect 27172 15502 27200 16050
rect 26976 15496 27028 15502
rect 26976 15438 27028 15444
rect 27160 15496 27212 15502
rect 27160 15438 27212 15444
rect 26238 15328 26294 15337
rect 26238 15263 26294 15272
rect 26252 15094 26280 15263
rect 26240 15088 26292 15094
rect 26240 15030 26292 15036
rect 26988 13938 27016 15438
rect 27158 15192 27214 15201
rect 27158 15127 27214 15136
rect 27172 14006 27200 15127
rect 27264 14346 27292 17632
rect 27356 17270 27384 17682
rect 27434 17640 27490 17649
rect 27434 17575 27436 17584
rect 27488 17575 27490 17584
rect 27436 17546 27488 17552
rect 27344 17264 27396 17270
rect 27344 17206 27396 17212
rect 27436 17196 27488 17202
rect 27436 17138 27488 17144
rect 27344 17128 27396 17134
rect 27344 17070 27396 17076
rect 27356 16658 27384 17070
rect 27448 16833 27476 17138
rect 27434 16824 27490 16833
rect 27434 16759 27490 16768
rect 27344 16652 27396 16658
rect 27344 16594 27396 16600
rect 27344 15904 27396 15910
rect 27344 15846 27396 15852
rect 27252 14340 27304 14346
rect 27252 14282 27304 14288
rect 27264 14006 27292 14282
rect 27160 14000 27212 14006
rect 27160 13942 27212 13948
rect 27252 14000 27304 14006
rect 27252 13942 27304 13948
rect 26332 13932 26384 13938
rect 26332 13874 26384 13880
rect 26976 13932 27028 13938
rect 26976 13874 27028 13880
rect 26344 12442 26372 13874
rect 26976 13728 27028 13734
rect 26976 13670 27028 13676
rect 26988 13394 27016 13670
rect 26976 13388 27028 13394
rect 26976 13330 27028 13336
rect 26332 12436 26384 12442
rect 26160 12406 26280 12434
rect 25964 12300 26016 12306
rect 26016 12260 26188 12288
rect 25964 12242 26016 12248
rect 25780 12164 25832 12170
rect 25780 12106 25832 12112
rect 25792 11898 25820 12106
rect 25872 12096 25924 12102
rect 25872 12038 25924 12044
rect 25780 11892 25832 11898
rect 25780 11834 25832 11840
rect 25780 11688 25832 11694
rect 25780 11630 25832 11636
rect 25688 10464 25740 10470
rect 25688 10406 25740 10412
rect 25228 9648 25280 9654
rect 25228 9590 25280 9596
rect 25240 9042 25268 9590
rect 25320 9512 25372 9518
rect 25320 9454 25372 9460
rect 25228 9036 25280 9042
rect 25228 8978 25280 8984
rect 25332 8838 25360 9454
rect 25688 9036 25740 9042
rect 25688 8978 25740 8984
rect 25320 8832 25372 8838
rect 25320 8774 25372 8780
rect 25136 6996 25188 7002
rect 25136 6938 25188 6944
rect 23848 6384 23900 6390
rect 23848 6326 23900 6332
rect 24400 6384 24452 6390
rect 24400 6326 24452 6332
rect 23860 5778 23888 6326
rect 24676 6316 24728 6322
rect 24676 6258 24728 6264
rect 23848 5772 23900 5778
rect 23848 5714 23900 5720
rect 23664 4752 23716 4758
rect 23664 4694 23716 4700
rect 23572 4684 23624 4690
rect 23572 4626 23624 4632
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 23584 4078 23612 4626
rect 23860 4486 23888 5714
rect 24584 5568 24636 5574
rect 24584 5510 24636 5516
rect 24596 5302 24624 5510
rect 24688 5370 24716 6258
rect 25332 5778 25360 8774
rect 25700 8430 25728 8978
rect 25688 8424 25740 8430
rect 25688 8366 25740 8372
rect 25792 6866 25820 11630
rect 25884 10266 25912 12038
rect 25964 11824 26016 11830
rect 25964 11766 26016 11772
rect 26056 11824 26108 11830
rect 26056 11766 26108 11772
rect 25976 11082 26004 11766
rect 25964 11076 26016 11082
rect 25964 11018 26016 11024
rect 25976 10810 26004 11018
rect 25964 10804 26016 10810
rect 25964 10746 26016 10752
rect 25872 10260 25924 10266
rect 25872 10202 25924 10208
rect 26068 9042 26096 11766
rect 26160 11694 26188 12260
rect 26252 11694 26280 12406
rect 26332 12378 26384 12384
rect 26148 11688 26200 11694
rect 26148 11630 26200 11636
rect 26240 11688 26292 11694
rect 26240 11630 26292 11636
rect 26148 11552 26200 11558
rect 26148 11494 26200 11500
rect 26056 9036 26108 9042
rect 26056 8978 26108 8984
rect 25872 8968 25924 8974
rect 25872 8910 25924 8916
rect 25884 8634 25912 8910
rect 25872 8628 25924 8634
rect 25872 8570 25924 8576
rect 26068 7546 26096 8978
rect 26160 8906 26188 11494
rect 26252 10674 26280 11630
rect 26700 11144 26752 11150
rect 26700 11086 26752 11092
rect 27252 11144 27304 11150
rect 27252 11086 27304 11092
rect 26712 10742 26740 11086
rect 27160 11076 27212 11082
rect 27160 11018 27212 11024
rect 27172 10810 27200 11018
rect 27160 10804 27212 10810
rect 27160 10746 27212 10752
rect 26700 10736 26752 10742
rect 26700 10678 26752 10684
rect 26240 10668 26292 10674
rect 26240 10610 26292 10616
rect 26712 10130 26740 10678
rect 27264 10606 27292 11086
rect 27252 10600 27304 10606
rect 27252 10542 27304 10548
rect 26332 10124 26384 10130
rect 26332 10066 26384 10072
rect 26700 10124 26752 10130
rect 26700 10066 26752 10072
rect 26240 9988 26292 9994
rect 26240 9930 26292 9936
rect 26252 9722 26280 9930
rect 26240 9716 26292 9722
rect 26240 9658 26292 9664
rect 26148 8900 26200 8906
rect 26148 8842 26200 8848
rect 26056 7540 26108 7546
rect 26056 7482 26108 7488
rect 26068 6934 26096 7482
rect 26056 6928 26108 6934
rect 26056 6870 26108 6876
rect 25780 6860 25832 6866
rect 25780 6802 25832 6808
rect 25412 6724 25464 6730
rect 25412 6666 25464 6672
rect 25424 6458 25452 6666
rect 25964 6656 26016 6662
rect 25964 6598 26016 6604
rect 25412 6452 25464 6458
rect 25412 6394 25464 6400
rect 25976 5914 26004 6598
rect 26068 6304 26096 6870
rect 26160 6866 26188 8842
rect 26148 6860 26200 6866
rect 26148 6802 26200 6808
rect 26160 6458 26188 6802
rect 26252 6798 26280 9658
rect 26344 9178 26372 10066
rect 26424 9648 26476 9654
rect 26424 9590 26476 9596
rect 26332 9172 26384 9178
rect 26332 9114 26384 9120
rect 26240 6792 26292 6798
rect 26240 6734 26292 6740
rect 26148 6452 26200 6458
rect 26148 6394 26200 6400
rect 26436 6390 26464 9590
rect 26712 9586 26740 10066
rect 26700 9580 26752 9586
rect 26620 9540 26700 9568
rect 26516 8424 26568 8430
rect 26516 8366 26568 8372
rect 26424 6384 26476 6390
rect 26424 6326 26476 6332
rect 26148 6316 26200 6322
rect 26068 6276 26148 6304
rect 26148 6258 26200 6264
rect 26240 6180 26292 6186
rect 26240 6122 26292 6128
rect 26056 6112 26108 6118
rect 26056 6054 26108 6060
rect 25964 5908 26016 5914
rect 25964 5850 26016 5856
rect 26068 5778 26096 6054
rect 24768 5772 24820 5778
rect 24768 5714 24820 5720
rect 25320 5772 25372 5778
rect 25320 5714 25372 5720
rect 26056 5772 26108 5778
rect 26056 5714 26108 5720
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 24780 5302 24808 5714
rect 24952 5568 25004 5574
rect 24952 5510 25004 5516
rect 24964 5370 24992 5510
rect 24952 5364 25004 5370
rect 24952 5306 25004 5312
rect 24584 5296 24636 5302
rect 24584 5238 24636 5244
rect 24768 5296 24820 5302
rect 24768 5238 24820 5244
rect 26252 5234 26280 6122
rect 26436 5846 26464 6326
rect 26424 5840 26476 5846
rect 26424 5782 26476 5788
rect 26240 5228 26292 5234
rect 26240 5170 26292 5176
rect 26528 5166 26556 8366
rect 26620 7886 26648 9540
rect 26700 9522 26752 9528
rect 27160 8288 27212 8294
rect 27160 8230 27212 8236
rect 27172 7886 27200 8230
rect 26608 7880 26660 7886
rect 26608 7822 26660 7828
rect 27160 7880 27212 7886
rect 27160 7822 27212 7828
rect 27264 6118 27292 10542
rect 27252 6112 27304 6118
rect 27252 6054 27304 6060
rect 27264 5846 27292 6054
rect 27252 5840 27304 5846
rect 27252 5782 27304 5788
rect 26976 5228 27028 5234
rect 26976 5170 27028 5176
rect 24032 5160 24084 5166
rect 24032 5102 24084 5108
rect 26516 5160 26568 5166
rect 26516 5102 26568 5108
rect 24044 4622 24072 5102
rect 25872 5024 25924 5030
rect 25872 4966 25924 4972
rect 24032 4616 24084 4622
rect 24032 4558 24084 4564
rect 25884 4554 25912 4966
rect 26988 4826 27016 5170
rect 26976 4820 27028 4826
rect 26976 4762 27028 4768
rect 25872 4548 25924 4554
rect 25872 4490 25924 4496
rect 23848 4480 23900 4486
rect 23848 4422 23900 4428
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 23572 4072 23624 4078
rect 23572 4014 23624 4020
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 27356 2446 27384 15846
rect 27448 14958 27476 16759
rect 27540 16046 27568 18686
rect 27712 18284 27764 18290
rect 27712 18226 27764 18232
rect 27724 17270 27752 18226
rect 27908 18154 27936 18770
rect 27896 18148 27948 18154
rect 27896 18090 27948 18096
rect 28080 17672 28132 17678
rect 28080 17614 28132 17620
rect 27988 17536 28040 17542
rect 27988 17478 28040 17484
rect 27712 17264 27764 17270
rect 27712 17206 27764 17212
rect 27894 17096 27950 17105
rect 27894 17031 27950 17040
rect 27712 16992 27764 16998
rect 27712 16934 27764 16940
rect 27724 16794 27752 16934
rect 27712 16788 27764 16794
rect 27712 16730 27764 16736
rect 27908 16726 27936 17031
rect 27896 16720 27948 16726
rect 27896 16662 27948 16668
rect 27620 16448 27672 16454
rect 27620 16390 27672 16396
rect 27804 16448 27856 16454
rect 27804 16390 27856 16396
rect 27632 16114 27660 16390
rect 27620 16108 27672 16114
rect 27620 16050 27672 16056
rect 27528 16040 27580 16046
rect 27528 15982 27580 15988
rect 27816 15178 27844 16390
rect 27896 16108 27948 16114
rect 27896 16050 27948 16056
rect 27908 15706 27936 16050
rect 27896 15700 27948 15706
rect 27896 15642 27948 15648
rect 27724 15150 27844 15178
rect 27436 14952 27488 14958
rect 27436 14894 27488 14900
rect 27620 13864 27672 13870
rect 27620 13806 27672 13812
rect 27632 13394 27660 13806
rect 27620 13388 27672 13394
rect 27620 13330 27672 13336
rect 27620 13252 27672 13258
rect 27620 13194 27672 13200
rect 27632 12238 27660 13194
rect 27620 12232 27672 12238
rect 27620 12174 27672 12180
rect 27528 10668 27580 10674
rect 27528 10610 27580 10616
rect 27540 9042 27568 10610
rect 27528 9036 27580 9042
rect 27528 8978 27580 8984
rect 27540 8634 27568 8978
rect 27528 8628 27580 8634
rect 27528 8570 27580 8576
rect 27436 6724 27488 6730
rect 27436 6666 27488 6672
rect 27448 6254 27476 6666
rect 27436 6248 27488 6254
rect 27436 6190 27488 6196
rect 27448 4622 27476 6190
rect 27436 4616 27488 4622
rect 27436 4558 27488 4564
rect 27724 3058 27752 15150
rect 27804 15020 27856 15026
rect 27804 14962 27856 14968
rect 27816 14618 27844 14962
rect 27896 14816 27948 14822
rect 27896 14758 27948 14764
rect 27804 14612 27856 14618
rect 27804 14554 27856 14560
rect 27804 14408 27856 14414
rect 27804 14350 27856 14356
rect 27816 13802 27844 14350
rect 27804 13796 27856 13802
rect 27804 13738 27856 13744
rect 27816 13326 27844 13738
rect 27804 13320 27856 13326
rect 27804 13262 27856 13268
rect 27816 12850 27844 13262
rect 27804 12844 27856 12850
rect 27804 12786 27856 12792
rect 27804 12640 27856 12646
rect 27802 12608 27804 12617
rect 27856 12608 27858 12617
rect 27802 12543 27858 12552
rect 27802 12336 27858 12345
rect 27802 12271 27858 12280
rect 27816 12102 27844 12271
rect 27804 12096 27856 12102
rect 27804 12038 27856 12044
rect 27908 8650 27936 14758
rect 28000 13938 28028 17478
rect 28092 17134 28120 17614
rect 28080 17128 28132 17134
rect 28080 17070 28132 17076
rect 28184 15502 28212 25638
rect 28448 25288 28500 25294
rect 28552 25276 28580 26386
rect 28644 25294 28672 26454
rect 28816 25832 28868 25838
rect 28816 25774 28868 25780
rect 28500 25248 28580 25276
rect 28632 25288 28684 25294
rect 28448 25230 28500 25236
rect 28632 25230 28684 25236
rect 28264 25152 28316 25158
rect 28264 25094 28316 25100
rect 28276 24993 28304 25094
rect 28262 24984 28318 24993
rect 28262 24919 28318 24928
rect 28540 24744 28592 24750
rect 28540 24686 28592 24692
rect 28264 24676 28316 24682
rect 28264 24618 28316 24624
rect 28276 23225 28304 24618
rect 28356 24132 28408 24138
rect 28356 24074 28408 24080
rect 28368 23526 28396 24074
rect 28552 24070 28580 24686
rect 28540 24064 28592 24070
rect 28540 24006 28592 24012
rect 28356 23520 28408 23526
rect 28552 23508 28580 24006
rect 28828 23866 28856 25774
rect 28920 25430 28948 26522
rect 29012 25838 29040 26930
rect 29000 25832 29052 25838
rect 29000 25774 29052 25780
rect 28908 25424 28960 25430
rect 28908 25366 28960 25372
rect 29000 25288 29052 25294
rect 29000 25230 29052 25236
rect 29012 24682 29040 25230
rect 29090 25120 29146 25129
rect 29090 25055 29146 25064
rect 29000 24676 29052 24682
rect 29000 24618 29052 24624
rect 28816 23860 28868 23866
rect 28816 23802 28868 23808
rect 28632 23792 28684 23798
rect 28684 23769 28764 23780
rect 28684 23760 28778 23769
rect 28684 23752 28722 23760
rect 28632 23734 28684 23740
rect 28722 23695 28778 23704
rect 28632 23520 28684 23526
rect 28552 23480 28632 23508
rect 28356 23462 28408 23468
rect 28954 23520 29006 23526
rect 28632 23462 28684 23468
rect 28828 23480 28954 23508
rect 28630 23352 28686 23361
rect 28630 23287 28686 23296
rect 28262 23216 28318 23225
rect 28262 23151 28318 23160
rect 28644 23118 28672 23287
rect 28632 23112 28684 23118
rect 28632 23054 28684 23060
rect 28724 23112 28776 23118
rect 28724 23054 28776 23060
rect 28540 22772 28592 22778
rect 28540 22714 28592 22720
rect 28262 22672 28318 22681
rect 28262 22607 28264 22616
rect 28316 22607 28318 22616
rect 28264 22578 28316 22584
rect 28552 22098 28580 22714
rect 28540 22092 28592 22098
rect 28540 22034 28592 22040
rect 28356 22024 28408 22030
rect 28356 21966 28408 21972
rect 28448 22024 28500 22030
rect 28448 21966 28500 21972
rect 28276 20398 28304 20429
rect 28264 20392 28316 20398
rect 28262 20360 28264 20369
rect 28316 20360 28318 20369
rect 28262 20295 28318 20304
rect 28276 20262 28304 20295
rect 28264 20256 28316 20262
rect 28264 20198 28316 20204
rect 28080 15496 28132 15502
rect 28080 15438 28132 15444
rect 28172 15496 28224 15502
rect 28172 15438 28224 15444
rect 28092 15026 28120 15438
rect 28080 15020 28132 15026
rect 28080 14962 28132 14968
rect 27988 13932 28040 13938
rect 27988 13874 28040 13880
rect 28172 13728 28224 13734
rect 28172 13670 28224 13676
rect 27988 12776 28040 12782
rect 27988 12718 28040 12724
rect 28000 12442 28028 12718
rect 27988 12436 28040 12442
rect 27988 12378 28040 12384
rect 28080 11008 28132 11014
rect 28080 10950 28132 10956
rect 28092 10810 28120 10950
rect 28080 10804 28132 10810
rect 28080 10746 28132 10752
rect 27988 9580 28040 9586
rect 27988 9522 28040 9528
rect 28000 9178 28028 9522
rect 27988 9172 28040 9178
rect 27988 9114 28040 9120
rect 27908 8622 28028 8650
rect 27896 8492 27948 8498
rect 27896 8434 27948 8440
rect 27908 8090 27936 8434
rect 27896 8084 27948 8090
rect 27896 8026 27948 8032
rect 27908 7886 27936 8026
rect 27896 7880 27948 7886
rect 27896 7822 27948 7828
rect 28000 5778 28028 8622
rect 28080 6316 28132 6322
rect 28080 6258 28132 6264
rect 28092 5914 28120 6258
rect 28080 5908 28132 5914
rect 28080 5850 28132 5856
rect 27988 5772 28040 5778
rect 27988 5714 28040 5720
rect 27896 4548 27948 4554
rect 27896 4490 27948 4496
rect 27908 4282 27936 4490
rect 28184 4486 28212 13670
rect 28276 13258 28304 20198
rect 28368 14414 28396 21966
rect 28460 20398 28488 21966
rect 28644 21894 28672 23054
rect 28632 21888 28684 21894
rect 28538 21856 28594 21865
rect 28632 21830 28684 21836
rect 28538 21791 28594 21800
rect 28552 21554 28580 21791
rect 28632 21616 28684 21622
rect 28632 21558 28684 21564
rect 28540 21548 28592 21554
rect 28540 21490 28592 21496
rect 28448 20392 28500 20398
rect 28448 20334 28500 20340
rect 28356 14408 28408 14414
rect 28356 14350 28408 14356
rect 28354 13696 28410 13705
rect 28354 13631 28410 13640
rect 28368 13326 28396 13631
rect 28356 13320 28408 13326
rect 28356 13262 28408 13268
rect 28264 13252 28316 13258
rect 28264 13194 28316 13200
rect 28262 12336 28318 12345
rect 28460 12306 28488 20334
rect 28644 19718 28672 21558
rect 28632 19712 28684 19718
rect 28632 19654 28684 19660
rect 28540 19168 28592 19174
rect 28540 19110 28592 19116
rect 28552 16697 28580 19110
rect 28736 18850 28764 23054
rect 28828 22273 28856 23480
rect 28954 23462 29006 23468
rect 28908 23112 28960 23118
rect 28908 23054 28960 23060
rect 28920 22642 28948 23054
rect 28908 22636 28960 22642
rect 28908 22578 28960 22584
rect 29000 22432 29052 22438
rect 29000 22374 29052 22380
rect 28814 22264 28870 22273
rect 28814 22199 28870 22208
rect 28816 22092 28868 22098
rect 28816 22034 28868 22040
rect 28828 20466 28856 22034
rect 28908 21072 28960 21078
rect 28908 21014 28960 21020
rect 28816 20460 28868 20466
rect 28816 20402 28868 20408
rect 28920 19394 28948 21014
rect 28828 19378 28948 19394
rect 28816 19372 28948 19378
rect 28868 19366 28948 19372
rect 29012 19357 29040 22374
rect 29104 21418 29132 25055
rect 29196 24070 29224 31282
rect 29288 27538 29316 34002
rect 29644 33992 29696 33998
rect 29644 33934 29696 33940
rect 30196 33992 30248 33998
rect 30196 33934 30248 33940
rect 29656 32434 29684 33934
rect 30012 33924 30064 33930
rect 30012 33866 30064 33872
rect 30104 33924 30156 33930
rect 30104 33866 30156 33872
rect 29828 33448 29880 33454
rect 29828 33390 29880 33396
rect 29840 32774 29868 33390
rect 29920 33380 29972 33386
rect 29920 33322 29972 33328
rect 29932 32910 29960 33322
rect 29920 32904 29972 32910
rect 29920 32846 29972 32852
rect 29828 32768 29880 32774
rect 29828 32710 29880 32716
rect 29644 32428 29696 32434
rect 29644 32370 29696 32376
rect 29656 30938 29684 32370
rect 29736 32360 29788 32366
rect 29736 32302 29788 32308
rect 29644 30932 29696 30938
rect 29644 30874 29696 30880
rect 29656 30258 29684 30874
rect 29644 30252 29696 30258
rect 29644 30194 29696 30200
rect 29368 30116 29420 30122
rect 29368 30058 29420 30064
rect 29380 29238 29408 30058
rect 29460 30048 29512 30054
rect 29460 29990 29512 29996
rect 29368 29232 29420 29238
rect 29366 29200 29368 29209
rect 29420 29200 29422 29209
rect 29366 29135 29422 29144
rect 29368 28960 29420 28966
rect 29368 28902 29420 28908
rect 29276 27532 29328 27538
rect 29276 27474 29328 27480
rect 29380 27334 29408 28902
rect 29368 27328 29420 27334
rect 29368 27270 29420 27276
rect 29276 24812 29328 24818
rect 29276 24754 29328 24760
rect 29288 24206 29316 24754
rect 29276 24200 29328 24206
rect 29276 24142 29328 24148
rect 29184 24064 29236 24070
rect 29184 24006 29236 24012
rect 29288 23118 29316 24142
rect 29276 23112 29328 23118
rect 29276 23054 29328 23060
rect 29380 22760 29408 27270
rect 29472 23866 29500 29990
rect 29656 29646 29684 30194
rect 29644 29640 29696 29646
rect 29644 29582 29696 29588
rect 29552 29572 29604 29578
rect 29552 29514 29604 29520
rect 29564 29073 29592 29514
rect 29656 29170 29684 29582
rect 29644 29164 29696 29170
rect 29644 29106 29696 29112
rect 29550 29064 29606 29073
rect 29550 28999 29606 29008
rect 29656 28082 29684 29106
rect 29644 28076 29696 28082
rect 29644 28018 29696 28024
rect 29748 27614 29776 32302
rect 29932 28150 29960 32846
rect 30024 32756 30052 33866
rect 30116 33833 30144 33866
rect 30102 33824 30158 33833
rect 30102 33759 30158 33768
rect 30208 33046 30236 33934
rect 30668 33114 30696 35022
rect 31024 35022 31076 35028
rect 31668 35080 31720 35086
rect 31668 35022 31720 35028
rect 31760 35080 31812 35086
rect 31760 35022 31812 35028
rect 31944 35080 31996 35086
rect 32048 35068 32076 35702
rect 32128 35148 32180 35154
rect 32128 35090 32180 35096
rect 31996 35040 32076 35068
rect 31944 35022 31996 35028
rect 30746 34983 30802 34992
rect 30760 34746 30788 34983
rect 31116 34944 31168 34950
rect 31116 34886 31168 34892
rect 30748 34740 30800 34746
rect 30748 34682 30800 34688
rect 30748 34400 30800 34406
rect 30748 34342 30800 34348
rect 30760 33454 30788 34342
rect 31128 33930 31156 34886
rect 31390 34096 31446 34105
rect 31390 34031 31446 34040
rect 31208 33992 31260 33998
rect 31300 33992 31352 33998
rect 31208 33934 31260 33940
rect 31298 33960 31300 33969
rect 31352 33960 31354 33969
rect 31116 33924 31168 33930
rect 30944 33884 31116 33912
rect 30944 33590 30972 33884
rect 31116 33866 31168 33872
rect 31116 33652 31168 33658
rect 31116 33594 31168 33600
rect 30932 33584 30984 33590
rect 30932 33526 30984 33532
rect 30748 33448 30800 33454
rect 30746 33416 30748 33425
rect 30800 33416 30802 33425
rect 30746 33351 30802 33360
rect 30656 33108 30708 33114
rect 30656 33050 30708 33056
rect 30196 33040 30248 33046
rect 30196 32982 30248 32988
rect 30104 32904 30156 32910
rect 30102 32872 30104 32881
rect 30380 32904 30432 32910
rect 30156 32872 30158 32881
rect 30102 32807 30158 32816
rect 30208 32864 30380 32892
rect 30104 32768 30156 32774
rect 30024 32736 30104 32756
rect 30156 32736 30158 32745
rect 30024 32728 30102 32736
rect 30102 32671 30158 32680
rect 30116 32502 30144 32671
rect 30104 32496 30156 32502
rect 30104 32438 30156 32444
rect 30012 30252 30064 30258
rect 30116 30240 30144 32438
rect 30208 32434 30236 32864
rect 30380 32846 30432 32852
rect 30288 32768 30340 32774
rect 30288 32710 30340 32716
rect 30196 32428 30248 32434
rect 30196 32370 30248 32376
rect 30300 32416 30328 32710
rect 30380 32428 30432 32434
rect 30300 32388 30380 32416
rect 30196 30660 30248 30666
rect 30196 30602 30248 30608
rect 30064 30212 30144 30240
rect 30012 30194 30064 30200
rect 30116 29646 30144 30212
rect 30012 29640 30064 29646
rect 30012 29582 30064 29588
rect 30104 29640 30156 29646
rect 30104 29582 30156 29588
rect 30024 28626 30052 29582
rect 30012 28620 30064 28626
rect 30012 28562 30064 28568
rect 30024 28422 30052 28562
rect 30012 28416 30064 28422
rect 30012 28358 30064 28364
rect 30116 28218 30144 29582
rect 30208 28762 30236 30602
rect 30300 30258 30328 32388
rect 30380 32370 30432 32376
rect 30748 31476 30800 31482
rect 30748 31418 30800 31424
rect 30564 31408 30616 31414
rect 30564 31350 30616 31356
rect 30470 30968 30526 30977
rect 30470 30903 30526 30912
rect 30484 30258 30512 30903
rect 30288 30252 30340 30258
rect 30288 30194 30340 30200
rect 30472 30252 30524 30258
rect 30472 30194 30524 30200
rect 30300 29628 30328 30194
rect 30380 30116 30432 30122
rect 30380 30058 30432 30064
rect 30392 30025 30420 30058
rect 30378 30016 30434 30025
rect 30378 29951 30434 29960
rect 30380 29640 30432 29646
rect 30300 29600 30380 29628
rect 30380 29582 30432 29588
rect 30392 29209 30420 29582
rect 30576 29306 30604 31350
rect 30760 31346 30788 31418
rect 30944 31346 30972 33526
rect 31024 33516 31076 33522
rect 31024 33458 31076 33464
rect 31036 32570 31064 33458
rect 31024 32564 31076 32570
rect 31024 32506 31076 32512
rect 30656 31340 30708 31346
rect 30656 31282 30708 31288
rect 30748 31340 30800 31346
rect 30748 31282 30800 31288
rect 30932 31340 30984 31346
rect 30932 31282 30984 31288
rect 30668 30394 30696 31282
rect 30760 31249 30788 31282
rect 30746 31240 30802 31249
rect 30746 31175 30802 31184
rect 30748 30728 30800 30734
rect 30748 30670 30800 30676
rect 30840 30728 30892 30734
rect 30840 30670 30892 30676
rect 30656 30388 30708 30394
rect 30656 30330 30708 30336
rect 30760 29850 30788 30670
rect 30852 30394 30880 30670
rect 30944 30666 30972 31282
rect 31128 30938 31156 33594
rect 31220 33114 31248 33934
rect 31298 33895 31354 33904
rect 31404 33590 31432 34031
rect 31680 33998 31708 35022
rect 31772 34202 31800 35022
rect 31852 34944 31904 34950
rect 31852 34886 31904 34892
rect 31864 34202 31892 34886
rect 31760 34196 31812 34202
rect 31760 34138 31812 34144
rect 31852 34196 31904 34202
rect 31852 34138 31904 34144
rect 31944 34128 31996 34134
rect 31864 34076 31944 34082
rect 31864 34070 31996 34076
rect 31864 34054 31984 34070
rect 31668 33992 31720 33998
rect 31496 33940 31668 33946
rect 31496 33934 31720 33940
rect 31496 33918 31708 33934
rect 31392 33584 31444 33590
rect 31392 33526 31444 33532
rect 31496 33522 31524 33918
rect 31484 33516 31536 33522
rect 31484 33458 31536 33464
rect 31496 33402 31524 33458
rect 31404 33374 31524 33402
rect 31208 33108 31260 33114
rect 31208 33050 31260 33056
rect 31300 32904 31352 32910
rect 31220 32864 31300 32892
rect 31220 32434 31248 32864
rect 31300 32846 31352 32852
rect 31300 32768 31352 32774
rect 31298 32736 31300 32745
rect 31352 32736 31354 32745
rect 31298 32671 31354 32680
rect 31208 32428 31260 32434
rect 31208 32370 31260 32376
rect 31404 32230 31432 33374
rect 31484 32972 31536 32978
rect 31484 32914 31536 32920
rect 31392 32224 31444 32230
rect 31392 32166 31444 32172
rect 31116 30932 31168 30938
rect 31116 30874 31168 30880
rect 30932 30660 30984 30666
rect 30932 30602 30984 30608
rect 31116 30660 31168 30666
rect 31116 30602 31168 30608
rect 31128 30410 31156 30602
rect 31392 30592 31444 30598
rect 31392 30534 31444 30540
rect 30840 30388 30892 30394
rect 30840 30330 30892 30336
rect 30944 30382 31156 30410
rect 30748 29844 30800 29850
rect 30748 29786 30800 29792
rect 30656 29776 30708 29782
rect 30656 29718 30708 29724
rect 30668 29510 30696 29718
rect 30656 29504 30708 29510
rect 30656 29446 30708 29452
rect 30564 29300 30616 29306
rect 30564 29242 30616 29248
rect 30472 29232 30524 29238
rect 30378 29200 30434 29209
rect 30472 29174 30524 29180
rect 30378 29135 30434 29144
rect 30196 28756 30248 28762
rect 30196 28698 30248 28704
rect 30392 28558 30420 29135
rect 30484 28626 30512 29174
rect 30472 28620 30524 28626
rect 30472 28562 30524 28568
rect 30380 28552 30432 28558
rect 30380 28494 30432 28500
rect 30104 28212 30156 28218
rect 30104 28154 30156 28160
rect 29920 28144 29972 28150
rect 29920 28086 29972 28092
rect 30012 28076 30064 28082
rect 30012 28018 30064 28024
rect 29656 27586 29776 27614
rect 29656 25226 29684 27586
rect 30024 27334 30052 28018
rect 30116 27538 30144 28154
rect 30196 28076 30248 28082
rect 30196 28018 30248 28024
rect 30104 27532 30156 27538
rect 30104 27474 30156 27480
rect 29736 27328 29788 27334
rect 29736 27270 29788 27276
rect 30012 27328 30064 27334
rect 30012 27270 30064 27276
rect 29748 26353 29776 27270
rect 30102 27024 30158 27033
rect 30102 26959 30158 26968
rect 29734 26344 29790 26353
rect 29734 26279 29790 26288
rect 29920 25492 29972 25498
rect 29920 25434 29972 25440
rect 29644 25220 29696 25226
rect 29644 25162 29696 25168
rect 29644 24812 29696 24818
rect 29644 24754 29696 24760
rect 29552 24064 29604 24070
rect 29552 24006 29604 24012
rect 29460 23860 29512 23866
rect 29460 23802 29512 23808
rect 29564 23236 29592 24006
rect 29656 23662 29684 24754
rect 29828 24676 29880 24682
rect 29828 24618 29880 24624
rect 29736 24608 29788 24614
rect 29736 24550 29788 24556
rect 29644 23656 29696 23662
rect 29644 23598 29696 23604
rect 29472 23208 29592 23236
rect 29472 22982 29500 23208
rect 29656 23186 29684 23598
rect 29644 23180 29696 23186
rect 29644 23122 29696 23128
rect 29460 22976 29512 22982
rect 29460 22918 29512 22924
rect 29380 22732 29500 22760
rect 29366 22672 29422 22681
rect 29366 22607 29368 22616
rect 29420 22607 29422 22616
rect 29368 22578 29420 22584
rect 29380 21729 29408 22578
rect 29472 22574 29500 22732
rect 29748 22642 29776 24550
rect 29840 24274 29868 24618
rect 29828 24268 29880 24274
rect 29828 24210 29880 24216
rect 29932 23730 29960 25434
rect 30012 24812 30064 24818
rect 30012 24754 30064 24760
rect 30024 24138 30052 24754
rect 30012 24132 30064 24138
rect 30012 24074 30064 24080
rect 29920 23724 29972 23730
rect 29920 23666 29972 23672
rect 29828 23656 29880 23662
rect 29828 23598 29880 23604
rect 29840 23118 29868 23598
rect 29932 23186 29960 23666
rect 30012 23588 30064 23594
rect 30012 23530 30064 23536
rect 29920 23180 29972 23186
rect 29920 23122 29972 23128
rect 30024 23118 30052 23530
rect 29828 23112 29880 23118
rect 29828 23054 29880 23060
rect 30012 23112 30064 23118
rect 30012 23054 30064 23060
rect 29840 22778 29868 23054
rect 29920 22976 29972 22982
rect 30116 22964 30144 26959
rect 30208 26897 30236 28018
rect 30380 28008 30432 28014
rect 30380 27950 30432 27956
rect 30392 27606 30420 27950
rect 30380 27600 30432 27606
rect 30380 27542 30432 27548
rect 30288 27396 30340 27402
rect 30392 27384 30420 27542
rect 30484 27470 30512 28562
rect 30564 28552 30616 28558
rect 30564 28494 30616 28500
rect 30576 28082 30604 28494
rect 30564 28076 30616 28082
rect 30564 28018 30616 28024
rect 30472 27464 30524 27470
rect 30472 27406 30524 27412
rect 30340 27356 30420 27384
rect 30288 27338 30340 27344
rect 30194 26888 30250 26897
rect 30194 26823 30250 26832
rect 30208 26586 30236 26823
rect 30196 26580 30248 26586
rect 30196 26522 30248 26528
rect 30300 26296 30328 27338
rect 30380 26920 30432 26926
rect 30380 26862 30432 26868
rect 29920 22918 29972 22924
rect 30024 22936 30144 22964
rect 30208 26268 30328 26296
rect 29828 22772 29880 22778
rect 29828 22714 29880 22720
rect 29736 22636 29788 22642
rect 29736 22578 29788 22584
rect 29460 22568 29512 22574
rect 29460 22510 29512 22516
rect 29460 22092 29512 22098
rect 29460 22034 29512 22040
rect 29366 21720 29422 21729
rect 29366 21655 29422 21664
rect 29092 21412 29144 21418
rect 29092 21354 29144 21360
rect 29276 20528 29328 20534
rect 29276 20470 29328 20476
rect 29184 20392 29236 20398
rect 29184 20334 29236 20340
rect 29196 19854 29224 20334
rect 29288 20058 29316 20470
rect 29368 20460 29420 20466
rect 29368 20402 29420 20408
rect 29276 20052 29328 20058
rect 29276 19994 29328 20000
rect 29184 19848 29236 19854
rect 29184 19790 29236 19796
rect 29276 19780 29328 19786
rect 29276 19722 29328 19728
rect 29288 19378 29316 19722
rect 29276 19372 29328 19378
rect 28816 19314 28868 19320
rect 28998 19348 29054 19357
rect 28644 18822 28764 18850
rect 28538 16688 28594 16697
rect 28538 16623 28594 16632
rect 28644 15502 28672 18822
rect 28724 18692 28776 18698
rect 28724 18634 28776 18640
rect 28736 18222 28764 18634
rect 28724 18216 28776 18222
rect 28724 18158 28776 18164
rect 28724 17808 28776 17814
rect 28724 17750 28776 17756
rect 28736 17270 28764 17750
rect 28724 17264 28776 17270
rect 28722 17232 28724 17241
rect 28776 17232 28778 17241
rect 28722 17167 28778 17176
rect 28724 17128 28776 17134
rect 28828 17116 28856 19314
rect 28908 19304 28960 19310
rect 29276 19314 29328 19320
rect 28998 19283 29054 19292
rect 28908 19246 28960 19252
rect 28920 18902 28948 19246
rect 29184 19168 29236 19174
rect 29184 19110 29236 19116
rect 28998 19000 29054 19009
rect 29196 18970 29224 19110
rect 28998 18935 29054 18944
rect 29184 18964 29236 18970
rect 28908 18896 28960 18902
rect 28908 18838 28960 18844
rect 28776 17088 28856 17116
rect 28724 17070 28776 17076
rect 28632 15496 28684 15502
rect 28632 15438 28684 15444
rect 28644 13870 28672 15438
rect 28736 15366 28764 17070
rect 28906 16824 28962 16833
rect 28906 16759 28908 16768
rect 28960 16759 28962 16768
rect 28908 16730 28960 16736
rect 28906 16688 28962 16697
rect 28906 16623 28962 16632
rect 28920 16590 28948 16623
rect 28908 16584 28960 16590
rect 28908 16526 28960 16532
rect 28908 16448 28960 16454
rect 28906 16416 28908 16425
rect 28960 16416 28962 16425
rect 28906 16351 28962 16360
rect 29012 16046 29040 18935
rect 29184 18906 29236 18912
rect 29380 18766 29408 20402
rect 29472 20262 29500 22034
rect 29736 21344 29788 21350
rect 29736 21286 29788 21292
rect 29642 20496 29698 20505
rect 29642 20431 29644 20440
rect 29696 20431 29698 20440
rect 29644 20402 29696 20408
rect 29460 20256 29512 20262
rect 29460 20198 29512 20204
rect 29748 19854 29776 21286
rect 29932 20942 29960 22918
rect 29920 20936 29972 20942
rect 29920 20878 29972 20884
rect 29828 20800 29880 20806
rect 29828 20742 29880 20748
rect 29840 19922 29868 20742
rect 29932 20398 29960 20878
rect 29920 20392 29972 20398
rect 29920 20334 29972 20340
rect 29828 19916 29880 19922
rect 29828 19858 29880 19864
rect 29460 19848 29512 19854
rect 29460 19790 29512 19796
rect 29736 19848 29788 19854
rect 29736 19790 29788 19796
rect 29368 18760 29420 18766
rect 29368 18702 29420 18708
rect 29092 18148 29144 18154
rect 29092 18090 29144 18096
rect 29104 17882 29132 18090
rect 29092 17876 29144 17882
rect 29092 17818 29144 17824
rect 29184 17264 29236 17270
rect 29184 17206 29236 17212
rect 29196 16946 29224 17206
rect 29104 16918 29224 16946
rect 29276 16992 29328 16998
rect 29276 16934 29328 16940
rect 29104 16658 29132 16918
rect 29092 16652 29144 16658
rect 29092 16594 29144 16600
rect 29000 16040 29052 16046
rect 29000 15982 29052 15988
rect 28724 15360 28776 15366
rect 28724 15302 28776 15308
rect 29104 14958 29132 16594
rect 29184 16584 29236 16590
rect 29184 16526 29236 16532
rect 29092 14952 29144 14958
rect 29092 14894 29144 14900
rect 29000 14884 29052 14890
rect 29000 14826 29052 14832
rect 28816 14612 28868 14618
rect 28816 14554 28868 14560
rect 28828 13938 28856 14554
rect 29012 14278 29040 14826
rect 29000 14272 29052 14278
rect 29000 14214 29052 14220
rect 28816 13932 28868 13938
rect 28816 13874 28868 13880
rect 28632 13864 28684 13870
rect 28632 13806 28684 13812
rect 28644 13258 28672 13806
rect 28828 13462 28856 13874
rect 29196 13734 29224 16526
rect 29288 16114 29316 16934
rect 29472 16658 29500 19790
rect 29552 19712 29604 19718
rect 29552 19654 29604 19660
rect 29460 16652 29512 16658
rect 29460 16594 29512 16600
rect 29276 16108 29328 16114
rect 29276 16050 29328 16056
rect 29460 16108 29512 16114
rect 29460 16050 29512 16056
rect 29276 15904 29328 15910
rect 29276 15846 29328 15852
rect 29184 13728 29236 13734
rect 29090 13696 29146 13705
rect 29184 13670 29236 13676
rect 29090 13631 29146 13640
rect 28816 13456 28868 13462
rect 28816 13398 28868 13404
rect 29000 13388 29052 13394
rect 29000 13330 29052 13336
rect 28632 13252 28684 13258
rect 28632 13194 28684 13200
rect 28262 12271 28318 12280
rect 28448 12300 28500 12306
rect 28276 12238 28304 12271
rect 28448 12242 28500 12248
rect 28644 12238 28672 13194
rect 28816 12776 28868 12782
rect 28816 12718 28868 12724
rect 28828 12306 28856 12718
rect 29012 12442 29040 13330
rect 29104 12918 29132 13631
rect 29092 12912 29144 12918
rect 29092 12854 29144 12860
rect 29196 12850 29224 13670
rect 29184 12844 29236 12850
rect 29184 12786 29236 12792
rect 29000 12436 29052 12442
rect 29288 12434 29316 15846
rect 29472 15706 29500 16050
rect 29460 15700 29512 15706
rect 29460 15642 29512 15648
rect 29288 12406 29408 12434
rect 29000 12378 29052 12384
rect 28816 12300 28868 12306
rect 28816 12242 28868 12248
rect 28264 12232 28316 12238
rect 28264 12174 28316 12180
rect 28632 12232 28684 12238
rect 28632 12174 28684 12180
rect 28908 12232 28960 12238
rect 28908 12174 28960 12180
rect 28264 12096 28316 12102
rect 28264 12038 28316 12044
rect 28276 5710 28304 12038
rect 28920 11286 28948 12174
rect 29000 11552 29052 11558
rect 29000 11494 29052 11500
rect 28908 11280 28960 11286
rect 28908 11222 28960 11228
rect 29012 10742 29040 11494
rect 29184 11144 29236 11150
rect 29184 11086 29236 11092
rect 29000 10736 29052 10742
rect 29000 10678 29052 10684
rect 29196 9654 29224 11086
rect 29184 9648 29236 9654
rect 29184 9590 29236 9596
rect 28356 9444 28408 9450
rect 28356 9386 28408 9392
rect 28368 8974 28396 9386
rect 28356 8968 28408 8974
rect 28356 8910 28408 8916
rect 28448 8832 28500 8838
rect 28448 8774 28500 8780
rect 28460 8566 28488 8774
rect 29184 8628 29236 8634
rect 29184 8570 29236 8576
rect 28448 8560 28500 8566
rect 28448 8502 28500 8508
rect 29196 8498 29224 8570
rect 29184 8492 29236 8498
rect 29184 8434 29236 8440
rect 28356 8424 28408 8430
rect 28356 8366 28408 8372
rect 28368 7818 28396 8366
rect 28356 7812 28408 7818
rect 28356 7754 28408 7760
rect 28368 6866 28396 7754
rect 29196 7478 29224 8434
rect 29184 7472 29236 7478
rect 29184 7414 29236 7420
rect 29092 7200 29144 7206
rect 29092 7142 29144 7148
rect 28356 6860 28408 6866
rect 28356 6802 28408 6808
rect 28448 6384 28500 6390
rect 28448 6326 28500 6332
rect 28356 5772 28408 5778
rect 28356 5714 28408 5720
rect 28264 5704 28316 5710
rect 28264 5646 28316 5652
rect 28368 5302 28396 5714
rect 28460 5710 28488 6326
rect 29104 6322 29132 7142
rect 29196 6662 29224 7414
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 29184 6656 29236 6662
rect 29184 6598 29236 6604
rect 29288 6458 29316 6734
rect 29276 6452 29328 6458
rect 29276 6394 29328 6400
rect 29092 6316 29144 6322
rect 29092 6258 29144 6264
rect 28448 5704 28500 5710
rect 28448 5646 28500 5652
rect 28356 5296 28408 5302
rect 28356 5238 28408 5244
rect 28172 4480 28224 4486
rect 28172 4422 28224 4428
rect 27896 4276 27948 4282
rect 27896 4218 27948 4224
rect 28368 4146 28396 5238
rect 29000 4820 29052 4826
rect 29000 4762 29052 4768
rect 29012 4282 29040 4762
rect 29000 4276 29052 4282
rect 29000 4218 29052 4224
rect 28356 4140 28408 4146
rect 28356 4082 28408 4088
rect 29380 3942 29408 12406
rect 29564 9178 29592 19654
rect 30024 19514 30052 22936
rect 30104 22772 30156 22778
rect 30104 22714 30156 22720
rect 30116 20466 30144 22714
rect 30208 21078 30236 26268
rect 30286 23488 30342 23497
rect 30286 23423 30342 23432
rect 30196 21072 30248 21078
rect 30196 21014 30248 21020
rect 30104 20460 30156 20466
rect 30104 20402 30156 20408
rect 30300 19938 30328 23423
rect 30392 20074 30420 26862
rect 30484 24614 30512 27406
rect 30668 26994 30696 29446
rect 30748 29232 30800 29238
rect 30748 29174 30800 29180
rect 30656 26988 30708 26994
rect 30656 26930 30708 26936
rect 30564 26240 30616 26246
rect 30564 26182 30616 26188
rect 30576 25226 30604 26182
rect 30564 25220 30616 25226
rect 30564 25162 30616 25168
rect 30668 24698 30696 26930
rect 30760 26790 30788 29174
rect 30748 26784 30800 26790
rect 30748 26726 30800 26732
rect 30576 24670 30696 24698
rect 30472 24608 30524 24614
rect 30472 24550 30524 24556
rect 30484 22642 30512 24550
rect 30576 24274 30604 24670
rect 30564 24268 30616 24274
rect 30564 24210 30616 24216
rect 30656 23656 30708 23662
rect 30656 23598 30708 23604
rect 30472 22636 30524 22642
rect 30472 22578 30524 22584
rect 30668 21894 30696 23598
rect 30760 22778 30788 26726
rect 30748 22772 30800 22778
rect 30748 22714 30800 22720
rect 30852 22710 30880 30330
rect 30944 28490 30972 30382
rect 31404 30326 31432 30534
rect 31024 30320 31076 30326
rect 31022 30288 31024 30297
rect 31392 30320 31444 30326
rect 31076 30288 31078 30297
rect 31392 30262 31444 30268
rect 31022 30223 31078 30232
rect 31116 30252 31168 30258
rect 31116 30194 31168 30200
rect 31300 30252 31352 30258
rect 31300 30194 31352 30200
rect 31024 30184 31076 30190
rect 31024 30126 31076 30132
rect 31036 29753 31064 30126
rect 31022 29744 31078 29753
rect 31022 29679 31078 29688
rect 31024 29572 31076 29578
rect 31024 29514 31076 29520
rect 30932 28484 30984 28490
rect 30932 28426 30984 28432
rect 30932 27464 30984 27470
rect 30932 27406 30984 27412
rect 30944 27334 30972 27406
rect 30932 27328 30984 27334
rect 30932 27270 30984 27276
rect 30944 26246 30972 27270
rect 30932 26240 30984 26246
rect 30932 26182 30984 26188
rect 31036 25974 31064 29514
rect 31128 28218 31156 30194
rect 31312 29170 31340 30194
rect 31404 30054 31432 30262
rect 31392 30048 31444 30054
rect 31392 29990 31444 29996
rect 31300 29164 31352 29170
rect 31300 29106 31352 29112
rect 31300 28552 31352 28558
rect 31300 28494 31352 28500
rect 31392 28552 31444 28558
rect 31392 28494 31444 28500
rect 31116 28212 31168 28218
rect 31116 28154 31168 28160
rect 31208 28076 31260 28082
rect 31208 28018 31260 28024
rect 31220 27538 31248 28018
rect 31312 27674 31340 28494
rect 31404 27946 31432 28494
rect 31392 27940 31444 27946
rect 31392 27882 31444 27888
rect 31300 27668 31352 27674
rect 31300 27610 31352 27616
rect 31208 27532 31260 27538
rect 31208 27474 31260 27480
rect 31208 27396 31260 27402
rect 31208 27338 31260 27344
rect 31220 26994 31248 27338
rect 31208 26988 31260 26994
rect 31208 26930 31260 26936
rect 31392 26988 31444 26994
rect 31392 26930 31444 26936
rect 31300 26240 31352 26246
rect 31300 26182 31352 26188
rect 31024 25968 31076 25974
rect 31024 25910 31076 25916
rect 31312 25158 31340 26182
rect 31300 25152 31352 25158
rect 31300 25094 31352 25100
rect 31312 24410 31340 25094
rect 31300 24404 31352 24410
rect 31300 24346 31352 24352
rect 31300 23860 31352 23866
rect 31300 23802 31352 23808
rect 31022 23760 31078 23769
rect 31022 23695 31078 23704
rect 30932 22976 30984 22982
rect 30932 22918 30984 22924
rect 30840 22704 30892 22710
rect 30840 22646 30892 22652
rect 30748 22568 30800 22574
rect 30748 22510 30800 22516
rect 30656 21888 30708 21894
rect 30656 21830 30708 21836
rect 30760 21554 30788 22510
rect 30944 22030 30972 22918
rect 30932 22024 30984 22030
rect 30932 21966 30984 21972
rect 30472 21548 30524 21554
rect 30472 21490 30524 21496
rect 30748 21548 30800 21554
rect 30748 21490 30800 21496
rect 30484 21146 30512 21490
rect 30564 21480 30616 21486
rect 30564 21422 30616 21428
rect 30472 21140 30524 21146
rect 30472 21082 30524 21088
rect 30392 20046 30512 20074
rect 30300 19922 30420 19938
rect 30300 19916 30432 19922
rect 30300 19910 30380 19916
rect 30380 19858 30432 19864
rect 30288 19780 30340 19786
rect 30288 19722 30340 19728
rect 30012 19508 30064 19514
rect 30012 19450 30064 19456
rect 30300 19378 30328 19722
rect 29828 19372 29880 19378
rect 29828 19314 29880 19320
rect 30012 19372 30064 19378
rect 30012 19314 30064 19320
rect 30288 19372 30340 19378
rect 30288 19314 30340 19320
rect 29736 19168 29788 19174
rect 29736 19110 29788 19116
rect 29748 18970 29776 19110
rect 29736 18964 29788 18970
rect 29736 18906 29788 18912
rect 29840 18902 29868 19314
rect 29828 18896 29880 18902
rect 29828 18838 29880 18844
rect 29840 17678 29868 18838
rect 30024 18834 30052 19314
rect 30288 19168 30340 19174
rect 30288 19110 30340 19116
rect 30012 18828 30064 18834
rect 30012 18770 30064 18776
rect 30012 18692 30064 18698
rect 30012 18634 30064 18640
rect 29828 17672 29880 17678
rect 29828 17614 29880 17620
rect 29918 17640 29974 17649
rect 29736 17536 29788 17542
rect 29736 17478 29788 17484
rect 29748 16697 29776 17478
rect 29734 16688 29790 16697
rect 29734 16623 29790 16632
rect 29840 16182 29868 17614
rect 29918 17575 29974 17584
rect 29932 17542 29960 17575
rect 29920 17536 29972 17542
rect 29920 17478 29972 17484
rect 29828 16176 29880 16182
rect 29828 16118 29880 16124
rect 29840 15502 29868 16118
rect 29736 15496 29788 15502
rect 29736 15438 29788 15444
rect 29828 15496 29880 15502
rect 29828 15438 29880 15444
rect 29748 12986 29776 15438
rect 29932 14498 29960 17478
rect 30024 17202 30052 18634
rect 30300 17882 30328 19110
rect 30484 18902 30512 20046
rect 30472 18896 30524 18902
rect 30472 18838 30524 18844
rect 30576 18290 30604 21422
rect 30840 21004 30892 21010
rect 30840 20946 30892 20952
rect 30656 20868 30708 20874
rect 30656 20810 30708 20816
rect 30668 20398 30696 20810
rect 30656 20392 30708 20398
rect 30656 20334 30708 20340
rect 30656 20256 30708 20262
rect 30656 20198 30708 20204
rect 30668 18358 30696 20198
rect 30748 19984 30800 19990
rect 30748 19926 30800 19932
rect 30760 19378 30788 19926
rect 30748 19372 30800 19378
rect 30748 19314 30800 19320
rect 30852 18766 30880 20946
rect 31036 19718 31064 23695
rect 31312 23186 31340 23802
rect 31404 23798 31432 26930
rect 31392 23792 31444 23798
rect 31392 23734 31444 23740
rect 31300 23180 31352 23186
rect 31300 23122 31352 23128
rect 31208 22636 31260 22642
rect 31208 22578 31260 22584
rect 31220 22234 31248 22578
rect 31208 22228 31260 22234
rect 31208 22170 31260 22176
rect 31116 22024 31168 22030
rect 31116 21966 31168 21972
rect 31128 21026 31156 21966
rect 31220 21554 31248 22170
rect 31312 22098 31340 23122
rect 31300 22092 31352 22098
rect 31300 22034 31352 22040
rect 31312 21842 31340 22034
rect 31404 21894 31432 23734
rect 31496 22506 31524 32914
rect 31760 32836 31812 32842
rect 31760 32778 31812 32784
rect 31668 32496 31720 32502
rect 31666 32464 31668 32473
rect 31720 32464 31722 32473
rect 31666 32399 31722 32408
rect 31576 32224 31628 32230
rect 31576 32166 31628 32172
rect 31588 31346 31616 32166
rect 31772 31385 31800 32778
rect 31864 31754 31892 34054
rect 31944 32904 31996 32910
rect 31942 32872 31944 32881
rect 31996 32872 31998 32881
rect 32048 32858 32076 35040
rect 32140 32978 32168 35090
rect 32324 35018 32352 36246
rect 32588 36168 32640 36174
rect 32588 36110 32640 36116
rect 32600 35290 32628 36110
rect 32680 35692 32732 35698
rect 32680 35634 32732 35640
rect 32588 35284 32640 35290
rect 32588 35226 32640 35232
rect 32312 35012 32364 35018
rect 32312 34954 32364 34960
rect 32692 34950 32720 35634
rect 32680 34944 32732 34950
rect 32680 34886 32732 34892
rect 32680 33856 32732 33862
rect 32680 33798 32732 33804
rect 32692 33590 32720 33798
rect 32680 33584 32732 33590
rect 32680 33526 32732 33532
rect 32128 32972 32180 32978
rect 32128 32914 32180 32920
rect 32312 32904 32364 32910
rect 32048 32830 32168 32858
rect 32312 32846 32364 32852
rect 31942 32807 31998 32816
rect 32140 31754 32168 32830
rect 32324 32570 32352 32846
rect 32312 32564 32364 32570
rect 32312 32506 32364 32512
rect 32324 32298 32352 32506
rect 32784 32366 32812 36790
rect 33692 36576 33744 36582
rect 33692 36518 33744 36524
rect 32956 35692 33008 35698
rect 32956 35634 33008 35640
rect 33048 35692 33100 35698
rect 33048 35634 33100 35640
rect 32864 35284 32916 35290
rect 32864 35226 32916 35232
rect 32876 34542 32904 35226
rect 32968 35018 32996 35634
rect 33060 35290 33088 35634
rect 33048 35284 33100 35290
rect 33048 35226 33100 35232
rect 32956 35012 33008 35018
rect 32956 34954 33008 34960
rect 32968 34610 32996 34954
rect 33704 34746 33732 36518
rect 33796 36378 33824 37198
rect 33968 37120 34020 37126
rect 33968 37062 34020 37068
rect 33980 36854 34008 37062
rect 33968 36848 34020 36854
rect 33968 36790 34020 36796
rect 34244 36712 34296 36718
rect 34244 36654 34296 36660
rect 33784 36372 33836 36378
rect 33784 36314 33836 36320
rect 34256 36242 34284 36654
rect 34244 36236 34296 36242
rect 34244 36178 34296 36184
rect 33784 36168 33836 36174
rect 33784 36110 33836 36116
rect 33796 35698 33824 36110
rect 33784 35692 33836 35698
rect 33784 35634 33836 35640
rect 33796 35290 33824 35634
rect 33784 35284 33836 35290
rect 33784 35226 33836 35232
rect 33692 34740 33744 34746
rect 33692 34682 33744 34688
rect 32956 34604 33008 34610
rect 32956 34546 33008 34552
rect 32864 34536 32916 34542
rect 32864 34478 32916 34484
rect 32876 33658 32904 34478
rect 32864 33652 32916 33658
rect 32864 33594 32916 33600
rect 32864 33516 32916 33522
rect 32864 33458 32916 33464
rect 32876 33114 32904 33458
rect 32864 33108 32916 33114
rect 32864 33050 32916 33056
rect 32864 32428 32916 32434
rect 32864 32370 32916 32376
rect 32588 32360 32640 32366
rect 32588 32302 32640 32308
rect 32772 32360 32824 32366
rect 32772 32302 32824 32308
rect 32312 32292 32364 32298
rect 32312 32234 32364 32240
rect 32496 31816 32548 31822
rect 32496 31758 32548 31764
rect 31864 31726 31984 31754
rect 31758 31376 31814 31385
rect 31576 31340 31628 31346
rect 31758 31311 31814 31320
rect 31576 31282 31628 31288
rect 31588 30734 31616 31282
rect 31576 30728 31628 30734
rect 31576 30670 31628 30676
rect 31588 30258 31616 30670
rect 31576 30252 31628 30258
rect 31576 30194 31628 30200
rect 31588 30138 31616 30194
rect 31588 30110 31708 30138
rect 31576 30048 31628 30054
rect 31576 29990 31628 29996
rect 31588 29102 31616 29990
rect 31576 29096 31628 29102
rect 31576 29038 31628 29044
rect 31588 28558 31616 29038
rect 31680 28694 31708 30110
rect 31772 29510 31800 31311
rect 31852 30660 31904 30666
rect 31852 30602 31904 30608
rect 31864 30122 31892 30602
rect 31956 30410 31984 31726
rect 32036 31748 32088 31754
rect 32140 31726 32352 31754
rect 32036 31690 32088 31696
rect 32048 31482 32076 31690
rect 32128 31680 32180 31686
rect 32128 31622 32180 31628
rect 32036 31476 32088 31482
rect 32036 31418 32088 31424
rect 32140 31414 32168 31622
rect 32128 31408 32180 31414
rect 32128 31350 32180 31356
rect 32140 30734 32168 31350
rect 32128 30728 32180 30734
rect 32128 30670 32180 30676
rect 31956 30382 32076 30410
rect 31852 30116 31904 30122
rect 31852 30058 31904 30064
rect 31760 29504 31812 29510
rect 31760 29446 31812 29452
rect 31760 29164 31812 29170
rect 31760 29106 31812 29112
rect 31668 28688 31720 28694
rect 31668 28630 31720 28636
rect 31576 28552 31628 28558
rect 31576 28494 31628 28500
rect 31668 27124 31720 27130
rect 31668 27066 31720 27072
rect 31680 24886 31708 27066
rect 31772 27033 31800 29106
rect 32048 27962 32076 30382
rect 32220 30184 32272 30190
rect 32220 30126 32272 30132
rect 32232 29714 32260 30126
rect 32220 29708 32272 29714
rect 32220 29650 32272 29656
rect 32220 28484 32272 28490
rect 32220 28426 32272 28432
rect 31864 27934 32076 27962
rect 31758 27024 31814 27033
rect 31758 26959 31814 26968
rect 31760 25832 31812 25838
rect 31760 25774 31812 25780
rect 31772 25294 31800 25774
rect 31760 25288 31812 25294
rect 31760 25230 31812 25236
rect 31668 24880 31720 24886
rect 31668 24822 31720 24828
rect 31758 24848 31814 24857
rect 31758 24783 31814 24792
rect 31668 24268 31720 24274
rect 31668 24210 31720 24216
rect 31576 22636 31628 22642
rect 31576 22578 31628 22584
rect 31484 22500 31536 22506
rect 31484 22442 31536 22448
rect 31392 21888 31444 21894
rect 31312 21814 31345 21842
rect 31392 21830 31444 21836
rect 31317 21706 31345 21814
rect 31317 21678 31432 21706
rect 31208 21548 31260 21554
rect 31208 21490 31260 21496
rect 31300 21412 31352 21418
rect 31300 21354 31352 21360
rect 31128 20998 31248 21026
rect 31116 19848 31168 19854
rect 31116 19790 31168 19796
rect 31024 19712 31076 19718
rect 31024 19654 31076 19660
rect 30840 18760 30892 18766
rect 30840 18702 30892 18708
rect 30748 18624 30800 18630
rect 30748 18566 30800 18572
rect 30656 18352 30708 18358
rect 30656 18294 30708 18300
rect 30564 18284 30616 18290
rect 30564 18226 30616 18232
rect 30288 17876 30340 17882
rect 30288 17818 30340 17824
rect 30576 17746 30604 18226
rect 30656 18216 30708 18222
rect 30760 18204 30788 18566
rect 30708 18176 30788 18204
rect 30656 18158 30708 18164
rect 30564 17740 30616 17746
rect 30564 17682 30616 17688
rect 30380 17672 30432 17678
rect 30668 17626 30696 18158
rect 30380 17614 30432 17620
rect 30392 17338 30420 17614
rect 30576 17598 30696 17626
rect 30380 17332 30432 17338
rect 30380 17274 30432 17280
rect 30012 17196 30064 17202
rect 30012 17138 30064 17144
rect 30024 15910 30052 17138
rect 30576 16182 30604 17598
rect 30656 17264 30708 17270
rect 30656 17206 30708 17212
rect 30668 16454 30696 17206
rect 30852 17202 30880 18702
rect 31128 18306 31156 19790
rect 31036 18278 31156 18306
rect 31036 17762 31064 18278
rect 31116 18216 31168 18222
rect 31116 18158 31168 18164
rect 31128 17882 31156 18158
rect 31116 17876 31168 17882
rect 31116 17818 31168 17824
rect 31036 17734 31156 17762
rect 30932 17672 30984 17678
rect 30932 17614 30984 17620
rect 30840 17196 30892 17202
rect 30840 17138 30892 17144
rect 30944 16522 30972 17614
rect 31024 17604 31076 17610
rect 31024 17546 31076 17552
rect 31036 17066 31064 17546
rect 31024 17060 31076 17066
rect 31024 17002 31076 17008
rect 30932 16516 30984 16522
rect 30932 16458 30984 16464
rect 30656 16448 30708 16454
rect 30656 16390 30708 16396
rect 30840 16448 30892 16454
rect 30840 16390 30892 16396
rect 30564 16176 30616 16182
rect 30564 16118 30616 16124
rect 30472 16108 30524 16114
rect 30472 16050 30524 16056
rect 30484 15978 30512 16050
rect 30472 15972 30524 15978
rect 30472 15914 30524 15920
rect 30012 15904 30064 15910
rect 30012 15846 30064 15852
rect 30852 15570 30880 16390
rect 31128 15706 31156 17734
rect 31220 16114 31248 20998
rect 31312 20942 31340 21354
rect 31404 21146 31432 21678
rect 31484 21548 31536 21554
rect 31588 21536 31616 22578
rect 31536 21508 31616 21536
rect 31484 21490 31536 21496
rect 31392 21140 31444 21146
rect 31392 21082 31444 21088
rect 31300 20936 31352 20942
rect 31300 20878 31352 20884
rect 31312 20330 31340 20878
rect 31300 20324 31352 20330
rect 31300 20266 31352 20272
rect 31300 18896 31352 18902
rect 31300 18838 31352 18844
rect 31312 17610 31340 18838
rect 31404 18766 31432 21082
rect 31576 20936 31628 20942
rect 31680 20924 31708 24210
rect 31772 22166 31800 24783
rect 31864 23050 31892 27934
rect 31944 27872 31996 27878
rect 31944 27814 31996 27820
rect 31956 24206 31984 27814
rect 32232 27402 32260 28426
rect 32036 27396 32088 27402
rect 32036 27338 32088 27344
rect 32220 27396 32272 27402
rect 32220 27338 32272 27344
rect 32048 27062 32076 27338
rect 32036 27056 32088 27062
rect 32036 26998 32088 27004
rect 32048 24682 32076 26998
rect 32126 26888 32182 26897
rect 32126 26823 32128 26832
rect 32180 26823 32182 26832
rect 32128 26794 32180 26800
rect 32140 26382 32168 26794
rect 32128 26376 32180 26382
rect 32128 26318 32180 26324
rect 32128 26036 32180 26042
rect 32128 25978 32180 25984
rect 32036 24676 32088 24682
rect 32036 24618 32088 24624
rect 32140 24206 32168 25978
rect 32232 24954 32260 27338
rect 32220 24948 32272 24954
rect 32220 24890 32272 24896
rect 31944 24200 31996 24206
rect 31944 24142 31996 24148
rect 32128 24200 32180 24206
rect 32128 24142 32180 24148
rect 31944 24064 31996 24070
rect 31944 24006 31996 24012
rect 31956 23866 31984 24006
rect 31944 23860 31996 23866
rect 31944 23802 31996 23808
rect 32128 23792 32180 23798
rect 32128 23734 32180 23740
rect 31944 23248 31996 23254
rect 31944 23190 31996 23196
rect 31852 23044 31904 23050
rect 31852 22986 31904 22992
rect 31760 22160 31812 22166
rect 31760 22102 31812 22108
rect 31760 21888 31812 21894
rect 31760 21830 31812 21836
rect 31772 21010 31800 21830
rect 31956 21146 31984 23190
rect 32140 21962 32168 23734
rect 32128 21956 32180 21962
rect 32128 21898 32180 21904
rect 32220 21888 32272 21894
rect 32220 21830 32272 21836
rect 31944 21140 31996 21146
rect 31944 21082 31996 21088
rect 31760 21004 31812 21010
rect 31760 20946 31812 20952
rect 31628 20896 31708 20924
rect 31576 20878 31628 20884
rect 31484 20392 31536 20398
rect 31484 20334 31536 20340
rect 31496 19854 31524 20334
rect 31484 19848 31536 19854
rect 31484 19790 31536 19796
rect 31588 19258 31616 20878
rect 32232 20534 32260 21830
rect 32220 20528 32272 20534
rect 32220 20470 32272 20476
rect 31944 20324 31996 20330
rect 31944 20266 31996 20272
rect 31588 19242 31800 19258
rect 31588 19236 31812 19242
rect 31588 19230 31760 19236
rect 31588 18766 31616 19230
rect 31760 19178 31812 19184
rect 31956 18766 31984 20266
rect 32036 19984 32088 19990
rect 32036 19926 32088 19932
rect 31392 18760 31444 18766
rect 31392 18702 31444 18708
rect 31576 18760 31628 18766
rect 31576 18702 31628 18708
rect 31944 18760 31996 18766
rect 31944 18702 31996 18708
rect 31300 17604 31352 17610
rect 31300 17546 31352 17552
rect 31312 17270 31340 17546
rect 31300 17264 31352 17270
rect 31300 17206 31352 17212
rect 31588 16658 31616 18702
rect 31956 17954 31984 18702
rect 31864 17926 31984 17954
rect 31864 16674 31892 17926
rect 31944 17604 31996 17610
rect 31944 17546 31996 17552
rect 31956 17134 31984 17546
rect 31944 17128 31996 17134
rect 31944 17070 31996 17076
rect 31576 16652 31628 16658
rect 31864 16646 31984 16674
rect 31576 16594 31628 16600
rect 31300 16584 31352 16590
rect 31300 16526 31352 16532
rect 31392 16584 31444 16590
rect 31852 16584 31904 16590
rect 31392 16526 31444 16532
rect 31850 16552 31852 16561
rect 31904 16552 31906 16561
rect 31208 16108 31260 16114
rect 31208 16050 31260 16056
rect 31116 15700 31168 15706
rect 31116 15642 31168 15648
rect 30840 15564 30892 15570
rect 30840 15506 30892 15512
rect 31128 15450 31156 15642
rect 31036 15422 31156 15450
rect 30656 14952 30708 14958
rect 30656 14894 30708 14900
rect 29932 14470 30052 14498
rect 29920 14408 29972 14414
rect 29920 14350 29972 14356
rect 29932 14074 29960 14350
rect 29920 14068 29972 14074
rect 29920 14010 29972 14016
rect 30024 13190 30052 14470
rect 30380 13864 30432 13870
rect 30380 13806 30432 13812
rect 30196 13524 30248 13530
rect 30196 13466 30248 13472
rect 30012 13184 30064 13190
rect 30012 13126 30064 13132
rect 29736 12980 29788 12986
rect 29736 12922 29788 12928
rect 30104 11756 30156 11762
rect 30104 11698 30156 11704
rect 30116 11082 30144 11698
rect 30104 11076 30156 11082
rect 30104 11018 30156 11024
rect 30116 10810 30144 11018
rect 30104 10804 30156 10810
rect 30104 10746 30156 10752
rect 30208 9654 30236 13466
rect 30392 12238 30420 13806
rect 30380 12232 30432 12238
rect 30380 12174 30432 12180
rect 30392 11762 30420 12174
rect 30380 11756 30432 11762
rect 30380 11698 30432 11704
rect 30472 11756 30524 11762
rect 30472 11698 30524 11704
rect 30288 11144 30340 11150
rect 30288 11086 30340 11092
rect 30196 9648 30248 9654
rect 30196 9590 30248 9596
rect 29644 9580 29696 9586
rect 29644 9522 29696 9528
rect 29828 9580 29880 9586
rect 29828 9522 29880 9528
rect 29552 9172 29604 9178
rect 29552 9114 29604 9120
rect 29656 9110 29684 9522
rect 29644 9104 29696 9110
rect 29644 9046 29696 9052
rect 29656 8650 29684 9046
rect 29656 8622 29776 8650
rect 29644 8492 29696 8498
rect 29644 8434 29696 8440
rect 29552 8356 29604 8362
rect 29552 8298 29604 8304
rect 29564 7206 29592 8298
rect 29656 7410 29684 8434
rect 29644 7404 29696 7410
rect 29644 7346 29696 7352
rect 29552 7200 29604 7206
rect 29552 7142 29604 7148
rect 29564 4078 29592 7142
rect 29748 6866 29776 8622
rect 29840 8090 29868 9522
rect 29920 9444 29972 9450
rect 29920 9386 29972 9392
rect 29828 8084 29880 8090
rect 29828 8026 29880 8032
rect 29736 6860 29788 6866
rect 29736 6802 29788 6808
rect 29932 6254 29960 9386
rect 30208 8974 30236 9590
rect 30300 9586 30328 11086
rect 30288 9580 30340 9586
rect 30288 9522 30340 9528
rect 30196 8968 30248 8974
rect 30196 8910 30248 8916
rect 30208 8498 30236 8910
rect 30484 8906 30512 11698
rect 30472 8900 30524 8906
rect 30472 8842 30524 8848
rect 30196 8492 30248 8498
rect 30196 8434 30248 8440
rect 30104 6792 30156 6798
rect 30104 6734 30156 6740
rect 30116 6458 30144 6734
rect 30104 6452 30156 6458
rect 30104 6394 30156 6400
rect 29736 6248 29788 6254
rect 29736 6190 29788 6196
rect 29920 6248 29972 6254
rect 29920 6190 29972 6196
rect 29748 4826 29776 6190
rect 29736 4820 29788 4826
rect 29736 4762 29788 4768
rect 30288 4616 30340 4622
rect 30288 4558 30340 4564
rect 30012 4548 30064 4554
rect 30012 4490 30064 4496
rect 30024 4282 30052 4490
rect 30012 4276 30064 4282
rect 30012 4218 30064 4224
rect 30300 4078 30328 4558
rect 30484 4214 30512 8842
rect 30668 6866 30696 14894
rect 30930 14512 30986 14521
rect 30930 14447 30986 14456
rect 30840 14272 30892 14278
rect 30840 14214 30892 14220
rect 30852 13394 30880 14214
rect 30944 13462 30972 14447
rect 30932 13456 30984 13462
rect 30932 13398 30984 13404
rect 30840 13388 30892 13394
rect 30840 13330 30892 13336
rect 30944 13326 30972 13398
rect 31036 13326 31064 15422
rect 31116 15360 31168 15366
rect 31116 15302 31168 15308
rect 31128 13938 31156 15302
rect 31220 13938 31248 16050
rect 31312 15978 31340 16526
rect 31404 16250 31432 16526
rect 31668 16516 31720 16522
rect 31850 16487 31906 16496
rect 31668 16458 31720 16464
rect 31482 16416 31538 16425
rect 31482 16351 31538 16360
rect 31392 16244 31444 16250
rect 31392 16186 31444 16192
rect 31496 16182 31524 16351
rect 31484 16176 31536 16182
rect 31484 16118 31536 16124
rect 31300 15972 31352 15978
rect 31300 15914 31352 15920
rect 31496 15094 31524 16118
rect 31576 15564 31628 15570
rect 31576 15506 31628 15512
rect 31588 15162 31616 15506
rect 31680 15366 31708 16458
rect 31956 16182 31984 16646
rect 31944 16176 31996 16182
rect 31944 16118 31996 16124
rect 31668 15360 31720 15366
rect 31668 15302 31720 15308
rect 31576 15156 31628 15162
rect 31576 15098 31628 15104
rect 31484 15088 31536 15094
rect 31484 15030 31536 15036
rect 31680 14074 31708 15302
rect 31668 14068 31720 14074
rect 31668 14010 31720 14016
rect 31116 13932 31168 13938
rect 31116 13874 31168 13880
rect 31208 13932 31260 13938
rect 31208 13874 31260 13880
rect 30932 13320 30984 13326
rect 30932 13262 30984 13268
rect 31024 13320 31076 13326
rect 31024 13262 31076 13268
rect 31668 13252 31720 13258
rect 31668 13194 31720 13200
rect 30840 12300 30892 12306
rect 30840 12242 30892 12248
rect 30852 11354 30880 12242
rect 31116 12096 31168 12102
rect 31116 12038 31168 12044
rect 31484 12096 31536 12102
rect 31484 12038 31536 12044
rect 31128 11830 31156 12038
rect 31116 11824 31168 11830
rect 31116 11766 31168 11772
rect 31496 11694 31524 12038
rect 31484 11688 31536 11694
rect 31484 11630 31536 11636
rect 30840 11348 30892 11354
rect 30840 11290 30892 11296
rect 30852 9654 30880 11290
rect 31392 11144 31444 11150
rect 31392 11086 31444 11092
rect 30840 9648 30892 9654
rect 30840 9590 30892 9596
rect 30748 9512 30800 9518
rect 30748 9454 30800 9460
rect 30760 8566 30788 9454
rect 31208 8968 31260 8974
rect 31208 8910 31260 8916
rect 30932 8900 30984 8906
rect 30932 8842 30984 8848
rect 30748 8560 30800 8566
rect 30748 8502 30800 8508
rect 30656 6860 30708 6866
rect 30656 6802 30708 6808
rect 30564 5636 30616 5642
rect 30564 5578 30616 5584
rect 30576 5370 30604 5578
rect 30564 5364 30616 5370
rect 30564 5306 30616 5312
rect 30760 5166 30788 8502
rect 30944 8498 30972 8842
rect 30932 8492 30984 8498
rect 30932 8434 30984 8440
rect 31220 7886 31248 8910
rect 31404 8838 31432 11086
rect 31484 9172 31536 9178
rect 31484 9114 31536 9120
rect 31496 8838 31524 9114
rect 31392 8832 31444 8838
rect 31392 8774 31444 8780
rect 31484 8832 31536 8838
rect 31484 8774 31536 8780
rect 31404 8634 31432 8774
rect 31392 8628 31444 8634
rect 31392 8570 31444 8576
rect 31404 8430 31432 8570
rect 31392 8424 31444 8430
rect 31392 8366 31444 8372
rect 31680 8022 31708 13194
rect 32048 12986 32076 19926
rect 32324 19446 32352 31726
rect 32508 31142 32536 31758
rect 32600 31754 32628 32302
rect 32588 31748 32640 31754
rect 32588 31690 32640 31696
rect 32496 31136 32548 31142
rect 32496 31078 32548 31084
rect 32508 30870 32536 31078
rect 32496 30864 32548 30870
rect 32496 30806 32548 30812
rect 32588 30728 32640 30734
rect 32588 30670 32640 30676
rect 32404 30048 32456 30054
rect 32404 29990 32456 29996
rect 32416 29646 32444 29990
rect 32600 29782 32628 30670
rect 32784 30190 32812 32302
rect 32876 32026 32904 32370
rect 32864 32020 32916 32026
rect 32864 31962 32916 31968
rect 32968 31822 32996 34546
rect 33048 34128 33100 34134
rect 33048 34070 33100 34076
rect 33060 33522 33088 34070
rect 33704 33590 33732 34682
rect 34256 34610 34284 36178
rect 34520 36100 34572 36106
rect 34520 36042 34572 36048
rect 34532 35834 34560 36042
rect 34520 35828 34572 35834
rect 34520 35770 34572 35776
rect 34808 35193 34836 37726
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 36452 37256 36504 37262
rect 36452 37198 36504 37204
rect 35992 36780 36044 36786
rect 35992 36722 36044 36728
rect 35624 36576 35676 36582
rect 35624 36518 35676 36524
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35636 35766 35664 36518
rect 35624 35760 35676 35766
rect 35624 35702 35676 35708
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34794 35184 34850 35193
rect 34794 35119 34850 35128
rect 34704 35080 34756 35086
rect 34704 35022 34756 35028
rect 34244 34604 34296 34610
rect 34244 34546 34296 34552
rect 34520 33924 34572 33930
rect 34520 33866 34572 33872
rect 34426 33824 34482 33833
rect 34426 33759 34482 33768
rect 33692 33584 33744 33590
rect 33692 33526 33744 33532
rect 34334 33552 34390 33561
rect 33048 33516 33100 33522
rect 34440 33522 34468 33759
rect 34334 33487 34336 33496
rect 33048 33458 33100 33464
rect 34388 33487 34390 33496
rect 34428 33516 34480 33522
rect 34336 33458 34388 33464
rect 34428 33458 34480 33464
rect 34532 32910 34560 33866
rect 34716 33590 34744 35022
rect 35440 34944 35492 34950
rect 35440 34886 35492 34892
rect 35452 34610 35480 34886
rect 35440 34604 35492 34610
rect 35440 34546 35492 34552
rect 35348 34400 35400 34406
rect 35348 34342 35400 34348
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35256 34196 35308 34202
rect 35256 34138 35308 34144
rect 34704 33584 34756 33590
rect 34704 33526 34756 33532
rect 34612 33516 34664 33522
rect 34612 33458 34664 33464
rect 34520 32904 34572 32910
rect 34520 32846 34572 32852
rect 34624 32502 34652 33458
rect 34520 32496 34572 32502
rect 34520 32438 34572 32444
rect 34612 32496 34664 32502
rect 34612 32438 34664 32444
rect 34152 32224 34204 32230
rect 34152 32166 34204 32172
rect 32956 31816 33008 31822
rect 32956 31758 33008 31764
rect 32968 31482 32996 31758
rect 32956 31476 33008 31482
rect 32956 31418 33008 31424
rect 34164 31346 34192 32166
rect 34532 31346 34560 32438
rect 34624 31414 34652 32438
rect 34612 31408 34664 31414
rect 34610 31376 34612 31385
rect 34664 31376 34666 31385
rect 34152 31340 34204 31346
rect 34152 31282 34204 31288
rect 34520 31340 34572 31346
rect 34610 31311 34666 31320
rect 34520 31282 34572 31288
rect 34612 31272 34664 31278
rect 34612 31214 34664 31220
rect 34244 30932 34296 30938
rect 34244 30874 34296 30880
rect 34060 30796 34112 30802
rect 34060 30738 34112 30744
rect 34072 30326 34100 30738
rect 34060 30320 34112 30326
rect 34060 30262 34112 30268
rect 32772 30184 32824 30190
rect 32772 30126 32824 30132
rect 32588 29776 32640 29782
rect 32588 29718 32640 29724
rect 32404 29640 32456 29646
rect 32404 29582 32456 29588
rect 32496 29640 32548 29646
rect 32496 29582 32548 29588
rect 32416 29306 32444 29582
rect 32404 29300 32456 29306
rect 32404 29242 32456 29248
rect 32508 28966 32536 29582
rect 32600 29306 32628 29718
rect 32772 29504 32824 29510
rect 32772 29446 32824 29452
rect 33232 29504 33284 29510
rect 33232 29446 33284 29452
rect 32588 29300 32640 29306
rect 32588 29242 32640 29248
rect 32784 29238 32812 29446
rect 33244 29238 33272 29446
rect 32772 29232 32824 29238
rect 32772 29174 32824 29180
rect 33232 29232 33284 29238
rect 33232 29174 33284 29180
rect 32496 28960 32548 28966
rect 32496 28902 32548 28908
rect 32508 28694 32536 28902
rect 32588 28756 32640 28762
rect 32588 28698 32640 28704
rect 32496 28688 32548 28694
rect 32496 28630 32548 28636
rect 32496 27328 32548 27334
rect 32496 27270 32548 27276
rect 32402 26480 32458 26489
rect 32508 26450 32536 27270
rect 32402 26415 32404 26424
rect 32456 26415 32458 26424
rect 32496 26444 32548 26450
rect 32404 26386 32456 26392
rect 32496 26386 32548 26392
rect 32496 25152 32548 25158
rect 32496 25094 32548 25100
rect 32405 24812 32457 24818
rect 32405 24754 32457 24760
rect 32416 24721 32444 24754
rect 32402 24712 32458 24721
rect 32402 24647 32458 24656
rect 32416 24070 32444 24647
rect 32404 24064 32456 24070
rect 32404 24006 32456 24012
rect 32508 22710 32536 25094
rect 32600 24274 32628 28698
rect 32784 28558 32812 29174
rect 33048 29096 33100 29102
rect 33048 29038 33100 29044
rect 32772 28552 32824 28558
rect 32772 28494 32824 28500
rect 32680 28076 32732 28082
rect 32680 28018 32732 28024
rect 32692 26994 32720 28018
rect 32784 27402 32812 28494
rect 33060 28082 33088 29038
rect 33140 28620 33192 28626
rect 33140 28562 33192 28568
rect 33152 28150 33180 28562
rect 33140 28144 33192 28150
rect 33140 28086 33192 28092
rect 33048 28076 33100 28082
rect 33048 28018 33100 28024
rect 33232 27872 33284 27878
rect 33232 27814 33284 27820
rect 32864 27464 32916 27470
rect 32864 27406 32916 27412
rect 32772 27396 32824 27402
rect 32772 27338 32824 27344
rect 32680 26988 32732 26994
rect 32680 26930 32732 26936
rect 32692 25838 32720 26930
rect 32784 26518 32812 27338
rect 32772 26512 32824 26518
rect 32772 26454 32824 26460
rect 32876 26042 32904 27406
rect 32956 27328 33008 27334
rect 32956 27270 33008 27276
rect 32968 27062 32996 27270
rect 32956 27056 33008 27062
rect 32956 26998 33008 27004
rect 33244 26382 33272 27814
rect 33876 26852 33928 26858
rect 33876 26794 33928 26800
rect 33416 26784 33468 26790
rect 33416 26726 33468 26732
rect 33428 26382 33456 26726
rect 33600 26444 33652 26450
rect 33600 26386 33652 26392
rect 33140 26376 33192 26382
rect 33060 26324 33140 26330
rect 33060 26318 33192 26324
rect 33232 26376 33284 26382
rect 33232 26318 33284 26324
rect 33416 26376 33468 26382
rect 33416 26318 33468 26324
rect 33060 26302 33180 26318
rect 32864 26036 32916 26042
rect 32864 25978 32916 25984
rect 32680 25832 32732 25838
rect 32680 25774 32732 25780
rect 32772 25288 32824 25294
rect 32772 25230 32824 25236
rect 32956 25288 33008 25294
rect 32956 25230 33008 25236
rect 32678 24848 32734 24857
rect 32678 24783 32734 24792
rect 32680 24676 32732 24682
rect 32680 24618 32732 24624
rect 32588 24268 32640 24274
rect 32588 24210 32640 24216
rect 32692 24206 32720 24618
rect 32680 24200 32732 24206
rect 32680 24142 32732 24148
rect 32588 24064 32640 24070
rect 32588 24006 32640 24012
rect 32600 23730 32628 24006
rect 32588 23724 32640 23730
rect 32588 23666 32640 23672
rect 32496 22704 32548 22710
rect 32548 22664 32628 22692
rect 32496 22646 32548 22652
rect 32496 22024 32548 22030
rect 32496 21966 32548 21972
rect 32508 21622 32536 21966
rect 32496 21616 32548 21622
rect 32496 21558 32548 21564
rect 32508 20466 32536 21558
rect 32600 21554 32628 22664
rect 32692 22166 32720 24142
rect 32784 23798 32812 25230
rect 32968 24954 32996 25230
rect 32956 24948 33008 24954
rect 32956 24890 33008 24896
rect 33060 23866 33088 26302
rect 33152 26228 33180 26302
rect 33612 26228 33640 26386
rect 33152 26200 33640 26228
rect 33140 25900 33192 25906
rect 33140 25842 33192 25848
rect 33152 25430 33180 25842
rect 33140 25424 33192 25430
rect 33140 25366 33192 25372
rect 33888 25362 33916 26794
rect 33968 26376 34020 26382
rect 33968 26318 34020 26324
rect 34152 26376 34204 26382
rect 34152 26318 34204 26324
rect 33980 25838 34008 26318
rect 34164 25906 34192 26318
rect 34152 25900 34204 25906
rect 34152 25842 34204 25848
rect 33968 25832 34020 25838
rect 33968 25774 34020 25780
rect 33876 25356 33928 25362
rect 33876 25298 33928 25304
rect 33692 25288 33744 25294
rect 33692 25230 33744 25236
rect 33232 24880 33284 24886
rect 33232 24822 33284 24828
rect 33140 24200 33192 24206
rect 33140 24142 33192 24148
rect 33152 23866 33180 24142
rect 33244 24138 33272 24822
rect 33704 24818 33732 25230
rect 33980 24954 34008 25774
rect 34060 25356 34112 25362
rect 34060 25298 34112 25304
rect 33968 24948 34020 24954
rect 33968 24890 34020 24896
rect 34072 24886 34100 25298
rect 34060 24880 34112 24886
rect 34060 24822 34112 24828
rect 33692 24812 33744 24818
rect 33692 24754 33744 24760
rect 33232 24132 33284 24138
rect 33232 24074 33284 24080
rect 33324 24132 33376 24138
rect 33324 24074 33376 24080
rect 33048 23860 33100 23866
rect 33048 23802 33100 23808
rect 33140 23860 33192 23866
rect 33140 23802 33192 23808
rect 32772 23792 32824 23798
rect 32772 23734 32824 23740
rect 33244 23610 33272 24074
rect 32876 23582 33272 23610
rect 32680 22160 32732 22166
rect 32680 22102 32732 22108
rect 32876 21962 32904 23582
rect 32956 23520 33008 23526
rect 32956 23462 33008 23468
rect 32968 23254 32996 23462
rect 33336 23361 33364 24074
rect 33322 23352 33378 23361
rect 33322 23287 33378 23296
rect 32956 23248 33008 23254
rect 32956 23190 33008 23196
rect 33704 22778 33732 24754
rect 34072 24682 34100 24822
rect 34060 24676 34112 24682
rect 34060 24618 34112 24624
rect 33692 22772 33744 22778
rect 33692 22714 33744 22720
rect 33140 22636 33192 22642
rect 33140 22578 33192 22584
rect 33968 22636 34020 22642
rect 33968 22578 34020 22584
rect 33048 22228 33100 22234
rect 33048 22170 33100 22176
rect 33060 22030 33088 22170
rect 33152 22166 33180 22578
rect 33140 22160 33192 22166
rect 33140 22102 33192 22108
rect 33048 22024 33100 22030
rect 33048 21966 33100 21972
rect 32864 21956 32916 21962
rect 32864 21898 32916 21904
rect 32588 21548 32640 21554
rect 32588 21490 32640 21496
rect 32772 20800 32824 20806
rect 32772 20742 32824 20748
rect 32784 20602 32812 20742
rect 32772 20596 32824 20602
rect 32772 20538 32824 20544
rect 32496 20460 32548 20466
rect 32496 20402 32548 20408
rect 32680 20460 32732 20466
rect 32680 20402 32732 20408
rect 32772 20460 32824 20466
rect 32876 20448 32904 21898
rect 32956 21548 33008 21554
rect 32956 21490 33008 21496
rect 32968 20942 32996 21490
rect 32956 20936 33008 20942
rect 32956 20878 33008 20884
rect 32824 20420 32904 20448
rect 32772 20402 32824 20408
rect 32312 19440 32364 19446
rect 32312 19382 32364 19388
rect 32312 18896 32364 18902
rect 32312 18838 32364 18844
rect 32128 17604 32180 17610
rect 32128 17546 32180 17552
rect 32140 14890 32168 17546
rect 32220 16788 32272 16794
rect 32220 16730 32272 16736
rect 32232 16590 32260 16730
rect 32220 16584 32272 16590
rect 32220 16526 32272 16532
rect 32232 16250 32260 16526
rect 32220 16244 32272 16250
rect 32220 16186 32272 16192
rect 32324 15026 32352 18838
rect 32508 18766 32536 20402
rect 32692 19514 32720 20402
rect 32772 20324 32824 20330
rect 32772 20266 32824 20272
rect 32680 19508 32732 19514
rect 32680 19450 32732 19456
rect 32678 19408 32734 19417
rect 32678 19343 32680 19352
rect 32732 19343 32734 19352
rect 32680 19314 32732 19320
rect 32496 18760 32548 18766
rect 32496 18702 32548 18708
rect 32588 17264 32640 17270
rect 32588 17206 32640 17212
rect 32404 17128 32456 17134
rect 32404 17070 32456 17076
rect 32416 16590 32444 17070
rect 32404 16584 32456 16590
rect 32404 16526 32456 16532
rect 32600 16182 32628 17206
rect 32588 16176 32640 16182
rect 32588 16118 32640 16124
rect 32680 16108 32732 16114
rect 32680 16050 32732 16056
rect 32692 15910 32720 16050
rect 32680 15904 32732 15910
rect 32680 15846 32732 15852
rect 32312 15020 32364 15026
rect 32312 14962 32364 14968
rect 32128 14884 32180 14890
rect 32128 14826 32180 14832
rect 32692 14346 32720 15846
rect 32680 14340 32732 14346
rect 32680 14282 32732 14288
rect 32784 14074 32812 20266
rect 32876 18630 32904 20420
rect 32968 19310 32996 20878
rect 33060 20466 33088 21966
rect 33152 21418 33180 22102
rect 33692 22092 33744 22098
rect 33692 22034 33744 22040
rect 33232 21888 33284 21894
rect 33232 21830 33284 21836
rect 33244 21622 33272 21830
rect 33704 21622 33732 22034
rect 33980 22030 34008 22578
rect 33968 22024 34020 22030
rect 33968 21966 34020 21972
rect 33232 21616 33284 21622
rect 33232 21558 33284 21564
rect 33692 21616 33744 21622
rect 33692 21558 33744 21564
rect 33140 21412 33192 21418
rect 33140 21354 33192 21360
rect 33600 21072 33652 21078
rect 33600 21014 33652 21020
rect 33140 20868 33192 20874
rect 33140 20810 33192 20816
rect 33152 20602 33180 20810
rect 33140 20596 33192 20602
rect 33140 20538 33192 20544
rect 33612 20534 33640 21014
rect 33980 20602 34008 21966
rect 33968 20596 34020 20602
rect 33968 20538 34020 20544
rect 33232 20528 33284 20534
rect 33232 20470 33284 20476
rect 33600 20528 33652 20534
rect 33600 20470 33652 20476
rect 33048 20460 33100 20466
rect 33048 20402 33100 20408
rect 33140 20460 33192 20466
rect 33140 20402 33192 20408
rect 32956 19304 33008 19310
rect 32956 19246 33008 19252
rect 33060 18902 33088 20402
rect 33152 19854 33180 20402
rect 33140 19848 33192 19854
rect 33140 19790 33192 19796
rect 32956 18896 33008 18902
rect 32956 18838 33008 18844
rect 33048 18896 33100 18902
rect 33048 18838 33100 18844
rect 32968 18630 32996 18838
rect 32864 18624 32916 18630
rect 32864 18566 32916 18572
rect 32956 18624 33008 18630
rect 32956 18566 33008 18572
rect 32876 17134 32904 18566
rect 33060 17746 33088 18838
rect 33152 18426 33180 19790
rect 33244 19786 33272 20470
rect 33612 19990 33640 20470
rect 33600 19984 33652 19990
rect 33600 19926 33652 19932
rect 33232 19780 33284 19786
rect 33232 19722 33284 19728
rect 33508 19440 33560 19446
rect 33322 19408 33378 19417
rect 33508 19382 33560 19388
rect 33322 19343 33324 19352
rect 33376 19343 33378 19352
rect 33324 19314 33376 19320
rect 33324 19168 33376 19174
rect 33324 19110 33376 19116
rect 33232 18896 33284 18902
rect 33232 18838 33284 18844
rect 33336 18850 33364 19110
rect 33520 18970 33548 19382
rect 33508 18964 33560 18970
rect 33508 18906 33560 18912
rect 33244 18766 33272 18838
rect 33336 18822 33456 18850
rect 33232 18760 33284 18766
rect 33232 18702 33284 18708
rect 33322 18728 33378 18737
rect 33322 18663 33324 18672
rect 33376 18663 33378 18672
rect 33324 18634 33376 18640
rect 33140 18420 33192 18426
rect 33140 18362 33192 18368
rect 33428 18290 33456 18822
rect 33600 18692 33652 18698
rect 33600 18634 33652 18640
rect 33784 18692 33836 18698
rect 33784 18634 33836 18640
rect 33416 18284 33468 18290
rect 33416 18226 33468 18232
rect 33048 17740 33100 17746
rect 33048 17682 33100 17688
rect 33140 17672 33192 17678
rect 33140 17614 33192 17620
rect 33324 17672 33376 17678
rect 33324 17614 33376 17620
rect 33152 17218 33180 17614
rect 33232 17536 33284 17542
rect 33232 17478 33284 17484
rect 33060 17190 33180 17218
rect 33244 17202 33272 17478
rect 33232 17196 33284 17202
rect 32864 17128 32916 17134
rect 32864 17070 32916 17076
rect 32876 16522 32904 17070
rect 32956 16992 33008 16998
rect 32956 16934 33008 16940
rect 33060 16946 33088 17190
rect 33232 17138 33284 17144
rect 33336 17066 33364 17614
rect 33324 17060 33376 17066
rect 33324 17002 33376 17008
rect 32864 16516 32916 16522
rect 32864 16458 32916 16464
rect 32968 16182 32996 16934
rect 33060 16918 33180 16946
rect 33152 16794 33180 16918
rect 33140 16788 33192 16794
rect 33140 16730 33192 16736
rect 32956 16176 33008 16182
rect 32956 16118 33008 16124
rect 33152 15638 33180 16730
rect 33140 15632 33192 15638
rect 33140 15574 33192 15580
rect 33336 14482 33364 17002
rect 33428 16658 33456 18226
rect 33612 18222 33640 18634
rect 33692 18284 33744 18290
rect 33692 18226 33744 18232
rect 33600 18216 33652 18222
rect 33600 18158 33652 18164
rect 33508 18080 33560 18086
rect 33508 18022 33560 18028
rect 33520 17882 33548 18022
rect 33508 17876 33560 17882
rect 33508 17818 33560 17824
rect 33416 16652 33468 16658
rect 33416 16594 33468 16600
rect 33520 15638 33548 17818
rect 33704 17542 33732 18226
rect 33692 17536 33744 17542
rect 33692 17478 33744 17484
rect 33704 16590 33732 17478
rect 33692 16584 33744 16590
rect 33692 16526 33744 16532
rect 33508 15632 33560 15638
rect 33508 15574 33560 15580
rect 33520 15502 33548 15574
rect 33508 15496 33560 15502
rect 33508 15438 33560 15444
rect 33416 15360 33468 15366
rect 33416 15302 33468 15308
rect 33508 15360 33560 15366
rect 33508 15302 33560 15308
rect 33428 15094 33456 15302
rect 33416 15088 33468 15094
rect 33416 15030 33468 15036
rect 33324 14476 33376 14482
rect 33324 14418 33376 14424
rect 33428 14414 33456 15030
rect 33520 15026 33548 15302
rect 33508 15020 33560 15026
rect 33508 14962 33560 14968
rect 33416 14408 33468 14414
rect 33046 14376 33102 14385
rect 33416 14350 33468 14356
rect 33046 14311 33102 14320
rect 33508 14340 33560 14346
rect 32772 14068 32824 14074
rect 32772 14010 32824 14016
rect 33060 13938 33088 14311
rect 33508 14282 33560 14288
rect 33520 14006 33548 14282
rect 33508 14000 33560 14006
rect 33508 13942 33560 13948
rect 33048 13932 33100 13938
rect 33048 13874 33100 13880
rect 32864 13864 32916 13870
rect 32864 13806 32916 13812
rect 33324 13864 33376 13870
rect 33324 13806 33376 13812
rect 32036 12980 32088 12986
rect 32036 12922 32088 12928
rect 32048 12170 32076 12922
rect 32876 12782 32904 13806
rect 32864 12776 32916 12782
rect 32864 12718 32916 12724
rect 33048 12776 33100 12782
rect 33048 12718 33100 12724
rect 32588 12640 32640 12646
rect 32588 12582 32640 12588
rect 32600 12238 32628 12582
rect 32496 12232 32548 12238
rect 32496 12174 32548 12180
rect 32588 12232 32640 12238
rect 32588 12174 32640 12180
rect 32036 12164 32088 12170
rect 32036 12106 32088 12112
rect 31852 11552 31904 11558
rect 31852 11494 31904 11500
rect 31760 9376 31812 9382
rect 31760 9318 31812 9324
rect 31772 8974 31800 9318
rect 31760 8968 31812 8974
rect 31760 8910 31812 8916
rect 31864 8430 31892 11494
rect 31944 9988 31996 9994
rect 31944 9930 31996 9936
rect 31852 8424 31904 8430
rect 31852 8366 31904 8372
rect 31668 8016 31720 8022
rect 31668 7958 31720 7964
rect 31208 7880 31260 7886
rect 31208 7822 31260 7828
rect 31668 7880 31720 7886
rect 31668 7822 31720 7828
rect 31680 7410 31708 7822
rect 31668 7404 31720 7410
rect 31668 7346 31720 7352
rect 31024 7200 31076 7206
rect 31024 7142 31076 7148
rect 30840 6316 30892 6322
rect 30840 6258 30892 6264
rect 30852 5574 30880 6258
rect 31036 6254 31064 7142
rect 30932 6248 30984 6254
rect 30932 6190 30984 6196
rect 31024 6248 31076 6254
rect 31024 6190 31076 6196
rect 30840 5568 30892 5574
rect 30840 5510 30892 5516
rect 30852 5370 30880 5510
rect 30840 5364 30892 5370
rect 30840 5306 30892 5312
rect 30748 5160 30800 5166
rect 30748 5102 30800 5108
rect 30944 4826 30972 6190
rect 31680 5710 31708 7346
rect 31956 7206 31984 9930
rect 32048 9586 32076 12106
rect 32312 11756 32364 11762
rect 32312 11698 32364 11704
rect 32324 10266 32352 11698
rect 32508 11218 32536 12174
rect 32876 11762 32904 12718
rect 33060 12238 33088 12718
rect 33232 12436 33284 12442
rect 33336 12434 33364 13806
rect 33796 13462 33824 18634
rect 34256 17202 34284 30874
rect 34624 30802 34652 31214
rect 34612 30796 34664 30802
rect 34612 30738 34664 30744
rect 34612 26852 34664 26858
rect 34612 26794 34664 26800
rect 34624 26761 34652 26794
rect 34610 26752 34666 26761
rect 34610 26687 34666 26696
rect 34612 25152 34664 25158
rect 34612 25094 34664 25100
rect 34624 24818 34652 25094
rect 34336 24812 34388 24818
rect 34336 24754 34388 24760
rect 34520 24812 34572 24818
rect 34520 24754 34572 24760
rect 34612 24812 34664 24818
rect 34612 24754 34664 24760
rect 34348 24410 34376 24754
rect 34532 24682 34560 24754
rect 34520 24676 34572 24682
rect 34520 24618 34572 24624
rect 34336 24404 34388 24410
rect 34336 24346 34388 24352
rect 34716 24290 34744 33526
rect 34888 33516 34940 33522
rect 34808 33476 34888 33504
rect 34808 32570 34836 33476
rect 34888 33458 34940 33464
rect 35268 33454 35296 34138
rect 35256 33448 35308 33454
rect 35256 33390 35308 33396
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35164 32904 35216 32910
rect 35164 32846 35216 32852
rect 34888 32768 34940 32774
rect 34888 32710 34940 32716
rect 34796 32564 34848 32570
rect 34796 32506 34848 32512
rect 34808 31464 34836 32506
rect 34900 32434 34928 32710
rect 35176 32502 35204 32846
rect 35256 32564 35308 32570
rect 35256 32506 35308 32512
rect 35164 32496 35216 32502
rect 35164 32438 35216 32444
rect 35268 32434 35296 32506
rect 35360 32450 35388 34342
rect 35452 34202 35480 34546
rect 35440 34196 35492 34202
rect 35440 34138 35492 34144
rect 35532 33856 35584 33862
rect 35532 33798 35584 33804
rect 35440 32904 35492 32910
rect 35440 32846 35492 32852
rect 35452 32570 35480 32846
rect 35440 32564 35492 32570
rect 35440 32506 35492 32512
rect 34888 32428 34940 32434
rect 34888 32370 34940 32376
rect 35256 32428 35308 32434
rect 35360 32422 35480 32450
rect 35256 32370 35308 32376
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35452 31822 35480 32422
rect 35256 31816 35308 31822
rect 35256 31758 35308 31764
rect 35440 31816 35492 31822
rect 35440 31758 35492 31764
rect 35268 31482 35296 31758
rect 35256 31476 35308 31482
rect 34808 31436 34928 31464
rect 34794 31376 34850 31385
rect 34900 31346 34928 31436
rect 35256 31418 35308 31424
rect 35348 31476 35400 31482
rect 35348 31418 35400 31424
rect 34794 31311 34850 31320
rect 34888 31340 34940 31346
rect 34808 30666 34836 31311
rect 34888 31282 34940 31288
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34796 30660 34848 30666
rect 34796 30602 34848 30608
rect 34808 29646 34836 30602
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34886 29744 34942 29753
rect 34886 29679 34942 29688
rect 34796 29640 34848 29646
rect 34796 29582 34848 29588
rect 34900 29050 34928 29679
rect 34808 29022 34928 29050
rect 34808 27538 34836 29022
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35360 28762 35388 31418
rect 35544 31414 35572 33798
rect 35636 33454 35664 35702
rect 36004 35698 36032 36722
rect 36268 36168 36320 36174
rect 36268 36110 36320 36116
rect 36084 36032 36136 36038
rect 36084 35974 36136 35980
rect 35992 35692 36044 35698
rect 35992 35634 36044 35640
rect 35716 33652 35768 33658
rect 35716 33594 35768 33600
rect 35728 33522 35756 33594
rect 35898 33552 35954 33561
rect 35716 33516 35768 33522
rect 35898 33487 35900 33496
rect 35716 33458 35768 33464
rect 35952 33487 35954 33496
rect 35900 33458 35952 33464
rect 35624 33448 35676 33454
rect 35624 33390 35676 33396
rect 35728 33114 35756 33458
rect 35716 33108 35768 33114
rect 35716 33050 35768 33056
rect 35624 32360 35676 32366
rect 35624 32302 35676 32308
rect 35636 31482 35664 32302
rect 35728 32298 35756 33050
rect 35808 32496 35860 32502
rect 35808 32438 35860 32444
rect 35716 32292 35768 32298
rect 35716 32234 35768 32240
rect 35728 31958 35756 32234
rect 35716 31952 35768 31958
rect 35716 31894 35768 31900
rect 35820 31754 35848 32438
rect 35912 31822 35940 33458
rect 35900 31816 35952 31822
rect 35900 31758 35952 31764
rect 35728 31726 35848 31754
rect 35624 31476 35676 31482
rect 35624 31418 35676 31424
rect 35532 31408 35584 31414
rect 35532 31350 35584 31356
rect 35440 31340 35492 31346
rect 35440 31282 35492 31288
rect 35452 30734 35480 31282
rect 35532 30796 35584 30802
rect 35532 30738 35584 30744
rect 35440 30728 35492 30734
rect 35544 30705 35572 30738
rect 35440 30670 35492 30676
rect 35530 30696 35586 30705
rect 35452 29753 35480 30670
rect 35530 30631 35586 30640
rect 35532 30592 35584 30598
rect 35532 30534 35584 30540
rect 35438 29744 35494 29753
rect 35438 29679 35440 29688
rect 35492 29679 35494 29688
rect 35440 29650 35492 29656
rect 35544 29646 35572 30534
rect 35532 29640 35584 29646
rect 35728 29594 35756 31726
rect 35808 30592 35860 30598
rect 35808 30534 35860 30540
rect 35820 30258 35848 30534
rect 35912 30394 35940 31758
rect 36004 31210 36032 35634
rect 36096 34066 36124 35974
rect 36280 35154 36308 36110
rect 36464 35834 36492 37198
rect 36728 37188 36780 37194
rect 36728 37130 36780 37136
rect 36740 36961 36768 37130
rect 36726 36952 36782 36961
rect 36726 36887 36782 36896
rect 36832 36854 36860 38247
rect 38212 37346 38240 39200
rect 38120 37318 38240 37346
rect 38120 37262 38148 37318
rect 38108 37256 38160 37262
rect 38108 37198 38160 37204
rect 38016 37188 38068 37194
rect 38016 37130 38068 37136
rect 38028 36922 38056 37130
rect 38016 36916 38068 36922
rect 38016 36858 38068 36864
rect 36820 36848 36872 36854
rect 36820 36790 36872 36796
rect 37740 36780 37792 36786
rect 37740 36722 37792 36728
rect 37464 36100 37516 36106
rect 37464 36042 37516 36048
rect 37476 35834 37504 36042
rect 36452 35828 36504 35834
rect 36452 35770 36504 35776
rect 37464 35828 37516 35834
rect 37464 35770 37516 35776
rect 37752 35630 37780 36722
rect 38108 36712 38160 36718
rect 38108 36654 38160 36660
rect 37832 36032 37884 36038
rect 37832 35974 37884 35980
rect 37844 35698 37872 35974
rect 37832 35692 37884 35698
rect 37832 35634 37884 35640
rect 37740 35624 37792 35630
rect 37740 35566 37792 35572
rect 36268 35148 36320 35154
rect 36268 35090 36320 35096
rect 36176 35012 36228 35018
rect 36176 34954 36228 34960
rect 36188 34746 36216 34954
rect 36176 34740 36228 34746
rect 36176 34682 36228 34688
rect 36084 34060 36136 34066
rect 36084 34002 36136 34008
rect 36096 32842 36124 34002
rect 36176 33516 36228 33522
rect 36176 33458 36228 33464
rect 36188 32910 36216 33458
rect 36280 33046 36308 35090
rect 36636 34536 36688 34542
rect 36636 34478 36688 34484
rect 36648 33658 36676 34478
rect 37188 33992 37240 33998
rect 37188 33934 37240 33940
rect 36636 33652 36688 33658
rect 36636 33594 36688 33600
rect 37200 33454 37228 33934
rect 36360 33448 36412 33454
rect 36360 33390 36412 33396
rect 37188 33448 37240 33454
rect 37188 33390 37240 33396
rect 36372 33114 36400 33390
rect 37752 33386 37780 35566
rect 37844 34134 37872 35634
rect 38016 35624 38068 35630
rect 38120 35601 38148 36654
rect 38016 35566 38068 35572
rect 38106 35592 38162 35601
rect 38028 34474 38056 35566
rect 38106 35527 38162 35536
rect 38108 34536 38160 34542
rect 38108 34478 38160 34484
rect 38016 34468 38068 34474
rect 38016 34410 38068 34416
rect 37832 34128 37884 34134
rect 37832 34070 37884 34076
rect 37832 33516 37884 33522
rect 37832 33458 37884 33464
rect 37740 33380 37792 33386
rect 37740 33322 37792 33328
rect 37096 33312 37148 33318
rect 37096 33254 37148 33260
rect 36360 33108 36412 33114
rect 36360 33050 36412 33056
rect 36268 33040 36320 33046
rect 36268 32982 36320 32988
rect 36176 32904 36228 32910
rect 36176 32846 36228 32852
rect 36084 32836 36136 32842
rect 36084 32778 36136 32784
rect 36084 32292 36136 32298
rect 36084 32234 36136 32240
rect 35992 31204 36044 31210
rect 35992 31146 36044 31152
rect 35900 30388 35952 30394
rect 35900 30330 35952 30336
rect 35898 30288 35954 30297
rect 35808 30252 35860 30258
rect 36096 30258 36124 32234
rect 36176 32224 36228 32230
rect 36176 32166 36228 32172
rect 36188 30326 36216 32166
rect 36280 31906 36308 32982
rect 37108 32910 37136 33254
rect 37096 32904 37148 32910
rect 37096 32846 37148 32852
rect 37844 32774 37872 33458
rect 38028 33454 38056 34410
rect 38120 34241 38148 34478
rect 38106 34232 38162 34241
rect 38106 34167 38162 34176
rect 38108 33924 38160 33930
rect 38108 33866 38160 33872
rect 38016 33448 38068 33454
rect 38016 33390 38068 33396
rect 37832 32768 37884 32774
rect 37832 32710 37884 32716
rect 37832 32428 37884 32434
rect 37832 32370 37884 32376
rect 37844 32026 37872 32370
rect 37832 32020 37884 32026
rect 37832 31962 37884 31968
rect 36280 31890 36400 31906
rect 36268 31884 36400 31890
rect 36320 31878 36400 31884
rect 36268 31826 36320 31832
rect 36176 30320 36228 30326
rect 36176 30262 36228 30268
rect 36084 30252 36136 30258
rect 35898 30223 35900 30232
rect 35808 30194 35860 30200
rect 35952 30223 35954 30232
rect 35900 30194 35952 30200
rect 36004 30212 36084 30240
rect 35532 29582 35584 29588
rect 35440 29572 35492 29578
rect 35440 29514 35492 29520
rect 35636 29566 35756 29594
rect 35348 28756 35400 28762
rect 35348 28698 35400 28704
rect 35348 28484 35400 28490
rect 35348 28426 35400 28432
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34796 27532 34848 27538
rect 34796 27474 34848 27480
rect 34796 26988 34848 26994
rect 34796 26930 34848 26936
rect 34808 26586 34836 26930
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34796 26580 34848 26586
rect 34796 26522 34848 26528
rect 35360 25974 35388 28426
rect 35452 26382 35480 29514
rect 35532 27600 35584 27606
rect 35532 27542 35584 27548
rect 35544 26382 35572 27542
rect 35440 26376 35492 26382
rect 35440 26318 35492 26324
rect 35532 26376 35584 26382
rect 35532 26318 35584 26324
rect 35348 25968 35400 25974
rect 35348 25910 35400 25916
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35360 24818 35388 25910
rect 35348 24812 35400 24818
rect 35348 24754 35400 24760
rect 35636 24698 35664 29566
rect 35716 29504 35768 29510
rect 35716 29446 35768 29452
rect 35728 29170 35756 29446
rect 36004 29170 36032 30212
rect 36084 30194 36136 30200
rect 36268 30252 36320 30258
rect 36268 30194 36320 30200
rect 36084 30116 36136 30122
rect 36084 30058 36136 30064
rect 36096 29238 36124 30058
rect 36084 29232 36136 29238
rect 36084 29174 36136 29180
rect 36280 29170 36308 30194
rect 36372 29714 36400 31878
rect 37464 31816 37516 31822
rect 37464 31758 37516 31764
rect 37476 31482 37504 31758
rect 37740 31680 37792 31686
rect 37740 31622 37792 31628
rect 37464 31476 37516 31482
rect 37464 31418 37516 31424
rect 37752 31346 37780 31622
rect 37844 31482 37872 31962
rect 37832 31476 37884 31482
rect 37832 31418 37884 31424
rect 37740 31340 37792 31346
rect 37740 31282 37792 31288
rect 38028 31278 38056 33390
rect 38120 32881 38148 33866
rect 38106 32872 38162 32881
rect 38106 32807 38162 32816
rect 38108 32360 38160 32366
rect 38108 32302 38160 32308
rect 38120 31521 38148 32302
rect 38106 31512 38162 31521
rect 38106 31447 38162 31456
rect 38016 31272 38068 31278
rect 38016 31214 38068 31220
rect 36728 30728 36780 30734
rect 36728 30670 36780 30676
rect 36740 30326 36768 30670
rect 37004 30660 37056 30666
rect 37004 30602 37056 30608
rect 37280 30660 37332 30666
rect 37280 30602 37332 30608
rect 36728 30320 36780 30326
rect 36728 30262 36780 30268
rect 37016 30161 37044 30602
rect 37002 30152 37058 30161
rect 37002 30087 37058 30096
rect 36360 29708 36412 29714
rect 36360 29650 36412 29656
rect 36820 29708 36872 29714
rect 36820 29650 36872 29656
rect 35716 29164 35768 29170
rect 35716 29106 35768 29112
rect 35808 29164 35860 29170
rect 35808 29106 35860 29112
rect 35992 29164 36044 29170
rect 35992 29106 36044 29112
rect 36268 29164 36320 29170
rect 36268 29106 36320 29112
rect 35716 28756 35768 28762
rect 35716 28698 35768 28704
rect 35360 24670 35664 24698
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35256 24336 35308 24342
rect 34716 24262 34928 24290
rect 35256 24278 35308 24284
rect 34428 23792 34480 23798
rect 34428 23734 34480 23740
rect 34440 21486 34468 23734
rect 34900 23730 34928 24262
rect 35268 23730 35296 24278
rect 34796 23724 34848 23730
rect 34796 23666 34848 23672
rect 34888 23724 34940 23730
rect 34888 23666 34940 23672
rect 35256 23724 35308 23730
rect 35256 23666 35308 23672
rect 34520 23112 34572 23118
rect 34518 23080 34520 23089
rect 34572 23080 34574 23089
rect 34518 23015 34574 23024
rect 34612 22568 34664 22574
rect 34612 22510 34664 22516
rect 34428 21480 34480 21486
rect 34428 21422 34480 21428
rect 34520 21480 34572 21486
rect 34520 21422 34572 21428
rect 34440 21350 34468 21422
rect 34428 21344 34480 21350
rect 34428 21286 34480 21292
rect 34440 19446 34468 21286
rect 34532 20262 34560 21422
rect 34624 21010 34652 22510
rect 34808 21554 34836 23666
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34796 21548 34848 21554
rect 34796 21490 34848 21496
rect 35256 21548 35308 21554
rect 35256 21490 35308 21496
rect 34612 21004 34664 21010
rect 34612 20946 34664 20952
rect 34520 20256 34572 20262
rect 34520 20198 34572 20204
rect 34428 19440 34480 19446
rect 34428 19382 34480 19388
rect 34428 18352 34480 18358
rect 34428 18294 34480 18300
rect 34244 17196 34296 17202
rect 34244 17138 34296 17144
rect 33968 14816 34020 14822
rect 33968 14758 34020 14764
rect 33980 13938 34008 14758
rect 33968 13932 34020 13938
rect 33968 13874 34020 13880
rect 33784 13456 33836 13462
rect 33784 13398 33836 13404
rect 33876 12844 33928 12850
rect 33876 12786 33928 12792
rect 33888 12442 33916 12786
rect 33284 12406 33364 12434
rect 33876 12436 33928 12442
rect 33232 12378 33284 12384
rect 34440 12434 34468 18294
rect 34520 15700 34572 15706
rect 34520 15642 34572 15648
rect 34532 14482 34560 15642
rect 34520 14476 34572 14482
rect 34520 14418 34572 14424
rect 34520 13184 34572 13190
rect 34520 13126 34572 13132
rect 33876 12378 33928 12384
rect 34348 12406 34468 12434
rect 33048 12232 33100 12238
rect 33048 12174 33100 12180
rect 33060 11830 33088 12174
rect 33048 11824 33100 11830
rect 33048 11766 33100 11772
rect 33888 11762 33916 12378
rect 34348 12170 34376 12406
rect 34428 12300 34480 12306
rect 34428 12242 34480 12248
rect 34336 12164 34388 12170
rect 34336 12106 34388 12112
rect 32864 11756 32916 11762
rect 32864 11698 32916 11704
rect 33140 11756 33192 11762
rect 33140 11698 33192 11704
rect 33876 11756 33928 11762
rect 33876 11698 33928 11704
rect 33152 11286 33180 11698
rect 34440 11354 34468 12242
rect 34428 11348 34480 11354
rect 34428 11290 34480 11296
rect 33140 11280 33192 11286
rect 33140 11222 33192 11228
rect 33600 11280 33652 11286
rect 33600 11222 33652 11228
rect 32496 11212 32548 11218
rect 32496 11154 32548 11160
rect 32956 11212 33008 11218
rect 32956 11154 33008 11160
rect 32312 10260 32364 10266
rect 32312 10202 32364 10208
rect 32968 10130 32996 11154
rect 33232 11076 33284 11082
rect 33232 11018 33284 11024
rect 32956 10124 33008 10130
rect 32956 10066 33008 10072
rect 32128 10056 32180 10062
rect 32128 9998 32180 10004
rect 32140 9654 32168 9998
rect 32772 9920 32824 9926
rect 32772 9862 32824 9868
rect 32784 9654 32812 9862
rect 33244 9722 33272 11018
rect 33324 10600 33376 10606
rect 33324 10542 33376 10548
rect 33232 9716 33284 9722
rect 33232 9658 33284 9664
rect 32128 9648 32180 9654
rect 32128 9590 32180 9596
rect 32588 9648 32640 9654
rect 32772 9648 32824 9654
rect 32588 9590 32640 9596
rect 32692 9596 32772 9602
rect 32692 9590 32824 9596
rect 32036 9580 32088 9586
rect 32036 9522 32088 9528
rect 32600 9178 32628 9590
rect 32692 9574 32812 9590
rect 32588 9172 32640 9178
rect 32588 9114 32640 9120
rect 32692 8498 32720 9574
rect 32772 9512 32824 9518
rect 32772 9454 32824 9460
rect 32784 8634 32812 9454
rect 32864 8968 32916 8974
rect 32864 8910 32916 8916
rect 32772 8628 32824 8634
rect 32772 8570 32824 8576
rect 32876 8498 32904 8910
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 32864 8492 32916 8498
rect 32864 8434 32916 8440
rect 32496 8288 32548 8294
rect 32496 8230 32548 8236
rect 32508 7818 32536 8230
rect 32876 8090 32904 8434
rect 32864 8084 32916 8090
rect 32864 8026 32916 8032
rect 33244 7886 33272 9658
rect 33232 7880 33284 7886
rect 33232 7822 33284 7828
rect 32496 7812 32548 7818
rect 32496 7754 32548 7760
rect 32956 7404 33008 7410
rect 32956 7346 33008 7352
rect 31944 7200 31996 7206
rect 31944 7142 31996 7148
rect 32968 7002 32996 7346
rect 32956 6996 33008 7002
rect 32956 6938 33008 6944
rect 33048 6860 33100 6866
rect 33048 6802 33100 6808
rect 33060 5778 33088 6802
rect 33336 6662 33364 10542
rect 33508 10464 33560 10470
rect 33508 10406 33560 10412
rect 33520 10062 33548 10406
rect 33508 10056 33560 10062
rect 33508 9998 33560 10004
rect 33612 9994 33640 11222
rect 34244 10668 34296 10674
rect 34244 10610 34296 10616
rect 34256 10198 34284 10610
rect 34440 10606 34468 11290
rect 34428 10600 34480 10606
rect 34428 10542 34480 10548
rect 34244 10192 34296 10198
rect 34244 10134 34296 10140
rect 33416 9988 33468 9994
rect 33416 9930 33468 9936
rect 33600 9988 33652 9994
rect 33600 9930 33652 9936
rect 33428 9178 33456 9930
rect 33612 9722 33640 9930
rect 33600 9716 33652 9722
rect 33600 9658 33652 9664
rect 34152 9580 34204 9586
rect 34152 9522 34204 9528
rect 34164 9382 34192 9522
rect 34152 9376 34204 9382
rect 34152 9318 34204 9324
rect 33416 9172 33468 9178
rect 33416 9114 33468 9120
rect 33876 8900 33928 8906
rect 33876 8842 33928 8848
rect 33888 8566 33916 8842
rect 33876 8560 33928 8566
rect 33876 8502 33928 8508
rect 33324 6656 33376 6662
rect 33324 6598 33376 6604
rect 33888 6390 33916 8502
rect 33968 8492 34020 8498
rect 33968 8434 34020 8440
rect 33980 7546 34008 8434
rect 33968 7540 34020 7546
rect 33968 7482 34020 7488
rect 33980 6798 34008 7482
rect 34164 6934 34192 9318
rect 34440 8022 34468 10542
rect 34532 10198 34560 13126
rect 34624 11898 34652 20946
rect 34808 19334 34836 21490
rect 35268 21350 35296 21490
rect 35360 21418 35388 24670
rect 35624 23588 35676 23594
rect 35624 23530 35676 23536
rect 35530 23216 35586 23225
rect 35530 23151 35586 23160
rect 35544 23118 35572 23151
rect 35532 23112 35584 23118
rect 35532 23054 35584 23060
rect 35440 22976 35492 22982
rect 35440 22918 35492 22924
rect 35452 22642 35480 22918
rect 35440 22636 35492 22642
rect 35440 22578 35492 22584
rect 35532 22636 35584 22642
rect 35532 22578 35584 22584
rect 35544 22234 35572 22578
rect 35532 22228 35584 22234
rect 35532 22170 35584 22176
rect 35636 22094 35664 23530
rect 35728 22642 35756 28698
rect 35820 28422 35848 29106
rect 35808 28416 35860 28422
rect 35808 28358 35860 28364
rect 35820 28150 35848 28358
rect 35808 28144 35860 28150
rect 35808 28086 35860 28092
rect 35808 27532 35860 27538
rect 35808 27474 35860 27480
rect 35820 26994 35848 27474
rect 36004 27130 36032 29106
rect 36280 28218 36308 29106
rect 36636 29028 36688 29034
rect 36636 28970 36688 28976
rect 36268 28212 36320 28218
rect 36268 28154 36320 28160
rect 36084 28076 36136 28082
rect 36084 28018 36136 28024
rect 35992 27124 36044 27130
rect 35992 27066 36044 27072
rect 35808 26988 35860 26994
rect 35808 26930 35860 26936
rect 35808 26784 35860 26790
rect 35808 26726 35860 26732
rect 35820 26382 35848 26726
rect 35808 26376 35860 26382
rect 35808 26318 35860 26324
rect 35808 23180 35860 23186
rect 35808 23122 35860 23128
rect 35820 22710 35848 23122
rect 35808 22704 35860 22710
rect 35808 22646 35860 22652
rect 35716 22636 35768 22642
rect 35716 22578 35768 22584
rect 35452 22066 35664 22094
rect 35348 21412 35400 21418
rect 35348 21354 35400 21360
rect 35256 21344 35308 21350
rect 35256 21286 35308 21292
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34980 19712 35032 19718
rect 35032 19672 35112 19700
rect 34980 19654 35032 19660
rect 35084 19378 35112 19672
rect 35164 19440 35216 19446
rect 35216 19400 35388 19428
rect 35164 19382 35216 19388
rect 34888 19372 34940 19378
rect 34808 19320 34888 19334
rect 34808 19314 34940 19320
rect 35072 19372 35124 19378
rect 35072 19314 35124 19320
rect 34808 19306 34928 19314
rect 34808 18766 34836 19306
rect 35164 19304 35216 19310
rect 34992 19252 35164 19258
rect 34992 19246 35216 19252
rect 34992 19242 35204 19246
rect 34980 19236 35204 19242
rect 35032 19230 35204 19236
rect 34980 19178 35032 19184
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34888 18896 34940 18902
rect 34888 18838 34940 18844
rect 35162 18864 35218 18873
rect 34796 18760 34848 18766
rect 34796 18702 34848 18708
rect 34808 17202 34836 18702
rect 34900 18630 34928 18838
rect 35162 18799 35218 18808
rect 35176 18766 35204 18799
rect 35360 18766 35388 19400
rect 35164 18760 35216 18766
rect 35164 18702 35216 18708
rect 35348 18760 35400 18766
rect 35348 18702 35400 18708
rect 34888 18624 34940 18630
rect 34888 18566 34940 18572
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35360 17202 35388 18702
rect 35452 18154 35480 22066
rect 35532 21888 35584 21894
rect 35532 21830 35584 21836
rect 35544 21690 35572 21830
rect 35532 21684 35584 21690
rect 35532 21626 35584 21632
rect 35532 21548 35584 21554
rect 35584 21508 35664 21536
rect 35532 21490 35584 21496
rect 35532 20460 35584 20466
rect 35532 20402 35584 20408
rect 35544 19514 35572 20402
rect 35532 19508 35584 19514
rect 35532 19450 35584 19456
rect 35532 19372 35584 19378
rect 35636 19334 35664 21508
rect 35900 20800 35952 20806
rect 35900 20742 35952 20748
rect 35912 20466 35940 20742
rect 35900 20460 35952 20466
rect 35900 20402 35952 20408
rect 35912 20058 35940 20402
rect 35992 20324 36044 20330
rect 35992 20266 36044 20272
rect 35900 20052 35952 20058
rect 35900 19994 35952 20000
rect 35584 19320 35664 19334
rect 35532 19314 35664 19320
rect 35544 19306 35664 19314
rect 35544 18766 35572 19306
rect 35532 18760 35584 18766
rect 35532 18702 35584 18708
rect 35440 18148 35492 18154
rect 35440 18090 35492 18096
rect 35544 17202 35572 18702
rect 35716 18624 35768 18630
rect 35716 18566 35768 18572
rect 35728 18290 35756 18566
rect 35716 18284 35768 18290
rect 35716 18226 35768 18232
rect 35808 18284 35860 18290
rect 35808 18226 35860 18232
rect 34796 17196 34848 17202
rect 34796 17138 34848 17144
rect 35164 17196 35216 17202
rect 35164 17138 35216 17144
rect 35348 17196 35400 17202
rect 35532 17196 35584 17202
rect 35400 17156 35480 17184
rect 35348 17138 35400 17144
rect 34704 16652 34756 16658
rect 34704 16594 34756 16600
rect 34716 15434 34744 16594
rect 34808 16590 34836 17138
rect 35176 17105 35204 17138
rect 35162 17096 35218 17105
rect 35162 17031 35218 17040
rect 35348 16992 35400 16998
rect 35348 16934 35400 16940
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34796 16584 34848 16590
rect 34796 16526 34848 16532
rect 35072 16584 35124 16590
rect 35164 16584 35216 16590
rect 35072 16526 35124 16532
rect 35162 16552 35164 16561
rect 35216 16552 35218 16561
rect 35084 16425 35112 16526
rect 35162 16487 35218 16496
rect 35070 16416 35126 16425
rect 35070 16351 35126 16360
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34796 15496 34848 15502
rect 34796 15438 34848 15444
rect 34704 15428 34756 15434
rect 34704 15370 34756 15376
rect 34704 14272 34756 14278
rect 34704 14214 34756 14220
rect 34716 13326 34744 14214
rect 34808 14006 34836 15438
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35360 14618 35388 16934
rect 35452 16658 35480 17156
rect 35532 17138 35584 17144
rect 35440 16652 35492 16658
rect 35440 16594 35492 16600
rect 35544 16590 35572 17138
rect 35532 16584 35584 16590
rect 35532 16526 35584 16532
rect 35716 16448 35768 16454
rect 35716 16390 35768 16396
rect 35532 16244 35584 16250
rect 35532 16186 35584 16192
rect 35440 14884 35492 14890
rect 35440 14826 35492 14832
rect 35348 14612 35400 14618
rect 35348 14554 35400 14560
rect 35452 14482 35480 14826
rect 35440 14476 35492 14482
rect 35440 14418 35492 14424
rect 35164 14408 35216 14414
rect 35162 14376 35164 14385
rect 35216 14376 35218 14385
rect 35162 14311 35218 14320
rect 34796 14000 34848 14006
rect 34796 13942 34848 13948
rect 35176 13938 35204 14311
rect 35544 14074 35572 16186
rect 35728 16114 35756 16390
rect 35716 16108 35768 16114
rect 35716 16050 35768 16056
rect 35624 14544 35676 14550
rect 35624 14486 35676 14492
rect 35532 14068 35584 14074
rect 35532 14010 35584 14016
rect 35164 13932 35216 13938
rect 35164 13874 35216 13880
rect 35636 13870 35664 14486
rect 35716 14408 35768 14414
rect 35716 14350 35768 14356
rect 35728 14006 35756 14350
rect 35716 14000 35768 14006
rect 35716 13942 35768 13948
rect 35348 13864 35400 13870
rect 35348 13806 35400 13812
rect 35624 13864 35676 13870
rect 35624 13806 35676 13812
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34704 13320 34756 13326
rect 34704 13262 34756 13268
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34796 12096 34848 12102
rect 34796 12038 34848 12044
rect 34612 11892 34664 11898
rect 34612 11834 34664 11840
rect 34704 11756 34756 11762
rect 34704 11698 34756 11704
rect 34520 10192 34572 10198
rect 34520 10134 34572 10140
rect 34520 10056 34572 10062
rect 34520 9998 34572 10004
rect 34428 8016 34480 8022
rect 34428 7958 34480 7964
rect 34532 7546 34560 9998
rect 34612 8356 34664 8362
rect 34612 8298 34664 8304
rect 34624 7750 34652 8298
rect 34612 7744 34664 7750
rect 34612 7686 34664 7692
rect 34520 7540 34572 7546
rect 34520 7482 34572 7488
rect 34152 6928 34204 6934
rect 34152 6870 34204 6876
rect 33968 6792 34020 6798
rect 33968 6734 34020 6740
rect 34716 6390 34744 11698
rect 34808 11082 34836 12038
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34796 11076 34848 11082
rect 34796 11018 34848 11024
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 35360 9110 35388 13806
rect 35728 13394 35756 13942
rect 35820 13802 35848 18226
rect 36004 18154 36032 20266
rect 36096 18902 36124 28018
rect 36648 26994 36676 28970
rect 36832 28626 36860 29650
rect 36820 28620 36872 28626
rect 36820 28562 36872 28568
rect 36912 27464 36964 27470
rect 36912 27406 36964 27412
rect 37096 27464 37148 27470
rect 37096 27406 37148 27412
rect 37186 27432 37242 27441
rect 36924 27130 36952 27406
rect 36912 27124 36964 27130
rect 36912 27066 36964 27072
rect 36360 26988 36412 26994
rect 36360 26930 36412 26936
rect 36636 26988 36688 26994
rect 36636 26930 36688 26936
rect 36372 26586 36400 26930
rect 36544 26784 36596 26790
rect 36544 26726 36596 26732
rect 36360 26580 36412 26586
rect 36360 26522 36412 26528
rect 36268 25152 36320 25158
rect 36268 25094 36320 25100
rect 36280 24682 36308 25094
rect 36268 24676 36320 24682
rect 36268 24618 36320 24624
rect 36176 23724 36228 23730
rect 36176 23666 36228 23672
rect 36188 23322 36216 23666
rect 36280 23594 36308 24618
rect 36556 23662 36584 26726
rect 36820 26376 36872 26382
rect 36820 26318 36872 26324
rect 36832 25294 36860 26318
rect 37108 26314 37136 27406
rect 37186 27367 37188 27376
rect 37240 27367 37242 27376
rect 37188 27338 37240 27344
rect 37292 26897 37320 30602
rect 38028 30598 38056 31214
rect 38016 30592 38068 30598
rect 38016 30534 38068 30540
rect 37832 30388 37884 30394
rect 37832 30330 37884 30336
rect 37844 30297 37872 30330
rect 37830 30288 37886 30297
rect 37830 30223 37886 30232
rect 37464 30048 37516 30054
rect 37464 29990 37516 29996
rect 37476 29646 37504 29990
rect 37844 29850 37872 30223
rect 38028 30190 38056 30534
rect 38016 30184 38068 30190
rect 38016 30126 38068 30132
rect 37832 29844 37884 29850
rect 37832 29786 37884 29792
rect 37464 29640 37516 29646
rect 37464 29582 37516 29588
rect 37924 29164 37976 29170
rect 37924 29106 37976 29112
rect 37740 29096 37792 29102
rect 37740 29038 37792 29044
rect 37752 28801 37780 29038
rect 37738 28792 37794 28801
rect 37738 28727 37794 28736
rect 37464 28484 37516 28490
rect 37464 28426 37516 28432
rect 37476 28218 37504 28426
rect 37936 28218 37964 29106
rect 37464 28212 37516 28218
rect 37464 28154 37516 28160
rect 37924 28212 37976 28218
rect 37924 28154 37976 28160
rect 38028 28014 38056 30126
rect 38200 28416 38252 28422
rect 38200 28358 38252 28364
rect 38212 28150 38240 28358
rect 38200 28144 38252 28150
rect 38200 28086 38252 28092
rect 38016 28008 38068 28014
rect 38016 27950 38068 27956
rect 38108 27396 38160 27402
rect 38108 27338 38160 27344
rect 37832 27056 37884 27062
rect 37832 26998 37884 27004
rect 37278 26888 37334 26897
rect 37278 26823 37334 26832
rect 37464 26784 37516 26790
rect 37464 26726 37516 26732
rect 37476 26382 37504 26726
rect 37844 26586 37872 26998
rect 38016 26920 38068 26926
rect 38016 26862 38068 26868
rect 37832 26580 37884 26586
rect 37832 26522 37884 26528
rect 38028 26489 38056 26862
rect 38014 26480 38070 26489
rect 38014 26415 38070 26424
rect 37464 26376 37516 26382
rect 37464 26318 37516 26324
rect 37096 26308 37148 26314
rect 37096 26250 37148 26256
rect 37924 25900 37976 25906
rect 37924 25842 37976 25848
rect 36820 25288 36872 25294
rect 36820 25230 36872 25236
rect 36832 24886 36860 25230
rect 37464 25220 37516 25226
rect 37464 25162 37516 25168
rect 37476 24954 37504 25162
rect 37832 25152 37884 25158
rect 37832 25094 37884 25100
rect 37844 24954 37872 25094
rect 37464 24948 37516 24954
rect 37464 24890 37516 24896
rect 37832 24948 37884 24954
rect 37832 24890 37884 24896
rect 36820 24880 36872 24886
rect 36820 24822 36872 24828
rect 36544 23656 36596 23662
rect 36544 23598 36596 23604
rect 36268 23588 36320 23594
rect 36268 23530 36320 23536
rect 36176 23316 36228 23322
rect 36176 23258 36228 23264
rect 36556 23254 36584 23598
rect 36544 23248 36596 23254
rect 36544 23190 36596 23196
rect 36360 22432 36412 22438
rect 36360 22374 36412 22380
rect 36372 21554 36400 22374
rect 36360 21548 36412 21554
rect 36360 21490 36412 21496
rect 36556 21418 36584 23190
rect 36832 23118 36860 24822
rect 37844 24721 37872 24890
rect 37936 24750 37964 25842
rect 38028 24750 38056 26415
rect 38120 26081 38148 27338
rect 38106 26072 38162 26081
rect 38106 26007 38162 26016
rect 38108 25832 38160 25838
rect 38108 25774 38160 25780
rect 37924 24744 37976 24750
rect 37830 24712 37886 24721
rect 37924 24686 37976 24692
rect 38016 24744 38068 24750
rect 38120 24721 38148 25774
rect 38016 24686 38068 24692
rect 38106 24712 38162 24721
rect 37830 24647 37886 24656
rect 37832 24200 37884 24206
rect 37832 24142 37884 24148
rect 37844 23866 37872 24142
rect 37740 23860 37792 23866
rect 37740 23802 37792 23808
rect 37832 23860 37884 23866
rect 37832 23802 37884 23808
rect 37752 23730 37780 23802
rect 37740 23724 37792 23730
rect 37740 23666 37792 23672
rect 37004 23520 37056 23526
rect 37004 23462 37056 23468
rect 37016 23118 37044 23462
rect 37752 23322 37780 23666
rect 37936 23594 37964 24686
rect 38028 23662 38056 24686
rect 38106 24647 38162 24656
rect 38108 24132 38160 24138
rect 38108 24074 38160 24080
rect 38016 23656 38068 23662
rect 38016 23598 38068 23604
rect 37924 23588 37976 23594
rect 37924 23530 37976 23536
rect 37740 23316 37792 23322
rect 37740 23258 37792 23264
rect 36820 23112 36872 23118
rect 36820 23054 36872 23060
rect 37004 23112 37056 23118
rect 37004 23054 37056 23060
rect 36832 22030 36860 23054
rect 37740 22636 37792 22642
rect 37740 22578 37792 22584
rect 36820 22024 36872 22030
rect 36820 21966 36872 21972
rect 36636 21888 36688 21894
rect 36636 21830 36688 21836
rect 36648 21554 36676 21830
rect 36636 21548 36688 21554
rect 36636 21490 36688 21496
rect 36544 21412 36596 21418
rect 36544 21354 36596 21360
rect 36556 20330 36584 21354
rect 36832 20942 36860 21966
rect 37464 21956 37516 21962
rect 37464 21898 37516 21904
rect 37476 21690 37504 21898
rect 37464 21684 37516 21690
rect 37464 21626 37516 21632
rect 37752 21622 37780 22578
rect 37740 21616 37792 21622
rect 37740 21558 37792 21564
rect 38028 21486 38056 23598
rect 38120 23361 38148 24074
rect 38106 23352 38162 23361
rect 38106 23287 38162 23296
rect 38108 22568 38160 22574
rect 38108 22510 38160 22516
rect 38120 22001 38148 22510
rect 38106 21992 38162 22001
rect 38106 21927 38162 21936
rect 38292 21888 38344 21894
rect 38292 21830 38344 21836
rect 38304 21554 38332 21830
rect 38292 21548 38344 21554
rect 38292 21490 38344 21496
rect 38016 21480 38068 21486
rect 38016 21422 38068 21428
rect 36820 20936 36872 20942
rect 36820 20878 36872 20884
rect 36544 20324 36596 20330
rect 36544 20266 36596 20272
rect 36832 19854 36860 20878
rect 37464 20868 37516 20874
rect 37464 20810 37516 20816
rect 37476 20602 37504 20810
rect 37648 20800 37700 20806
rect 37648 20742 37700 20748
rect 37464 20596 37516 20602
rect 37464 20538 37516 20544
rect 37660 20466 37688 20742
rect 37648 20460 37700 20466
rect 37648 20402 37700 20408
rect 36820 19848 36872 19854
rect 36820 19790 36872 19796
rect 36360 19236 36412 19242
rect 36360 19178 36412 19184
rect 36084 18896 36136 18902
rect 36084 18838 36136 18844
rect 36372 18290 36400 19178
rect 36832 18766 36860 19790
rect 37660 19446 37688 20402
rect 38028 20398 38056 21422
rect 38106 20632 38162 20641
rect 38106 20567 38162 20576
rect 38016 20392 38068 20398
rect 38016 20334 38068 20340
rect 37832 20324 37884 20330
rect 37832 20266 37884 20272
rect 37844 19854 37872 20266
rect 37832 19848 37884 19854
rect 37832 19790 37884 19796
rect 37648 19440 37700 19446
rect 37648 19382 37700 19388
rect 37740 19372 37792 19378
rect 37740 19314 37792 19320
rect 36820 18760 36872 18766
rect 36820 18702 36872 18708
rect 36360 18284 36412 18290
rect 36360 18226 36412 18232
rect 36176 18216 36228 18222
rect 36176 18158 36228 18164
rect 35992 18148 36044 18154
rect 35992 18090 36044 18096
rect 36188 13938 36216 18158
rect 36372 15706 36400 18226
rect 36636 18148 36688 18154
rect 36636 18090 36688 18096
rect 36648 17134 36676 18090
rect 36728 17808 36780 17814
rect 36728 17750 36780 17756
rect 36740 17202 36768 17750
rect 36728 17196 36780 17202
rect 36728 17138 36780 17144
rect 36636 17128 36688 17134
rect 36636 17070 36688 17076
rect 36648 15978 36676 17070
rect 36636 15972 36688 15978
rect 36636 15914 36688 15920
rect 36360 15700 36412 15706
rect 36360 15642 36412 15648
rect 36452 14340 36504 14346
rect 36452 14282 36504 14288
rect 36464 14006 36492 14282
rect 36452 14000 36504 14006
rect 36452 13942 36504 13948
rect 36176 13932 36228 13938
rect 36176 13874 36228 13880
rect 35808 13796 35860 13802
rect 35808 13738 35860 13744
rect 36740 13530 36768 17138
rect 36832 16658 36860 18702
rect 37464 18692 37516 18698
rect 37464 18634 37516 18640
rect 37476 18426 37504 18634
rect 37464 18420 37516 18426
rect 37464 18362 37516 18368
rect 37752 18358 37780 19314
rect 37832 18624 37884 18630
rect 37832 18566 37884 18572
rect 37844 18426 37872 18566
rect 37832 18420 37884 18426
rect 37832 18362 37884 18368
rect 37740 18352 37792 18358
rect 37740 18294 37792 18300
rect 38028 18222 38056 20334
rect 38120 19922 38148 20567
rect 38108 19916 38160 19922
rect 38108 19858 38160 19864
rect 38108 19372 38160 19378
rect 38108 19314 38160 19320
rect 38120 19281 38148 19314
rect 38106 19272 38162 19281
rect 38106 19207 38162 19216
rect 38016 18216 38068 18222
rect 38016 18158 38068 18164
rect 37832 17672 37884 17678
rect 37832 17614 37884 17620
rect 37844 17338 37872 17614
rect 37740 17332 37792 17338
rect 37740 17274 37792 17280
rect 37832 17332 37884 17338
rect 37832 17274 37884 17280
rect 37752 17202 37780 17274
rect 37740 17196 37792 17202
rect 37740 17138 37792 17144
rect 37096 16992 37148 16998
rect 37096 16934 37148 16940
rect 36820 16652 36872 16658
rect 36820 16594 36872 16600
rect 37108 16590 37136 16934
rect 37752 16794 37780 17138
rect 38028 17134 38056 18158
rect 38106 17912 38162 17921
rect 38106 17847 38162 17856
rect 38120 17746 38148 17847
rect 38108 17740 38160 17746
rect 38108 17682 38160 17688
rect 38016 17128 38068 17134
rect 38016 17070 38068 17076
rect 37740 16788 37792 16794
rect 37740 16730 37792 16736
rect 37096 16584 37148 16590
rect 37096 16526 37148 16532
rect 37832 16516 37884 16522
rect 37832 16458 37884 16464
rect 37844 16250 37872 16458
rect 37832 16244 37884 16250
rect 37884 16204 37964 16232
rect 37832 16186 37884 16192
rect 37832 15972 37884 15978
rect 37832 15914 37884 15920
rect 37188 15904 37240 15910
rect 37188 15846 37240 15852
rect 37200 14414 37228 15846
rect 37844 15502 37872 15914
rect 37832 15496 37884 15502
rect 37832 15438 37884 15444
rect 37936 14618 37964 16204
rect 38028 16046 38056 17070
rect 38106 16552 38162 16561
rect 38106 16487 38162 16496
rect 38016 16040 38068 16046
rect 38016 15982 38068 15988
rect 38028 15366 38056 15982
rect 38120 15570 38148 16487
rect 38108 15564 38160 15570
rect 38108 15506 38160 15512
rect 38016 15360 38068 15366
rect 38016 15302 38068 15308
rect 38106 15192 38162 15201
rect 38106 15127 38162 15136
rect 38120 15094 38148 15127
rect 38108 15088 38160 15094
rect 38108 15030 38160 15036
rect 37924 14612 37976 14618
rect 37924 14554 37976 14560
rect 37188 14408 37240 14414
rect 37188 14350 37240 14356
rect 38292 13864 38344 13870
rect 38290 13832 38292 13841
rect 38344 13832 38346 13841
rect 38290 13767 38346 13776
rect 36728 13524 36780 13530
rect 36728 13466 36780 13472
rect 35716 13388 35768 13394
rect 35716 13330 35768 13336
rect 35532 12640 35584 12646
rect 35532 12582 35584 12588
rect 35544 12434 35572 12582
rect 35544 12406 35664 12434
rect 35532 9580 35584 9586
rect 35532 9522 35584 9528
rect 35348 9104 35400 9110
rect 35348 9046 35400 9052
rect 35440 8968 35492 8974
rect 35440 8910 35492 8916
rect 35348 8492 35400 8498
rect 35348 8434 35400 8440
rect 34796 8424 34848 8430
rect 34796 8366 34848 8372
rect 34808 7818 34836 8366
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35360 8090 35388 8434
rect 35348 8084 35400 8090
rect 35348 8026 35400 8032
rect 35256 7948 35308 7954
rect 35256 7890 35308 7896
rect 35348 7948 35400 7954
rect 35348 7890 35400 7896
rect 34796 7812 34848 7818
rect 34796 7754 34848 7760
rect 35268 7750 35296 7890
rect 35164 7744 35216 7750
rect 35164 7686 35216 7692
rect 35256 7744 35308 7750
rect 35256 7686 35308 7692
rect 35176 7410 35204 7686
rect 35072 7404 35124 7410
rect 35072 7346 35124 7352
rect 35164 7404 35216 7410
rect 35164 7346 35216 7352
rect 35084 7290 35112 7346
rect 35360 7290 35388 7890
rect 35084 7262 35388 7290
rect 34796 7200 34848 7206
rect 34796 7142 34848 7148
rect 34808 6474 34836 7142
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35072 6792 35124 6798
rect 35072 6734 35124 6740
rect 34808 6446 34928 6474
rect 34900 6390 34928 6446
rect 33876 6384 33928 6390
rect 33876 6326 33928 6332
rect 34704 6384 34756 6390
rect 34704 6326 34756 6332
rect 34888 6384 34940 6390
rect 34888 6326 34940 6332
rect 33784 6316 33836 6322
rect 33784 6258 33836 6264
rect 33048 5772 33100 5778
rect 33048 5714 33100 5720
rect 31668 5704 31720 5710
rect 31668 5646 31720 5652
rect 31680 5250 31708 5646
rect 31680 5234 31800 5250
rect 31680 5228 31812 5234
rect 31680 5222 31760 5228
rect 31760 5170 31812 5176
rect 32588 5228 32640 5234
rect 32588 5170 32640 5176
rect 32220 5160 32272 5166
rect 32220 5102 32272 5108
rect 30932 4820 30984 4826
rect 30932 4762 30984 4768
rect 30944 4282 30972 4762
rect 32232 4758 32260 5102
rect 32600 4826 32628 5170
rect 32588 4820 32640 4826
rect 32588 4762 32640 4768
rect 32220 4752 32272 4758
rect 32220 4694 32272 4700
rect 33060 4690 33088 5714
rect 33692 5568 33744 5574
rect 33692 5510 33744 5516
rect 33600 5160 33652 5166
rect 33600 5102 33652 5108
rect 33048 4684 33100 4690
rect 33048 4626 33100 4632
rect 30932 4276 30984 4282
rect 30932 4218 30984 4224
rect 30472 4208 30524 4214
rect 30472 4150 30524 4156
rect 33612 4146 33640 5102
rect 33704 4146 33732 5510
rect 33796 5370 33824 6258
rect 33888 5642 33916 6326
rect 35084 6118 35112 6734
rect 35360 6390 35388 7262
rect 35452 7002 35480 8910
rect 35544 7954 35572 9522
rect 35532 7948 35584 7954
rect 35532 7890 35584 7896
rect 35440 6996 35492 7002
rect 35440 6938 35492 6944
rect 35532 6792 35584 6798
rect 35532 6734 35584 6740
rect 35544 6458 35572 6734
rect 35532 6452 35584 6458
rect 35532 6394 35584 6400
rect 35348 6384 35400 6390
rect 35348 6326 35400 6332
rect 35636 6322 35664 12406
rect 35728 12306 35756 13330
rect 38292 12640 38344 12646
rect 38292 12582 38344 12588
rect 38304 12481 38332 12582
rect 38290 12472 38346 12481
rect 38290 12407 38346 12416
rect 35716 12300 35768 12306
rect 35716 12242 35768 12248
rect 38200 12232 38252 12238
rect 38200 12174 38252 12180
rect 35808 12164 35860 12170
rect 35808 12106 35860 12112
rect 37464 12164 37516 12170
rect 37464 12106 37516 12112
rect 35716 12096 35768 12102
rect 35716 12038 35768 12044
rect 35728 11558 35756 12038
rect 35820 11694 35848 12106
rect 37476 11898 37504 12106
rect 37832 12096 37884 12102
rect 37832 12038 37884 12044
rect 37844 11898 37872 12038
rect 37464 11892 37516 11898
rect 37464 11834 37516 11840
rect 37832 11892 37884 11898
rect 37832 11834 37884 11840
rect 35900 11756 35952 11762
rect 35900 11698 35952 11704
rect 35808 11688 35860 11694
rect 35808 11630 35860 11636
rect 35716 11552 35768 11558
rect 35716 11494 35768 11500
rect 35440 6316 35492 6322
rect 35440 6258 35492 6264
rect 35624 6316 35676 6322
rect 35624 6258 35676 6264
rect 35072 6112 35124 6118
rect 35072 6054 35124 6060
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35452 5914 35480 6258
rect 35440 5908 35492 5914
rect 35440 5850 35492 5856
rect 33876 5636 33928 5642
rect 33876 5578 33928 5584
rect 35348 5636 35400 5642
rect 35348 5578 35400 5584
rect 33784 5364 33836 5370
rect 33784 5306 33836 5312
rect 33796 4622 33824 5306
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 33784 4616 33836 4622
rect 33784 4558 33836 4564
rect 33600 4140 33652 4146
rect 33600 4082 33652 4088
rect 33692 4140 33744 4146
rect 33692 4082 33744 4088
rect 29552 4072 29604 4078
rect 29552 4014 29604 4020
rect 30288 4072 30340 4078
rect 30288 4014 30340 4020
rect 35360 3942 35388 5578
rect 35728 5574 35756 11494
rect 35820 11354 35848 11630
rect 35808 11348 35860 11354
rect 35808 11290 35860 11296
rect 35912 10062 35940 11698
rect 38212 11694 38240 12174
rect 38200 11688 38252 11694
rect 38200 11630 38252 11636
rect 36176 11620 36228 11626
rect 36176 11562 36228 11568
rect 36188 10130 36216 11562
rect 38106 11112 38162 11121
rect 37464 11076 37516 11082
rect 38106 11047 38162 11056
rect 37464 11018 37516 11024
rect 37476 10810 37504 11018
rect 37832 11008 37884 11014
rect 37832 10950 37884 10956
rect 37464 10804 37516 10810
rect 37464 10746 37516 10752
rect 37844 10674 37872 10950
rect 38016 10736 38068 10742
rect 38016 10678 38068 10684
rect 37372 10668 37424 10674
rect 37372 10610 37424 10616
rect 37832 10668 37884 10674
rect 37832 10610 37884 10616
rect 37384 10130 37412 10610
rect 37830 10160 37886 10169
rect 36176 10124 36228 10130
rect 36176 10066 36228 10072
rect 37372 10124 37424 10130
rect 37830 10095 37886 10104
rect 37372 10066 37424 10072
rect 35900 10056 35952 10062
rect 35900 9998 35952 10004
rect 35912 8974 35940 9998
rect 36188 9110 36216 10066
rect 37844 10062 37872 10095
rect 37832 10056 37884 10062
rect 37832 9998 37884 10004
rect 37830 9888 37886 9897
rect 37830 9823 37886 9832
rect 37844 9586 37872 9823
rect 37832 9580 37884 9586
rect 37832 9522 37884 9528
rect 36176 9104 36228 9110
rect 36176 9046 36228 9052
rect 36084 9036 36136 9042
rect 36084 8978 36136 8984
rect 35900 8968 35952 8974
rect 35900 8910 35952 8916
rect 36096 8634 36124 8978
rect 37740 8900 37792 8906
rect 37740 8842 37792 8848
rect 37752 8634 37780 8842
rect 36084 8628 36136 8634
rect 36084 8570 36136 8576
rect 37740 8628 37792 8634
rect 37740 8570 37792 8576
rect 36096 7818 36124 8570
rect 37188 8356 37240 8362
rect 37188 8298 37240 8304
rect 37200 7886 37228 8298
rect 37752 8106 37780 8570
rect 37924 8424 37976 8430
rect 37924 8366 37976 8372
rect 37752 8090 37872 8106
rect 37752 8084 37884 8090
rect 37752 8078 37832 8084
rect 37832 8026 37884 8032
rect 36728 7880 36780 7886
rect 36728 7822 36780 7828
rect 37188 7880 37240 7886
rect 37188 7822 37240 7828
rect 36084 7812 36136 7818
rect 36084 7754 36136 7760
rect 35900 7744 35952 7750
rect 35900 7686 35952 7692
rect 35716 5568 35768 5574
rect 35716 5510 35768 5516
rect 35532 5228 35584 5234
rect 35532 5170 35584 5176
rect 35544 4826 35572 5170
rect 35532 4820 35584 4826
rect 35532 4762 35584 4768
rect 35912 4690 35940 7686
rect 36740 6866 36768 7822
rect 37936 7750 37964 8366
rect 37924 7744 37976 7750
rect 37924 7686 37976 7692
rect 38028 7546 38056 10678
rect 38120 10130 38148 11047
rect 38212 10606 38240 11630
rect 38200 10600 38252 10606
rect 38200 10542 38252 10548
rect 38108 10124 38160 10130
rect 38108 10066 38160 10072
rect 38106 9752 38162 9761
rect 38106 9687 38162 9696
rect 38120 9654 38148 9687
rect 38108 9648 38160 9654
rect 38108 9590 38160 9596
rect 38108 8900 38160 8906
rect 38108 8842 38160 8848
rect 38120 8401 38148 8842
rect 38212 8430 38240 10542
rect 38200 8424 38252 8430
rect 38106 8392 38162 8401
rect 38200 8366 38252 8372
rect 38106 8327 38162 8336
rect 37832 7540 37884 7546
rect 37832 7482 37884 7488
rect 38016 7540 38068 7546
rect 38016 7482 38068 7488
rect 37004 7200 37056 7206
rect 37004 7142 37056 7148
rect 36728 6860 36780 6866
rect 36728 6802 36780 6808
rect 36636 6112 36688 6118
rect 36636 6054 36688 6060
rect 36648 5370 36676 6054
rect 36740 5778 36768 6802
rect 37016 6798 37044 7142
rect 37844 7002 37872 7482
rect 38016 7336 38068 7342
rect 38016 7278 38068 7284
rect 37832 6996 37884 7002
rect 37832 6938 37884 6944
rect 37004 6792 37056 6798
rect 37004 6734 37056 6740
rect 36728 5772 36780 5778
rect 36728 5714 36780 5720
rect 37464 5636 37516 5642
rect 37464 5578 37516 5584
rect 37476 5370 37504 5578
rect 37924 5568 37976 5574
rect 37924 5510 37976 5516
rect 36636 5364 36688 5370
rect 36636 5306 36688 5312
rect 37464 5364 37516 5370
rect 37464 5306 37516 5312
rect 35900 4684 35952 4690
rect 35900 4626 35952 4632
rect 35912 4486 35940 4626
rect 36648 4622 36676 5306
rect 37936 5302 37964 5510
rect 37924 5296 37976 5302
rect 37924 5238 37976 5244
rect 38028 5166 38056 7278
rect 38106 7032 38162 7041
rect 38106 6967 38162 6976
rect 38120 6390 38148 6967
rect 38108 6384 38160 6390
rect 38108 6326 38160 6332
rect 38292 6248 38344 6254
rect 38292 6190 38344 6196
rect 38304 5914 38332 6190
rect 38292 5908 38344 5914
rect 38292 5850 38344 5856
rect 38106 5672 38162 5681
rect 38106 5607 38162 5616
rect 38016 5160 38068 5166
rect 38016 5102 38068 5108
rect 38028 4758 38056 5102
rect 38016 4752 38068 4758
rect 38016 4694 38068 4700
rect 38120 4690 38148 5607
rect 38304 5370 38332 5850
rect 38292 5364 38344 5370
rect 38292 5306 38344 5312
rect 38108 4684 38160 4690
rect 38108 4626 38160 4632
rect 36636 4616 36688 4622
rect 36636 4558 36688 4564
rect 35900 4480 35952 4486
rect 35900 4422 35952 4428
rect 38106 4312 38162 4321
rect 38106 4247 38162 4256
rect 38120 4146 38148 4247
rect 38108 4140 38160 4146
rect 38108 4082 38160 4088
rect 29368 3936 29420 3942
rect 29368 3878 29420 3884
rect 35348 3936 35400 3942
rect 35348 3878 35400 3884
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 38108 2984 38160 2990
rect 38106 2952 38108 2961
rect 38160 2952 38162 2961
rect 38106 2887 38162 2896
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 27344 2440 27396 2446
rect 27344 2382 27396 2388
rect 38108 2372 38160 2378
rect 38108 2314 38160 2320
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 38120 1601 38148 2314
rect 38106 1592 38162 1601
rect 38106 1527 38162 1536
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 5722 33940 5724 33960
rect 5724 33940 5776 33960
rect 5776 33940 5778 33960
rect 5722 33904 5778 33940
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4066 28464 4122 28520
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4802 27104 4858 27160
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 5170 31728 5226 31784
rect 5446 28484 5502 28520
rect 5446 28464 5448 28484
rect 5448 28464 5500 28484
rect 5500 28464 5502 28484
rect 5814 28464 5870 28520
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 5170 27104 5226 27160
rect 5998 26424 6054 26480
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 9218 31728 9274 31784
rect 8482 28484 8538 28520
rect 8482 28464 8484 28484
rect 8484 28464 8536 28484
rect 8536 28464 8538 28484
rect 9494 32272 9550 32328
rect 9218 26732 9220 26752
rect 9220 26732 9272 26752
rect 9272 26732 9274 26752
rect 9218 26696 9274 26732
rect 9586 27396 9642 27432
rect 9586 27376 9588 27396
rect 9588 27376 9640 27396
rect 9640 27376 9642 27396
rect 9494 26424 9550 26480
rect 10414 31728 10470 31784
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 9862 22616 9918 22672
rect 11610 31728 11666 31784
rect 12162 31864 12218 31920
rect 12162 31728 12218 31784
rect 8850 15156 8906 15192
rect 8850 15136 8852 15156
rect 8852 15136 8904 15156
rect 8904 15136 8906 15156
rect 10414 20304 10470 20360
rect 11794 22636 11850 22672
rect 11794 22616 11796 22636
rect 11796 22616 11848 22636
rect 11848 22616 11850 22636
rect 12346 31864 12402 31920
rect 12622 32408 12678 32464
rect 13542 32272 13598 32328
rect 13726 30640 13782 30696
rect 13726 27376 13782 27432
rect 14370 32308 14372 32328
rect 14372 32308 14424 32328
rect 14424 32308 14426 32328
rect 14370 32272 14426 32308
rect 14554 30232 14610 30288
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 16026 34040 16082 34096
rect 15750 29588 15752 29608
rect 15752 29588 15804 29608
rect 15804 29588 15806 29608
rect 15750 29552 15806 29588
rect 15106 25472 15162 25528
rect 17590 32272 17646 32328
rect 17406 32172 17408 32192
rect 17408 32172 17460 32192
rect 17460 32172 17462 32192
rect 17406 32136 17462 32172
rect 17314 31764 17316 31784
rect 17316 31764 17368 31784
rect 17368 31764 17370 31784
rect 17314 31728 17370 31764
rect 17682 32136 17738 32192
rect 16670 29552 16726 29608
rect 17406 29044 17408 29064
rect 17408 29044 17460 29064
rect 17460 29044 17462 29064
rect 17406 29008 17462 29044
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 14002 12280 14058 12336
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 15198 15020 15254 15056
rect 15198 15000 15200 15020
rect 15200 15000 15252 15020
rect 15252 15000 15254 15020
rect 15750 20304 15806 20360
rect 17222 22616 17278 22672
rect 19706 34992 19762 35048
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19522 34176 19578 34232
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19706 31728 19762 31784
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19890 30912 19946 30968
rect 19706 30776 19762 30832
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19430 29164 19486 29200
rect 19430 29144 19432 29164
rect 19432 29144 19484 29164
rect 19484 29144 19486 29164
rect 19982 28872 20038 28928
rect 19338 26288 19394 26344
rect 14370 6704 14426 6760
rect 14738 6740 14740 6760
rect 14740 6740 14792 6760
rect 14792 6740 14794 6760
rect 14738 6704 14794 6740
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 17222 17856 17278 17912
rect 17222 12300 17278 12336
rect 17222 12280 17224 12300
rect 17224 12280 17276 12300
rect 17276 12280 17278 12300
rect 17866 15036 17868 15056
rect 17868 15036 17920 15056
rect 17920 15036 17922 15056
rect 17866 15000 17922 15036
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19982 28076 20038 28112
rect 19982 28056 19984 28076
rect 19984 28056 20036 28076
rect 20036 28056 20038 28076
rect 20166 31048 20222 31104
rect 20258 29028 20314 29064
rect 20258 29008 20260 29028
rect 20260 29008 20312 29028
rect 20312 29008 20314 29028
rect 19982 27376 20038 27432
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 20166 26832 20222 26888
rect 20534 30676 20536 30696
rect 20536 30676 20588 30696
rect 20588 30676 20590 30696
rect 20534 30640 20590 30676
rect 20902 32680 20958 32736
rect 20810 30776 20866 30832
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19430 20440 19486 20496
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 20718 23160 20774 23216
rect 20534 21936 20590 21992
rect 20534 20032 20590 20088
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 20074 18400 20130 18456
rect 19522 17620 19524 17640
rect 19524 17620 19576 17640
rect 19576 17620 19578 17640
rect 19522 17584 19578 17620
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19522 14320 19578 14376
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19430 13912 19486 13968
rect 18694 6704 18750 6760
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19706 12844 19762 12880
rect 19706 12824 19708 12844
rect 19708 12824 19760 12844
rect 19760 12824 19762 12844
rect 20258 12824 20314 12880
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 20994 26424 21050 26480
rect 21178 26832 21234 26888
rect 21822 33904 21878 33960
rect 22742 33940 22744 33960
rect 22744 33940 22796 33960
rect 22796 33940 22798 33960
rect 21822 32292 21878 32328
rect 21822 32272 21824 32292
rect 21824 32272 21876 32292
rect 21876 32272 21878 32292
rect 22742 33904 22798 33940
rect 21178 25880 21234 25936
rect 21086 24112 21142 24168
rect 21546 25744 21602 25800
rect 21638 22924 21640 22944
rect 21640 22924 21692 22944
rect 21692 22924 21694 22944
rect 21638 22888 21694 22924
rect 22374 30640 22430 30696
rect 21914 29008 21970 29064
rect 21914 25064 21970 25120
rect 23754 34176 23810 34232
rect 23110 32272 23166 32328
rect 22374 26732 22376 26752
rect 22376 26732 22428 26752
rect 22428 26732 22430 26752
rect 22374 26696 22430 26732
rect 23386 30640 23442 30696
rect 21362 20304 21418 20360
rect 21270 17448 21326 17504
rect 21086 17176 21142 17232
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 22742 24656 22798 24712
rect 22742 24384 22798 24440
rect 21914 19780 21970 19816
rect 21914 19760 21916 19780
rect 21916 19760 21968 19780
rect 21968 19760 21970 19780
rect 21914 18808 21970 18864
rect 22006 17720 22062 17776
rect 23018 27104 23074 27160
rect 23294 28056 23350 28112
rect 23478 27412 23480 27432
rect 23480 27412 23532 27432
rect 23532 27412 23534 27432
rect 23478 27376 23534 27412
rect 23386 27104 23442 27160
rect 23294 26732 23296 26752
rect 23296 26732 23348 26752
rect 23348 26732 23350 26752
rect 23294 26696 23350 26732
rect 23662 26288 23718 26344
rect 23294 23432 23350 23488
rect 22834 21664 22890 21720
rect 21454 14456 21510 14512
rect 21454 12588 21456 12608
rect 21456 12588 21508 12608
rect 21508 12588 21510 12608
rect 21454 12552 21510 12588
rect 22558 18400 22614 18456
rect 22650 17856 22706 17912
rect 24030 32272 24086 32328
rect 24306 29280 24362 29336
rect 23754 24656 23810 24712
rect 23478 22616 23534 22672
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 25042 34992 25098 35048
rect 24858 30776 24914 30832
rect 25226 32408 25282 32464
rect 25226 29280 25282 29336
rect 25134 29144 25190 29200
rect 25686 31728 25742 31784
rect 25502 29824 25558 29880
rect 24490 25900 24546 25936
rect 24490 25880 24492 25900
rect 24492 25880 24544 25900
rect 24544 25880 24546 25900
rect 24674 25472 24730 25528
rect 24950 27376 25006 27432
rect 25134 26832 25190 26888
rect 26238 32272 26294 32328
rect 26422 30776 26478 30832
rect 24858 25764 24914 25800
rect 24858 25744 24860 25764
rect 24860 25744 24912 25764
rect 24912 25744 24914 25764
rect 24030 20304 24086 20360
rect 23938 19760 23994 19816
rect 24306 19372 24362 19408
rect 24306 19352 24308 19372
rect 24308 19352 24360 19372
rect 24360 19352 24362 19372
rect 25778 26424 25834 26480
rect 25962 25880 26018 25936
rect 25686 24384 25742 24440
rect 24674 17448 24730 17504
rect 25226 20032 25282 20088
rect 26514 29844 26570 29880
rect 26514 29824 26516 29844
rect 26516 29824 26568 29844
rect 26568 29824 26570 29844
rect 26514 24112 26570 24168
rect 26054 20576 26110 20632
rect 25686 20032 25742 20088
rect 25410 12844 25466 12880
rect 25410 12824 25412 12844
rect 25412 12824 25464 12844
rect 25464 12824 25466 12844
rect 25870 13640 25926 13696
rect 26790 23160 26846 23216
rect 27710 30676 27712 30696
rect 27712 30676 27764 30696
rect 27764 30676 27766 30696
rect 27710 30640 27766 30676
rect 27710 30232 27766 30288
rect 27618 29008 27674 29064
rect 26974 22888 27030 22944
rect 26790 21972 26792 21992
rect 26792 21972 26844 21992
rect 26844 21972 26846 21992
rect 26790 21936 26846 21972
rect 26238 19352 26294 19408
rect 27618 27648 27674 27704
rect 27526 26832 27582 26888
rect 27618 26152 27674 26208
rect 27434 24792 27490 24848
rect 27342 23568 27398 23624
rect 27066 20748 27068 20768
rect 27068 20748 27120 20768
rect 27120 20748 27122 20768
rect 27066 20712 27122 20748
rect 27066 19352 27122 19408
rect 36818 38256 36874 38312
rect 28906 34584 28962 34640
rect 27986 26016 28042 26072
rect 28262 26152 28318 26208
rect 30746 35028 30748 35048
rect 30748 35028 30800 35048
rect 30800 35028 30802 35048
rect 28906 31748 28962 31784
rect 28906 31728 28908 31748
rect 28908 31728 28960 31748
rect 28960 31728 28962 31748
rect 28722 27784 28778 27840
rect 28814 27648 28870 27704
rect 27710 23060 27712 23080
rect 27712 23060 27764 23080
rect 27764 23060 27766 23080
rect 27710 23024 27766 23060
rect 27158 17720 27214 17776
rect 26514 16360 26570 16416
rect 26238 15272 26294 15328
rect 27158 15136 27214 15192
rect 27434 17604 27490 17640
rect 27434 17584 27436 17604
rect 27436 17584 27488 17604
rect 27488 17584 27490 17604
rect 27434 16768 27490 16824
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 27894 17040 27950 17096
rect 27802 12588 27804 12608
rect 27804 12588 27856 12608
rect 27856 12588 27858 12608
rect 27802 12552 27858 12588
rect 27802 12280 27858 12336
rect 28262 24928 28318 24984
rect 29090 25064 29146 25120
rect 28722 23704 28778 23760
rect 28630 23296 28686 23352
rect 28262 23160 28318 23216
rect 28262 22636 28318 22672
rect 28262 22616 28264 22636
rect 28264 22616 28316 22636
rect 28316 22616 28318 22636
rect 28262 20340 28264 20360
rect 28264 20340 28316 20360
rect 28316 20340 28318 20360
rect 28262 20304 28318 20340
rect 28538 21800 28594 21856
rect 28354 13640 28410 13696
rect 28262 12280 28318 12336
rect 28814 22208 28870 22264
rect 29366 29180 29368 29200
rect 29368 29180 29420 29200
rect 29420 29180 29422 29200
rect 29366 29144 29422 29180
rect 29550 29008 29606 29064
rect 30102 33768 30158 33824
rect 30746 34992 30802 35028
rect 31390 34040 31446 34096
rect 31298 33940 31300 33960
rect 31300 33940 31352 33960
rect 31352 33940 31354 33960
rect 30746 33396 30748 33416
rect 30748 33396 30800 33416
rect 30800 33396 30802 33416
rect 30746 33360 30802 33396
rect 30102 32852 30104 32872
rect 30104 32852 30156 32872
rect 30156 32852 30158 32872
rect 30102 32816 30158 32852
rect 30102 32716 30104 32736
rect 30104 32716 30156 32736
rect 30156 32716 30158 32736
rect 30102 32680 30158 32716
rect 30470 30912 30526 30968
rect 30378 29960 30434 30016
rect 30746 31184 30802 31240
rect 31298 33904 31354 33940
rect 31298 32716 31300 32736
rect 31300 32716 31352 32736
rect 31352 32716 31354 32736
rect 31298 32680 31354 32716
rect 30378 29144 30434 29200
rect 30102 26968 30158 27024
rect 29734 26288 29790 26344
rect 29366 22636 29422 22672
rect 29366 22616 29368 22636
rect 29368 22616 29420 22636
rect 29420 22616 29422 22636
rect 30194 26832 30250 26888
rect 29366 21664 29422 21720
rect 28538 16632 28594 16688
rect 28722 17212 28724 17232
rect 28724 17212 28776 17232
rect 28776 17212 28778 17232
rect 28722 17176 28778 17212
rect 28998 19292 29054 19348
rect 28998 18944 29054 19000
rect 28906 16788 28962 16824
rect 28906 16768 28908 16788
rect 28908 16768 28960 16788
rect 28960 16768 28962 16788
rect 28906 16632 28962 16688
rect 28906 16396 28908 16416
rect 28908 16396 28960 16416
rect 28960 16396 28962 16416
rect 28906 16360 28962 16396
rect 29642 20460 29698 20496
rect 29642 20440 29644 20460
rect 29644 20440 29696 20460
rect 29696 20440 29698 20460
rect 29090 13640 29146 13696
rect 30286 23432 30342 23488
rect 31022 30268 31024 30288
rect 31024 30268 31076 30288
rect 31076 30268 31078 30288
rect 31022 30232 31078 30268
rect 31022 29688 31078 29744
rect 31022 23704 31078 23760
rect 29734 16632 29790 16688
rect 29918 17584 29974 17640
rect 31666 32444 31668 32464
rect 31668 32444 31720 32464
rect 31720 32444 31722 32464
rect 31666 32408 31722 32444
rect 31942 32852 31944 32872
rect 31944 32852 31996 32872
rect 31996 32852 31998 32872
rect 31942 32816 31998 32852
rect 31758 31320 31814 31376
rect 31758 26968 31814 27024
rect 31758 24792 31814 24848
rect 32126 26852 32182 26888
rect 32126 26832 32128 26852
rect 32128 26832 32180 26852
rect 32180 26832 32182 26852
rect 31850 16532 31852 16552
rect 31852 16532 31904 16552
rect 31904 16532 31906 16552
rect 30930 14456 30986 14512
rect 31850 16496 31906 16532
rect 31482 16360 31538 16416
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34794 35128 34850 35184
rect 34426 33768 34482 33824
rect 34334 33516 34390 33552
rect 34334 33496 34336 33516
rect 34336 33496 34388 33516
rect 34388 33496 34390 33516
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34610 31356 34612 31376
rect 34612 31356 34664 31376
rect 34664 31356 34666 31376
rect 34610 31320 34666 31356
rect 32402 26444 32458 26480
rect 32402 26424 32404 26444
rect 32404 26424 32456 26444
rect 32456 26424 32458 26444
rect 32402 24656 32458 24712
rect 32678 24846 32734 24848
rect 32678 24794 32680 24846
rect 32680 24794 32732 24846
rect 32732 24794 32734 24846
rect 32678 24792 32734 24794
rect 33322 23296 33378 23352
rect 32678 19372 32734 19408
rect 32678 19352 32680 19372
rect 32680 19352 32732 19372
rect 32732 19352 32734 19372
rect 33322 19372 33378 19408
rect 33322 19352 33324 19372
rect 33324 19352 33376 19372
rect 33376 19352 33378 19372
rect 33322 18692 33378 18728
rect 33322 18672 33324 18692
rect 33324 18672 33376 18692
rect 33376 18672 33378 18692
rect 33046 14320 33102 14376
rect 34610 26696 34666 26752
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34794 31320 34850 31376
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34886 29688 34942 29744
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 35898 33516 35954 33552
rect 35898 33496 35900 33516
rect 35900 33496 35952 33516
rect 35952 33496 35954 33516
rect 35530 30640 35586 30696
rect 35438 29708 35494 29744
rect 35438 29688 35440 29708
rect 35440 29688 35492 29708
rect 35492 29688 35494 29708
rect 36726 36896 36782 36952
rect 38106 35536 38162 35592
rect 35898 30252 35954 30288
rect 38106 34176 38162 34232
rect 35898 30232 35900 30252
rect 35900 30232 35952 30252
rect 35952 30232 35954 30252
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 38106 32816 38162 32872
rect 38106 31456 38162 31512
rect 37002 30096 37058 30152
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34518 23060 34520 23080
rect 34520 23060 34572 23080
rect 34572 23060 34574 23080
rect 34518 23024 34574 23060
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 35530 23160 35586 23216
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35162 18808 35218 18864
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 35162 17040 35218 17096
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35162 16532 35164 16552
rect 35164 16532 35216 16552
rect 35216 16532 35218 16552
rect 35162 16496 35218 16532
rect 35070 16360 35126 16416
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 35162 14356 35164 14376
rect 35164 14356 35216 14376
rect 35216 14356 35218 14376
rect 35162 14320 35218 14356
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 37186 27396 37242 27432
rect 37186 27376 37188 27396
rect 37188 27376 37240 27396
rect 37240 27376 37242 27396
rect 37830 30232 37886 30288
rect 37738 28736 37794 28792
rect 37278 26832 37334 26888
rect 38014 26424 38070 26480
rect 38106 26016 38162 26072
rect 37830 24656 37886 24712
rect 38106 24656 38162 24712
rect 38106 23296 38162 23352
rect 38106 21936 38162 21992
rect 38106 20576 38162 20632
rect 38106 19216 38162 19272
rect 38106 17856 38162 17912
rect 38106 16496 38162 16552
rect 38106 15136 38162 15192
rect 38290 13812 38292 13832
rect 38292 13812 38344 13832
rect 38344 13812 38346 13832
rect 38290 13776 38346 13812
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 38290 12416 38346 12472
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 38106 11056 38162 11112
rect 37830 10104 37886 10160
rect 37830 9832 37886 9888
rect 38106 9696 38162 9752
rect 38106 8336 38162 8392
rect 38106 6976 38162 7032
rect 38106 5616 38162 5672
rect 38106 4256 38162 4312
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 38106 2932 38108 2952
rect 38108 2932 38160 2952
rect 38160 2932 38162 2952
rect 38106 2896 38162 2932
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 38106 1536 38162 1592
<< metal3 >>
rect 36813 38314 36879 38317
rect 39200 38314 40000 38344
rect 36813 38312 40000 38314
rect 36813 38256 36818 38312
rect 36874 38256 40000 38312
rect 36813 38254 40000 38256
rect 36813 38251 36879 38254
rect 39200 38224 40000 38254
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 36721 36954 36787 36957
rect 39200 36954 40000 36984
rect 36721 36952 40000 36954
rect 36721 36896 36726 36952
rect 36782 36896 40000 36952
rect 36721 36894 40000 36896
rect 36721 36891 36787 36894
rect 39200 36864 40000 36894
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 38101 35594 38167 35597
rect 39200 35594 40000 35624
rect 38101 35592 40000 35594
rect 38101 35536 38106 35592
rect 38162 35536 40000 35592
rect 38101 35534 40000 35536
rect 38101 35531 38167 35534
rect 39200 35504 40000 35534
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 23974 35124 23980 35188
rect 24044 35186 24050 35188
rect 34789 35186 34855 35189
rect 24044 35184 34855 35186
rect 24044 35128 34794 35184
rect 34850 35128 34855 35184
rect 24044 35126 34855 35128
rect 24044 35124 24050 35126
rect 34789 35123 34855 35126
rect 19701 35050 19767 35053
rect 25037 35050 25103 35053
rect 30741 35052 30807 35053
rect 30741 35050 30788 35052
rect 19701 35048 25103 35050
rect 19701 34992 19706 35048
rect 19762 34992 25042 35048
rect 25098 34992 25103 35048
rect 19701 34990 25103 34992
rect 30696 35048 30788 35050
rect 30696 34992 30746 35048
rect 30696 34990 30788 34992
rect 19701 34987 19767 34990
rect 25037 34987 25103 34990
rect 30741 34988 30788 34990
rect 30852 34988 30858 35052
rect 30741 34987 30807 34988
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 28022 34580 28028 34644
rect 28092 34642 28098 34644
rect 28901 34642 28967 34645
rect 28092 34640 28967 34642
rect 28092 34584 28906 34640
rect 28962 34584 28967 34640
rect 28092 34582 28967 34584
rect 28092 34580 28098 34582
rect 28901 34579 28967 34582
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19517 34234 19583 34237
rect 23749 34234 23815 34237
rect 19517 34232 23815 34234
rect 19517 34176 19522 34232
rect 19578 34176 23754 34232
rect 23810 34176 23815 34232
rect 19517 34174 23815 34176
rect 19517 34171 19583 34174
rect 23749 34171 23815 34174
rect 38101 34234 38167 34237
rect 39200 34234 40000 34264
rect 38101 34232 40000 34234
rect 38101 34176 38106 34232
rect 38162 34176 40000 34232
rect 38101 34174 40000 34176
rect 38101 34171 38167 34174
rect 39200 34144 40000 34174
rect 16021 34098 16087 34101
rect 28758 34098 28764 34100
rect 16021 34096 28764 34098
rect 16021 34040 16026 34096
rect 16082 34040 28764 34096
rect 16021 34038 28764 34040
rect 16021 34035 16087 34038
rect 28758 34036 28764 34038
rect 28828 34098 28834 34100
rect 31385 34098 31451 34101
rect 28828 34096 31451 34098
rect 28828 34040 31390 34096
rect 31446 34040 31451 34096
rect 28828 34038 31451 34040
rect 28828 34036 28834 34038
rect 31385 34035 31451 34038
rect 5717 33962 5783 33965
rect 20662 33962 20668 33964
rect 5717 33960 20668 33962
rect 5717 33904 5722 33960
rect 5778 33904 20668 33960
rect 5717 33902 20668 33904
rect 5717 33899 5783 33902
rect 20662 33900 20668 33902
rect 20732 33900 20738 33964
rect 21817 33962 21883 33965
rect 22737 33962 22803 33965
rect 31293 33964 31359 33965
rect 31293 33962 31340 33964
rect 21817 33960 22803 33962
rect 21817 33904 21822 33960
rect 21878 33904 22742 33960
rect 22798 33904 22803 33960
rect 21817 33902 22803 33904
rect 31248 33960 31340 33962
rect 31248 33904 31298 33960
rect 31248 33902 31340 33904
rect 21817 33899 21883 33902
rect 22737 33899 22803 33902
rect 31293 33900 31340 33902
rect 31404 33900 31410 33964
rect 31293 33899 31359 33900
rect 30097 33828 30163 33829
rect 30046 33764 30052 33828
rect 30116 33826 30163 33828
rect 34421 33826 34487 33829
rect 30116 33824 34487 33826
rect 30158 33768 34426 33824
rect 34482 33768 34487 33824
rect 30116 33766 34487 33768
rect 30116 33764 30163 33766
rect 30097 33763 30163 33764
rect 34421 33763 34487 33766
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 34329 33554 34395 33557
rect 35893 33554 35959 33557
rect 34329 33552 35959 33554
rect 34329 33496 34334 33552
rect 34390 33496 35898 33552
rect 35954 33496 35959 33552
rect 34329 33494 35959 33496
rect 34329 33491 34395 33494
rect 35893 33491 35959 33494
rect 27470 33356 27476 33420
rect 27540 33418 27546 33420
rect 30741 33418 30807 33421
rect 27540 33416 30807 33418
rect 27540 33360 30746 33416
rect 30802 33360 30807 33416
rect 27540 33358 30807 33360
rect 27540 33356 27546 33358
rect 30741 33355 30807 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 30097 32874 30163 32877
rect 31937 32874 32003 32877
rect 32806 32874 32812 32876
rect 30097 32872 32812 32874
rect 30097 32816 30102 32872
rect 30158 32816 31942 32872
rect 31998 32816 32812 32872
rect 30097 32814 32812 32816
rect 30097 32811 30163 32814
rect 31937 32811 32003 32814
rect 32806 32812 32812 32814
rect 32876 32812 32882 32876
rect 38101 32874 38167 32877
rect 39200 32874 40000 32904
rect 38101 32872 40000 32874
rect 38101 32816 38106 32872
rect 38162 32816 40000 32872
rect 38101 32814 40000 32816
rect 38101 32811 38167 32814
rect 39200 32784 40000 32814
rect 20478 32676 20484 32740
rect 20548 32738 20554 32740
rect 20897 32738 20963 32741
rect 20548 32736 20963 32738
rect 20548 32680 20902 32736
rect 20958 32680 20963 32736
rect 20548 32678 20963 32680
rect 20548 32676 20554 32678
rect 20897 32675 20963 32678
rect 30097 32738 30163 32741
rect 31293 32738 31359 32741
rect 30097 32736 31359 32738
rect 30097 32680 30102 32736
rect 30158 32680 31298 32736
rect 31354 32680 31359 32736
rect 30097 32678 31359 32680
rect 30097 32675 30163 32678
rect 31293 32675 31359 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 12617 32466 12683 32469
rect 25221 32466 25287 32469
rect 12617 32464 25287 32466
rect 12617 32408 12622 32464
rect 12678 32408 25226 32464
rect 25282 32408 25287 32464
rect 12617 32406 25287 32408
rect 12617 32403 12683 32406
rect 25221 32403 25287 32406
rect 30598 32404 30604 32468
rect 30668 32466 30674 32468
rect 31661 32466 31727 32469
rect 30668 32464 31727 32466
rect 30668 32408 31666 32464
rect 31722 32408 31727 32464
rect 30668 32406 31727 32408
rect 30668 32404 30674 32406
rect 31661 32403 31727 32406
rect 9489 32330 9555 32333
rect 13537 32330 13603 32333
rect 9489 32328 13603 32330
rect 9489 32272 9494 32328
rect 9550 32272 13542 32328
rect 13598 32272 13603 32328
rect 9489 32270 13603 32272
rect 9489 32267 9555 32270
rect 13537 32267 13603 32270
rect 14365 32330 14431 32333
rect 17585 32330 17651 32333
rect 14365 32328 17651 32330
rect 14365 32272 14370 32328
rect 14426 32272 17590 32328
rect 17646 32272 17651 32328
rect 14365 32270 17651 32272
rect 14365 32267 14431 32270
rect 17585 32267 17651 32270
rect 21817 32330 21883 32333
rect 23105 32330 23171 32333
rect 21817 32328 23171 32330
rect 21817 32272 21822 32328
rect 21878 32272 23110 32328
rect 23166 32272 23171 32328
rect 21817 32270 23171 32272
rect 21817 32267 21883 32270
rect 23105 32267 23171 32270
rect 24025 32330 24091 32333
rect 26233 32330 26299 32333
rect 24025 32328 26299 32330
rect 24025 32272 24030 32328
rect 24086 32272 26238 32328
rect 26294 32272 26299 32328
rect 24025 32270 26299 32272
rect 24025 32267 24091 32270
rect 26233 32267 26299 32270
rect 17401 32194 17467 32197
rect 17677 32194 17743 32197
rect 17401 32192 17743 32194
rect 17401 32136 17406 32192
rect 17462 32136 17682 32192
rect 17738 32136 17743 32192
rect 17401 32134 17743 32136
rect 17401 32131 17467 32134
rect 17677 32131 17743 32134
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 12157 31922 12223 31925
rect 12341 31922 12407 31925
rect 12157 31920 12407 31922
rect 12157 31864 12162 31920
rect 12218 31864 12346 31920
rect 12402 31864 12407 31920
rect 12157 31862 12407 31864
rect 12157 31859 12223 31862
rect 12341 31859 12407 31862
rect 5165 31786 5231 31789
rect 9213 31786 9279 31789
rect 10409 31786 10475 31789
rect 5165 31784 10475 31786
rect 5165 31728 5170 31784
rect 5226 31728 9218 31784
rect 9274 31728 10414 31784
rect 10470 31728 10475 31784
rect 5165 31726 10475 31728
rect 5165 31723 5231 31726
rect 9213 31723 9279 31726
rect 10409 31723 10475 31726
rect 11605 31786 11671 31789
rect 12157 31786 12223 31789
rect 11605 31784 12223 31786
rect 11605 31728 11610 31784
rect 11666 31728 12162 31784
rect 12218 31728 12223 31784
rect 11605 31726 12223 31728
rect 11605 31723 11671 31726
rect 12157 31723 12223 31726
rect 17166 31724 17172 31788
rect 17236 31786 17242 31788
rect 17309 31786 17375 31789
rect 17236 31784 17375 31786
rect 17236 31728 17314 31784
rect 17370 31728 17375 31784
rect 17236 31726 17375 31728
rect 17236 31724 17242 31726
rect 17309 31723 17375 31726
rect 19701 31786 19767 31789
rect 25681 31786 25747 31789
rect 28901 31786 28967 31789
rect 19701 31784 20040 31786
rect 19701 31728 19706 31784
rect 19762 31728 20040 31784
rect 19701 31726 20040 31728
rect 19701 31723 19767 31726
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 19980 31106 20040 31726
rect 25681 31784 28967 31786
rect 25681 31728 25686 31784
rect 25742 31728 28906 31784
rect 28962 31728 28967 31784
rect 25681 31726 28967 31728
rect 25681 31723 25747 31726
rect 28901 31723 28967 31726
rect 38101 31514 38167 31517
rect 39200 31514 40000 31544
rect 38101 31512 40000 31514
rect 38101 31456 38106 31512
rect 38162 31456 40000 31512
rect 38101 31454 40000 31456
rect 38101 31451 38167 31454
rect 39200 31424 40000 31454
rect 31753 31378 31819 31381
rect 34605 31378 34671 31381
rect 34789 31378 34855 31381
rect 31753 31376 34855 31378
rect 31753 31320 31758 31376
rect 31814 31320 34610 31376
rect 34666 31320 34794 31376
rect 34850 31320 34855 31376
rect 31753 31318 34855 31320
rect 31753 31315 31819 31318
rect 34605 31315 34671 31318
rect 34789 31315 34855 31318
rect 25814 31180 25820 31244
rect 25884 31242 25890 31244
rect 30741 31242 30807 31245
rect 25884 31240 30807 31242
rect 25884 31184 30746 31240
rect 30802 31184 30807 31240
rect 25884 31182 30807 31184
rect 25884 31180 25890 31182
rect 30741 31179 30807 31182
rect 20161 31106 20227 31109
rect 19980 31104 20227 31106
rect 19980 31048 20166 31104
rect 20222 31048 20227 31104
rect 19980 31046 20227 31048
rect 20161 31043 20227 31046
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19885 30970 19951 30973
rect 20478 30970 20484 30972
rect 19885 30968 20484 30970
rect 19885 30912 19890 30968
rect 19946 30912 20484 30968
rect 19885 30910 20484 30912
rect 19885 30907 19951 30910
rect 20478 30908 20484 30910
rect 20548 30908 20554 30972
rect 20662 30908 20668 30972
rect 20732 30970 20738 30972
rect 30465 30970 30531 30973
rect 20732 30968 30531 30970
rect 20732 30912 30470 30968
rect 30526 30912 30531 30968
rect 20732 30910 30531 30912
rect 20732 30908 20738 30910
rect 30465 30907 30531 30910
rect 19701 30834 19767 30837
rect 20805 30834 20871 30837
rect 19701 30832 20871 30834
rect 19701 30776 19706 30832
rect 19762 30776 20810 30832
rect 20866 30776 20871 30832
rect 19701 30774 20871 30776
rect 19701 30771 19767 30774
rect 20805 30771 20871 30774
rect 24853 30834 24919 30837
rect 26417 30834 26483 30837
rect 24853 30832 26483 30834
rect 24853 30776 24858 30832
rect 24914 30776 26422 30832
rect 26478 30776 26483 30832
rect 24853 30774 26483 30776
rect 24853 30771 24919 30774
rect 26417 30771 26483 30774
rect 13721 30698 13787 30701
rect 20110 30698 20116 30700
rect 13721 30696 20116 30698
rect 13721 30640 13726 30696
rect 13782 30640 20116 30696
rect 13721 30638 20116 30640
rect 13721 30635 13787 30638
rect 20110 30636 20116 30638
rect 20180 30636 20186 30700
rect 20529 30698 20595 30701
rect 22369 30698 22435 30701
rect 20529 30696 22435 30698
rect 20529 30640 20534 30696
rect 20590 30640 22374 30696
rect 22430 30640 22435 30696
rect 20529 30638 22435 30640
rect 20529 30635 20595 30638
rect 22369 30635 22435 30638
rect 23381 30698 23447 30701
rect 27705 30698 27771 30701
rect 35525 30700 35591 30701
rect 35525 30698 35572 30700
rect 23381 30696 27771 30698
rect 23381 30640 23386 30696
rect 23442 30640 27710 30696
rect 27766 30640 27771 30696
rect 23381 30638 27771 30640
rect 35480 30696 35572 30698
rect 35480 30640 35530 30696
rect 35480 30638 35572 30640
rect 23381 30635 23447 30638
rect 27705 30635 27771 30638
rect 35525 30636 35572 30638
rect 35636 30636 35642 30700
rect 35525 30635 35591 30636
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 14549 30290 14615 30293
rect 27705 30290 27771 30293
rect 28022 30290 28028 30292
rect 14549 30288 28028 30290
rect 14549 30232 14554 30288
rect 14610 30232 27710 30288
rect 27766 30232 28028 30288
rect 14549 30230 28028 30232
rect 14549 30227 14615 30230
rect 27705 30227 27771 30230
rect 28022 30228 28028 30230
rect 28092 30228 28098 30292
rect 31017 30290 31083 30293
rect 35893 30290 35959 30293
rect 37825 30290 37891 30293
rect 31017 30288 37891 30290
rect 31017 30232 31022 30288
rect 31078 30232 35898 30288
rect 35954 30232 37830 30288
rect 37886 30232 37891 30288
rect 31017 30230 37891 30232
rect 31017 30227 31083 30230
rect 35893 30227 35959 30230
rect 37825 30227 37891 30230
rect 36997 30154 37063 30157
rect 39200 30154 40000 30184
rect 36997 30152 40000 30154
rect 36997 30096 37002 30152
rect 37058 30096 40000 30152
rect 36997 30094 40000 30096
rect 36997 30091 37063 30094
rect 39200 30064 40000 30094
rect 30230 29956 30236 30020
rect 30300 30018 30306 30020
rect 30373 30018 30439 30021
rect 30300 30016 30439 30018
rect 30300 29960 30378 30016
rect 30434 29960 30439 30016
rect 30300 29958 30439 29960
rect 30300 29956 30306 29958
rect 30373 29955 30439 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 25497 29882 25563 29885
rect 26509 29882 26575 29885
rect 25497 29880 26575 29882
rect 25497 29824 25502 29880
rect 25558 29824 26514 29880
rect 26570 29824 26575 29880
rect 25497 29822 26575 29824
rect 25497 29819 25563 29822
rect 26509 29819 26575 29822
rect 31017 29746 31083 29749
rect 31150 29746 31156 29748
rect 31017 29744 31156 29746
rect 31017 29688 31022 29744
rect 31078 29688 31156 29744
rect 31017 29686 31156 29688
rect 31017 29683 31083 29686
rect 31150 29684 31156 29686
rect 31220 29684 31226 29748
rect 34881 29746 34947 29749
rect 35433 29746 35499 29749
rect 34881 29744 35499 29746
rect 34881 29688 34886 29744
rect 34942 29688 35438 29744
rect 35494 29688 35499 29744
rect 34881 29686 35499 29688
rect 34881 29683 34947 29686
rect 35433 29683 35499 29686
rect 15745 29610 15811 29613
rect 16665 29610 16731 29613
rect 15745 29608 16731 29610
rect 15745 29552 15750 29608
rect 15806 29552 16670 29608
rect 16726 29552 16731 29608
rect 15745 29550 16731 29552
rect 15745 29547 15811 29550
rect 16665 29547 16731 29550
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 24301 29338 24367 29341
rect 25221 29338 25287 29341
rect 24301 29336 25287 29338
rect 24301 29280 24306 29336
rect 24362 29280 25226 29336
rect 25282 29280 25287 29336
rect 24301 29278 25287 29280
rect 24301 29275 24367 29278
rect 25221 29275 25287 29278
rect 19425 29202 19491 29205
rect 25129 29202 25195 29205
rect 19425 29200 25195 29202
rect 19425 29144 19430 29200
rect 19486 29144 25134 29200
rect 25190 29144 25195 29200
rect 19425 29142 25195 29144
rect 19425 29139 19491 29142
rect 25129 29139 25195 29142
rect 29361 29202 29427 29205
rect 30373 29202 30439 29205
rect 29361 29200 30439 29202
rect 29361 29144 29366 29200
rect 29422 29144 30378 29200
rect 30434 29144 30439 29200
rect 29361 29142 30439 29144
rect 29361 29139 29427 29142
rect 30373 29139 30439 29142
rect 17401 29066 17467 29069
rect 17401 29064 19994 29066
rect 17401 29008 17406 29064
rect 17462 29008 19994 29064
rect 17401 29006 19994 29008
rect 17401 29003 17467 29006
rect 19934 28933 19994 29006
rect 20110 29004 20116 29068
rect 20180 29066 20186 29068
rect 20253 29066 20319 29069
rect 20180 29064 20319 29066
rect 20180 29008 20258 29064
rect 20314 29008 20319 29064
rect 20180 29006 20319 29008
rect 20180 29004 20186 29006
rect 20253 29003 20319 29006
rect 21909 29066 21975 29069
rect 27613 29066 27679 29069
rect 29545 29068 29611 29069
rect 29494 29066 29500 29068
rect 21909 29064 27679 29066
rect 21909 29008 21914 29064
rect 21970 29008 27618 29064
rect 27674 29008 27679 29064
rect 21909 29006 27679 29008
rect 29454 29006 29500 29066
rect 29564 29064 29611 29068
rect 29606 29008 29611 29064
rect 21909 29003 21975 29006
rect 27613 29003 27679 29006
rect 29494 29004 29500 29006
rect 29564 29004 29611 29008
rect 29545 29003 29611 29004
rect 19934 28928 20043 28933
rect 19934 28872 19982 28928
rect 20038 28872 20043 28928
rect 19934 28870 20043 28872
rect 19977 28867 20043 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 37733 28794 37799 28797
rect 39200 28794 40000 28824
rect 37733 28792 40000 28794
rect 37733 28736 37738 28792
rect 37794 28736 40000 28792
rect 37733 28734 40000 28736
rect 37733 28731 37799 28734
rect 39200 28704 40000 28734
rect 4061 28522 4127 28525
rect 5441 28522 5507 28525
rect 5809 28522 5875 28525
rect 8477 28522 8543 28525
rect 4061 28520 8543 28522
rect 4061 28464 4066 28520
rect 4122 28464 5446 28520
rect 5502 28464 5814 28520
rect 5870 28464 8482 28520
rect 8538 28464 8543 28520
rect 4061 28462 8543 28464
rect 4061 28459 4127 28462
rect 5441 28459 5507 28462
rect 5809 28459 5875 28462
rect 8477 28459 8543 28462
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 19977 28114 20043 28117
rect 22686 28114 22692 28116
rect 19977 28112 22692 28114
rect 19977 28056 19982 28112
rect 20038 28056 22692 28112
rect 19977 28054 22692 28056
rect 19977 28051 20043 28054
rect 22686 28052 22692 28054
rect 22756 28114 22762 28116
rect 23289 28114 23355 28117
rect 22756 28112 23355 28114
rect 22756 28056 23294 28112
rect 23350 28056 23355 28112
rect 22756 28054 23355 28056
rect 22756 28052 22762 28054
rect 23289 28051 23355 28054
rect 27286 27780 27292 27844
rect 27356 27842 27362 27844
rect 28717 27842 28783 27845
rect 27356 27840 28783 27842
rect 27356 27784 28722 27840
rect 28778 27784 28783 27840
rect 27356 27782 28783 27784
rect 27356 27780 27362 27782
rect 28717 27779 28783 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 25998 27644 26004 27708
rect 26068 27706 26074 27708
rect 27613 27706 27679 27709
rect 26068 27704 27679 27706
rect 26068 27648 27618 27704
rect 27674 27648 27679 27704
rect 26068 27646 27679 27648
rect 26068 27644 26074 27646
rect 27613 27643 27679 27646
rect 28390 27644 28396 27708
rect 28460 27706 28466 27708
rect 28809 27706 28875 27709
rect 28460 27704 28875 27706
rect 28460 27648 28814 27704
rect 28870 27648 28875 27704
rect 28460 27646 28875 27648
rect 28460 27644 28466 27646
rect 28809 27643 28875 27646
rect 9581 27434 9647 27437
rect 13721 27434 13787 27437
rect 9581 27432 13787 27434
rect 9581 27376 9586 27432
rect 9642 27376 13726 27432
rect 13782 27376 13787 27432
rect 9581 27374 13787 27376
rect 9581 27371 9647 27374
rect 13721 27371 13787 27374
rect 19977 27434 20043 27437
rect 23473 27434 23539 27437
rect 24945 27434 25011 27437
rect 19977 27432 25011 27434
rect 19977 27376 19982 27432
rect 20038 27376 23478 27432
rect 23534 27376 24950 27432
rect 25006 27376 25011 27432
rect 19977 27374 25011 27376
rect 19977 27371 20043 27374
rect 23473 27371 23539 27374
rect 24945 27371 25011 27374
rect 37181 27434 37247 27437
rect 39200 27434 40000 27464
rect 37181 27432 40000 27434
rect 37181 27376 37186 27432
rect 37242 27376 40000 27432
rect 37181 27374 40000 27376
rect 37181 27371 37247 27374
rect 39200 27344 40000 27374
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4797 27162 4863 27165
rect 5165 27162 5231 27165
rect 4797 27160 5231 27162
rect 4797 27104 4802 27160
rect 4858 27104 5170 27160
rect 5226 27104 5231 27160
rect 4797 27102 5231 27104
rect 4797 27099 4863 27102
rect 5165 27099 5231 27102
rect 23013 27162 23079 27165
rect 23381 27162 23447 27165
rect 23013 27160 23447 27162
rect 23013 27104 23018 27160
rect 23074 27104 23386 27160
rect 23442 27104 23447 27160
rect 23013 27102 23447 27104
rect 23013 27099 23079 27102
rect 23381 27099 23447 27102
rect 30097 27026 30163 27029
rect 31753 27026 31819 27029
rect 30097 27024 31819 27026
rect 30097 26968 30102 27024
rect 30158 26968 31758 27024
rect 31814 26968 31819 27024
rect 30097 26966 31819 26968
rect 30097 26963 30163 26966
rect 31753 26963 31819 26966
rect 20161 26890 20227 26893
rect 21173 26890 21239 26893
rect 25129 26890 25195 26893
rect 20161 26888 25195 26890
rect 20161 26832 20166 26888
rect 20222 26832 21178 26888
rect 21234 26832 25134 26888
rect 25190 26832 25195 26888
rect 20161 26830 25195 26832
rect 20161 26827 20227 26830
rect 21173 26827 21239 26830
rect 25129 26827 25195 26830
rect 27521 26890 27587 26893
rect 30189 26890 30255 26893
rect 27521 26888 30255 26890
rect 27521 26832 27526 26888
rect 27582 26832 30194 26888
rect 30250 26832 30255 26888
rect 27521 26830 30255 26832
rect 27521 26827 27587 26830
rect 30189 26827 30255 26830
rect 32121 26890 32187 26893
rect 37273 26890 37339 26893
rect 32121 26888 37339 26890
rect 32121 26832 32126 26888
rect 32182 26832 37278 26888
rect 37334 26832 37339 26888
rect 32121 26830 37339 26832
rect 32121 26827 32187 26830
rect 37273 26827 37339 26830
rect 8886 26692 8892 26756
rect 8956 26754 8962 26756
rect 9213 26754 9279 26757
rect 8956 26752 9279 26754
rect 8956 26696 9218 26752
rect 9274 26696 9279 26752
rect 8956 26694 9279 26696
rect 8956 26692 8962 26694
rect 9213 26691 9279 26694
rect 22369 26754 22435 26757
rect 23289 26754 23355 26757
rect 34605 26756 34671 26757
rect 34605 26754 34652 26756
rect 22369 26752 23355 26754
rect 22369 26696 22374 26752
rect 22430 26696 23294 26752
rect 23350 26696 23355 26752
rect 22369 26694 23355 26696
rect 34560 26752 34652 26754
rect 34560 26696 34610 26752
rect 34560 26694 34652 26696
rect 22369 26691 22435 26694
rect 23289 26691 23355 26694
rect 34605 26692 34652 26694
rect 34716 26692 34722 26756
rect 34605 26691 34671 26692
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 5993 26482 6059 26485
rect 9489 26482 9555 26485
rect 5993 26480 9555 26482
rect 5993 26424 5998 26480
rect 6054 26424 9494 26480
rect 9550 26424 9555 26480
rect 5993 26422 9555 26424
rect 5993 26419 6059 26422
rect 9489 26419 9555 26422
rect 20989 26482 21055 26485
rect 25773 26482 25839 26485
rect 20989 26480 25839 26482
rect 20989 26424 20994 26480
rect 21050 26424 25778 26480
rect 25834 26424 25839 26480
rect 20989 26422 25839 26424
rect 20989 26419 21055 26422
rect 25773 26419 25839 26422
rect 32397 26482 32463 26485
rect 38009 26482 38075 26485
rect 32397 26480 38075 26482
rect 32397 26424 32402 26480
rect 32458 26424 38014 26480
rect 38070 26424 38075 26480
rect 32397 26422 38075 26424
rect 32397 26419 32463 26422
rect 38009 26419 38075 26422
rect 19333 26346 19399 26349
rect 23657 26346 23723 26349
rect 19333 26344 23723 26346
rect 19333 26288 19338 26344
rect 19394 26288 23662 26344
rect 23718 26288 23723 26344
rect 19333 26286 23723 26288
rect 19333 26283 19399 26286
rect 23657 26283 23723 26286
rect 29729 26346 29795 26349
rect 29862 26346 29868 26348
rect 29729 26344 29868 26346
rect 29729 26288 29734 26344
rect 29790 26288 29868 26344
rect 29729 26286 29868 26288
rect 29729 26283 29795 26286
rect 29862 26284 29868 26286
rect 29932 26284 29938 26348
rect 34646 26346 34652 26348
rect 31710 26286 34652 26346
rect 27613 26210 27679 26213
rect 28257 26210 28323 26213
rect 27613 26208 28323 26210
rect 27613 26152 27618 26208
rect 27674 26152 28262 26208
rect 28318 26152 28323 26208
rect 27613 26150 28323 26152
rect 27613 26147 27679 26150
rect 28257 26147 28323 26150
rect 31150 26148 31156 26212
rect 31220 26210 31226 26212
rect 31710 26210 31770 26286
rect 34646 26284 34652 26286
rect 34716 26284 34722 26348
rect 31220 26150 31770 26210
rect 31220 26148 31226 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 27838 26012 27844 26076
rect 27908 26074 27914 26076
rect 27981 26074 28047 26077
rect 31158 26074 31218 26148
rect 27908 26072 31218 26074
rect 27908 26016 27986 26072
rect 28042 26016 31218 26072
rect 27908 26014 31218 26016
rect 38101 26074 38167 26077
rect 39200 26074 40000 26104
rect 38101 26072 40000 26074
rect 38101 26016 38106 26072
rect 38162 26016 40000 26072
rect 38101 26014 40000 26016
rect 27908 26012 27914 26014
rect 27981 26011 28047 26014
rect 38101 26011 38167 26014
rect 39200 25984 40000 26014
rect 17166 25876 17172 25940
rect 17236 25938 17242 25940
rect 21173 25938 21239 25941
rect 17236 25936 21239 25938
rect 17236 25880 21178 25936
rect 21234 25880 21239 25936
rect 17236 25878 21239 25880
rect 17236 25876 17242 25878
rect 21173 25875 21239 25878
rect 24485 25938 24551 25941
rect 25957 25938 26023 25941
rect 24485 25936 26023 25938
rect 24485 25880 24490 25936
rect 24546 25880 25962 25936
rect 26018 25880 26023 25936
rect 24485 25878 26023 25880
rect 24485 25875 24551 25878
rect 25957 25875 26023 25878
rect 21541 25802 21607 25805
rect 24853 25802 24919 25805
rect 21541 25800 24919 25802
rect 21541 25744 21546 25800
rect 21602 25744 24858 25800
rect 24914 25744 24919 25800
rect 21541 25742 24919 25744
rect 21541 25739 21607 25742
rect 24853 25739 24919 25742
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 15101 25530 15167 25533
rect 24669 25530 24735 25533
rect 15101 25528 24735 25530
rect 15101 25472 15106 25528
rect 15162 25472 24674 25528
rect 24730 25472 24735 25528
rect 15101 25470 24735 25472
rect 15101 25467 15167 25470
rect 24669 25467 24735 25470
rect 21909 25122 21975 25125
rect 29085 25122 29151 25125
rect 21909 25120 29151 25122
rect 21909 25064 21914 25120
rect 21970 25064 29090 25120
rect 29146 25064 29151 25120
rect 21909 25062 29151 25064
rect 21909 25059 21975 25062
rect 29085 25059 29151 25062
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 28257 24986 28323 24989
rect 28574 24986 28580 24988
rect 28257 24984 28580 24986
rect 28257 24928 28262 24984
rect 28318 24928 28580 24984
rect 28257 24926 28580 24928
rect 28257 24923 28323 24926
rect 28574 24924 28580 24926
rect 28644 24924 28650 24988
rect 27429 24852 27495 24853
rect 27429 24848 27476 24852
rect 27540 24850 27546 24852
rect 31753 24850 31819 24853
rect 32673 24850 32739 24853
rect 32806 24850 32812 24852
rect 27429 24792 27434 24848
rect 27429 24788 27476 24792
rect 27540 24790 27586 24850
rect 31753 24848 32812 24850
rect 31753 24792 31758 24848
rect 31814 24792 32678 24848
rect 32734 24792 32812 24848
rect 31753 24790 32812 24792
rect 27540 24788 27546 24790
rect 27429 24787 27495 24788
rect 31753 24787 31819 24790
rect 32673 24787 32739 24790
rect 32806 24788 32812 24790
rect 32876 24788 32882 24852
rect 22737 24716 22803 24717
rect 22686 24652 22692 24716
rect 22756 24714 22803 24716
rect 23749 24714 23815 24717
rect 28022 24714 28028 24716
rect 22756 24712 22848 24714
rect 22798 24656 22848 24712
rect 22756 24654 22848 24656
rect 23749 24712 28028 24714
rect 23749 24656 23754 24712
rect 23810 24656 28028 24712
rect 23749 24654 28028 24656
rect 22756 24652 22803 24654
rect 22737 24651 22803 24652
rect 23749 24651 23815 24654
rect 28022 24652 28028 24654
rect 28092 24652 28098 24716
rect 32397 24714 32463 24717
rect 37825 24714 37891 24717
rect 32397 24712 37891 24714
rect 32397 24656 32402 24712
rect 32458 24656 37830 24712
rect 37886 24656 37891 24712
rect 32397 24654 37891 24656
rect 32397 24651 32463 24654
rect 37825 24651 37891 24654
rect 38101 24714 38167 24717
rect 39200 24714 40000 24744
rect 38101 24712 40000 24714
rect 38101 24656 38106 24712
rect 38162 24656 40000 24712
rect 38101 24654 40000 24656
rect 38101 24651 38167 24654
rect 39200 24624 40000 24654
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 22737 24442 22803 24445
rect 25681 24442 25747 24445
rect 22737 24440 25747 24442
rect 22737 24384 22742 24440
rect 22798 24384 25686 24440
rect 25742 24384 25747 24440
rect 22737 24382 25747 24384
rect 22737 24379 22803 24382
rect 25681 24379 25747 24382
rect 21081 24170 21147 24173
rect 26509 24170 26575 24173
rect 21081 24168 26575 24170
rect 21081 24112 21086 24168
rect 21142 24112 26514 24168
rect 26570 24112 26575 24168
rect 21081 24110 26575 24112
rect 21081 24107 21147 24110
rect 26509 24107 26575 24110
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 28717 23764 28783 23765
rect 28717 23762 28764 23764
rect 23292 23760 28764 23762
rect 28828 23762 28834 23764
rect 31017 23762 31083 23765
rect 28828 23760 31083 23762
rect 23292 23704 28722 23760
rect 28828 23704 31022 23760
rect 31078 23704 31083 23760
rect 23292 23702 28764 23704
rect 23292 23493 23352 23702
rect 28717 23700 28764 23702
rect 28828 23702 31083 23704
rect 28828 23700 28834 23702
rect 28717 23699 28783 23700
rect 31017 23699 31083 23702
rect 26918 23564 26924 23628
rect 26988 23626 26994 23628
rect 27337 23626 27403 23629
rect 26988 23624 30298 23626
rect 26988 23568 27342 23624
rect 27398 23568 30298 23624
rect 26988 23566 30298 23568
rect 26988 23564 26994 23566
rect 27337 23563 27403 23566
rect 30238 23493 30298 23566
rect 23289 23488 23355 23493
rect 23289 23432 23294 23488
rect 23350 23432 23355 23488
rect 23289 23427 23355 23432
rect 30238 23490 30347 23493
rect 30598 23490 30604 23492
rect 30238 23488 30604 23490
rect 30238 23432 30286 23488
rect 30342 23432 30604 23488
rect 30238 23430 30604 23432
rect 30281 23427 30347 23430
rect 30598 23428 30604 23430
rect 30668 23428 30674 23492
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 28625 23354 28691 23357
rect 30046 23354 30052 23356
rect 28625 23352 30052 23354
rect 28625 23296 28630 23352
rect 28686 23296 30052 23352
rect 28625 23294 30052 23296
rect 28625 23291 28691 23294
rect 30046 23292 30052 23294
rect 30116 23354 30122 23356
rect 33317 23354 33383 23357
rect 30116 23352 33383 23354
rect 30116 23296 33322 23352
rect 33378 23296 33383 23352
rect 30116 23294 33383 23296
rect 30116 23292 30122 23294
rect 33317 23291 33383 23294
rect 38101 23354 38167 23357
rect 39200 23354 40000 23384
rect 38101 23352 40000 23354
rect 38101 23296 38106 23352
rect 38162 23296 40000 23352
rect 38101 23294 40000 23296
rect 38101 23291 38167 23294
rect 20713 23218 20779 23221
rect 26785 23218 26851 23221
rect 28257 23218 28323 23221
rect 20713 23216 28323 23218
rect 20713 23160 20718 23216
rect 20774 23160 26790 23216
rect 26846 23160 28262 23216
rect 28318 23160 28323 23216
rect 20713 23158 28323 23160
rect 33320 23218 33380 23291
rect 39200 23264 40000 23294
rect 35525 23218 35591 23221
rect 33320 23216 35591 23218
rect 33320 23160 35530 23216
rect 35586 23160 35591 23216
rect 33320 23158 35591 23160
rect 20713 23155 20779 23158
rect 26785 23155 26851 23158
rect 28257 23155 28323 23158
rect 35525 23155 35591 23158
rect 27705 23082 27771 23085
rect 30046 23082 30052 23084
rect 27705 23080 30052 23082
rect 27705 23024 27710 23080
rect 27766 23024 30052 23080
rect 27705 23022 30052 23024
rect 27705 23019 27771 23022
rect 30046 23020 30052 23022
rect 30116 23082 30122 23084
rect 34513 23082 34579 23085
rect 30116 23080 34579 23082
rect 30116 23024 34518 23080
rect 34574 23024 34579 23080
rect 30116 23022 34579 23024
rect 30116 23020 30122 23022
rect 34513 23019 34579 23022
rect 21633 22946 21699 22949
rect 26969 22946 27035 22949
rect 21633 22944 27035 22946
rect 21633 22888 21638 22944
rect 21694 22888 26974 22944
rect 27030 22888 27035 22944
rect 21633 22886 27035 22888
rect 21633 22883 21699 22886
rect 26969 22883 27035 22886
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 9857 22674 9923 22677
rect 11789 22674 11855 22677
rect 17217 22674 17283 22677
rect 9857 22672 17283 22674
rect 9857 22616 9862 22672
rect 9918 22616 11794 22672
rect 11850 22616 17222 22672
rect 17278 22616 17283 22672
rect 9857 22614 17283 22616
rect 9857 22611 9923 22614
rect 11789 22611 11855 22614
rect 17217 22611 17283 22614
rect 23473 22674 23539 22677
rect 28257 22674 28323 22677
rect 23473 22672 28323 22674
rect 23473 22616 23478 22672
rect 23534 22616 28262 22672
rect 28318 22616 28323 22672
rect 23473 22614 28323 22616
rect 23473 22611 23539 22614
rect 28257 22611 28323 22614
rect 29361 22674 29427 22677
rect 29494 22674 29500 22676
rect 29361 22672 29500 22674
rect 29361 22616 29366 22672
rect 29422 22616 29500 22672
rect 29361 22614 29500 22616
rect 29361 22611 29427 22614
rect 29494 22612 29500 22614
rect 29564 22612 29570 22676
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 28206 22204 28212 22268
rect 28276 22266 28282 22268
rect 28809 22266 28875 22269
rect 28276 22264 28875 22266
rect 28276 22208 28814 22264
rect 28870 22208 28875 22264
rect 28276 22206 28875 22208
rect 28276 22204 28282 22206
rect 28809 22203 28875 22206
rect 20529 21994 20595 21997
rect 23974 21994 23980 21996
rect 20529 21992 23980 21994
rect 20529 21936 20534 21992
rect 20590 21936 23980 21992
rect 20529 21934 23980 21936
rect 20529 21931 20595 21934
rect 23974 21932 23980 21934
rect 24044 21932 24050 21996
rect 26785 21994 26851 21997
rect 30782 21994 30788 21996
rect 26785 21992 30788 21994
rect 26785 21936 26790 21992
rect 26846 21936 30788 21992
rect 26785 21934 30788 21936
rect 26785 21931 26851 21934
rect 30782 21932 30788 21934
rect 30852 21932 30858 21996
rect 38101 21994 38167 21997
rect 39200 21994 40000 22024
rect 38101 21992 40000 21994
rect 38101 21936 38106 21992
rect 38162 21936 40000 21992
rect 38101 21934 40000 21936
rect 38101 21931 38167 21934
rect 39200 21904 40000 21934
rect 28533 21858 28599 21861
rect 31334 21858 31340 21860
rect 28533 21856 31340 21858
rect 28533 21800 28538 21856
rect 28594 21800 31340 21856
rect 28533 21798 31340 21800
rect 28533 21795 28599 21798
rect 31334 21796 31340 21798
rect 31404 21796 31410 21860
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 22829 21722 22895 21725
rect 29361 21722 29427 21725
rect 22829 21720 29427 21722
rect 22829 21664 22834 21720
rect 22890 21664 29366 21720
rect 29422 21664 29427 21720
rect 22829 21662 29427 21664
rect 22829 21659 22895 21662
rect 29361 21659 29427 21662
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 27061 20772 27127 20773
rect 27061 20768 27108 20772
rect 27172 20770 27178 20772
rect 27061 20712 27066 20768
rect 27061 20708 27108 20712
rect 27172 20710 27218 20770
rect 27172 20708 27178 20710
rect 27061 20707 27127 20708
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 25814 20572 25820 20636
rect 25884 20634 25890 20636
rect 26049 20634 26115 20637
rect 25884 20632 26115 20634
rect 25884 20576 26054 20632
rect 26110 20576 26115 20632
rect 25884 20574 26115 20576
rect 25884 20572 25890 20574
rect 26049 20571 26115 20574
rect 38101 20634 38167 20637
rect 39200 20634 40000 20664
rect 38101 20632 40000 20634
rect 38101 20576 38106 20632
rect 38162 20576 40000 20632
rect 38101 20574 40000 20576
rect 38101 20571 38167 20574
rect 39200 20544 40000 20574
rect 19425 20498 19491 20501
rect 29637 20498 29703 20501
rect 19425 20496 29703 20498
rect 19425 20440 19430 20496
rect 19486 20440 29642 20496
rect 29698 20440 29703 20496
rect 19425 20438 29703 20440
rect 19425 20435 19491 20438
rect 29637 20435 29703 20438
rect 10409 20362 10475 20365
rect 15745 20362 15811 20365
rect 10409 20360 15811 20362
rect 10409 20304 10414 20360
rect 10470 20304 15750 20360
rect 15806 20304 15811 20360
rect 10409 20302 15811 20304
rect 10409 20299 10475 20302
rect 15745 20299 15811 20302
rect 21357 20362 21423 20365
rect 24025 20362 24091 20365
rect 28257 20362 28323 20365
rect 21357 20360 28323 20362
rect 21357 20304 21362 20360
rect 21418 20304 24030 20360
rect 24086 20304 28262 20360
rect 28318 20304 28323 20360
rect 21357 20302 28323 20304
rect 21357 20299 21423 20302
rect 24025 20299 24091 20302
rect 28257 20299 28323 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 20529 20090 20595 20093
rect 25221 20090 25287 20093
rect 25681 20090 25747 20093
rect 20529 20088 25747 20090
rect 20529 20032 20534 20088
rect 20590 20032 25226 20088
rect 25282 20032 25686 20088
rect 25742 20032 25747 20088
rect 20529 20030 25747 20032
rect 20529 20027 20595 20030
rect 25221 20027 25287 20030
rect 25681 20027 25747 20030
rect 21909 19818 21975 19821
rect 23933 19818 23999 19821
rect 21909 19816 23999 19818
rect 21909 19760 21914 19816
rect 21970 19760 23938 19816
rect 23994 19760 23999 19816
rect 21909 19758 23999 19760
rect 21909 19755 21975 19758
rect 23933 19755 23999 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 24301 19410 24367 19413
rect 26233 19410 26299 19413
rect 27061 19410 27127 19413
rect 24301 19408 27127 19410
rect 24301 19352 24306 19408
rect 24362 19352 26238 19408
rect 26294 19352 27066 19408
rect 27122 19352 27127 19408
rect 32673 19410 32739 19413
rect 33317 19410 33383 19413
rect 32673 19408 33383 19410
rect 24301 19350 27127 19352
rect 28993 19350 29059 19353
rect 24301 19347 24367 19350
rect 26233 19347 26299 19350
rect 27061 19347 27127 19350
rect 28950 19348 29059 19350
rect 28950 19292 28998 19348
rect 29054 19292 29059 19348
rect 32673 19352 32678 19408
rect 32734 19352 33322 19408
rect 33378 19352 33383 19408
rect 32673 19350 33383 19352
rect 32673 19347 32739 19350
rect 33317 19347 33383 19350
rect 28950 19287 29059 19292
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 28950 19005 29010 19287
rect 38101 19274 38167 19277
rect 39200 19274 40000 19304
rect 38101 19272 40000 19274
rect 38101 19216 38106 19272
rect 38162 19216 40000 19272
rect 38101 19214 40000 19216
rect 38101 19211 38167 19214
rect 39200 19184 40000 19214
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 28950 19000 29059 19005
rect 28950 18944 28998 19000
rect 29054 18944 29059 19000
rect 28950 18942 29059 18944
rect 28993 18939 29059 18942
rect 21909 18866 21975 18869
rect 26918 18866 26924 18868
rect 21909 18864 26924 18866
rect 21909 18808 21914 18864
rect 21970 18808 26924 18864
rect 21909 18806 26924 18808
rect 21909 18803 21975 18806
rect 26918 18804 26924 18806
rect 26988 18804 26994 18868
rect 35157 18866 35223 18869
rect 35566 18866 35572 18868
rect 35157 18864 35572 18866
rect 35157 18808 35162 18864
rect 35218 18808 35572 18864
rect 35157 18806 35572 18808
rect 35157 18803 35223 18806
rect 35566 18804 35572 18806
rect 35636 18804 35642 18868
rect 30230 18668 30236 18732
rect 30300 18730 30306 18732
rect 33317 18730 33383 18733
rect 30300 18728 33383 18730
rect 30300 18672 33322 18728
rect 33378 18672 33383 18728
rect 30300 18670 33383 18672
rect 30300 18668 30306 18670
rect 33317 18667 33383 18670
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 20069 18458 20135 18461
rect 22553 18458 22619 18461
rect 20069 18456 22619 18458
rect 20069 18400 20074 18456
rect 20130 18400 22558 18456
rect 22614 18400 22619 18456
rect 20069 18398 22619 18400
rect 20069 18395 20135 18398
rect 22553 18395 22619 18398
rect 26918 17988 26924 18052
rect 26988 18050 26994 18052
rect 27470 18050 27476 18052
rect 26988 17990 27476 18050
rect 26988 17988 26994 17990
rect 27470 17988 27476 17990
rect 27540 17988 27546 18052
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 17217 17914 17283 17917
rect 22645 17914 22711 17917
rect 17217 17912 22711 17914
rect 17217 17856 17222 17912
rect 17278 17856 22650 17912
rect 22706 17856 22711 17912
rect 17217 17854 22711 17856
rect 17217 17851 17283 17854
rect 22645 17851 22711 17854
rect 38101 17914 38167 17917
rect 39200 17914 40000 17944
rect 38101 17912 40000 17914
rect 38101 17856 38106 17912
rect 38162 17856 40000 17912
rect 38101 17854 40000 17856
rect 38101 17851 38167 17854
rect 39200 17824 40000 17854
rect 22001 17778 22067 17781
rect 27153 17778 27219 17781
rect 30230 17778 30236 17780
rect 22001 17776 30236 17778
rect 22001 17720 22006 17776
rect 22062 17720 27158 17776
rect 27214 17720 30236 17776
rect 22001 17718 30236 17720
rect 22001 17715 22067 17718
rect 27153 17715 27219 17718
rect 30230 17716 30236 17718
rect 30300 17716 30306 17780
rect 19517 17642 19583 17645
rect 27429 17642 27495 17645
rect 19517 17640 27495 17642
rect 19517 17584 19522 17640
rect 19578 17584 27434 17640
rect 27490 17584 27495 17640
rect 19517 17582 27495 17584
rect 19517 17579 19583 17582
rect 27429 17579 27495 17582
rect 29913 17642 29979 17645
rect 30046 17642 30052 17644
rect 29913 17640 30052 17642
rect 29913 17584 29918 17640
rect 29974 17584 30052 17640
rect 29913 17582 30052 17584
rect 29913 17579 29979 17582
rect 30046 17580 30052 17582
rect 30116 17580 30122 17644
rect 21265 17506 21331 17509
rect 24669 17506 24735 17509
rect 21265 17504 24735 17506
rect 21265 17448 21270 17504
rect 21326 17448 24674 17504
rect 24730 17448 24735 17504
rect 21265 17446 24735 17448
rect 21265 17443 21331 17446
rect 24669 17443 24735 17446
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 21081 17234 21147 17237
rect 28717 17234 28783 17237
rect 21081 17232 28783 17234
rect 21081 17176 21086 17232
rect 21142 17176 28722 17232
rect 28778 17176 28783 17232
rect 21081 17174 28783 17176
rect 21081 17171 21147 17174
rect 28717 17171 28783 17174
rect 27889 17098 27955 17101
rect 35157 17098 35223 17101
rect 27889 17096 35223 17098
rect 27889 17040 27894 17096
rect 27950 17040 35162 17096
rect 35218 17040 35223 17096
rect 27889 17038 35223 17040
rect 27889 17035 27955 17038
rect 35157 17035 35223 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 27429 16826 27495 16829
rect 28901 16826 28967 16829
rect 27429 16824 28967 16826
rect 27429 16768 27434 16824
rect 27490 16768 28906 16824
rect 28962 16768 28967 16824
rect 27429 16766 28967 16768
rect 27429 16763 27495 16766
rect 28901 16763 28967 16766
rect 28533 16690 28599 16693
rect 28901 16690 28967 16693
rect 28533 16688 28967 16690
rect 28533 16632 28538 16688
rect 28594 16632 28906 16688
rect 28962 16632 28967 16688
rect 28533 16630 28967 16632
rect 28533 16627 28599 16630
rect 28901 16627 28967 16630
rect 29729 16690 29795 16693
rect 30230 16690 30236 16692
rect 29729 16688 30236 16690
rect 29729 16632 29734 16688
rect 29790 16632 30236 16688
rect 29729 16630 30236 16632
rect 29729 16627 29795 16630
rect 30230 16628 30236 16630
rect 30300 16628 30306 16692
rect 29862 16492 29868 16556
rect 29932 16554 29938 16556
rect 31845 16554 31911 16557
rect 29932 16552 31911 16554
rect 29932 16496 31850 16552
rect 31906 16496 31911 16552
rect 29932 16494 31911 16496
rect 29932 16492 29938 16494
rect 31845 16491 31911 16494
rect 34646 16492 34652 16556
rect 34716 16554 34722 16556
rect 35157 16554 35223 16557
rect 34716 16552 35223 16554
rect 34716 16496 35162 16552
rect 35218 16496 35223 16552
rect 34716 16494 35223 16496
rect 34716 16492 34722 16494
rect 35157 16491 35223 16494
rect 38101 16554 38167 16557
rect 39200 16554 40000 16584
rect 38101 16552 40000 16554
rect 38101 16496 38106 16552
rect 38162 16496 40000 16552
rect 38101 16494 40000 16496
rect 38101 16491 38167 16494
rect 39200 16464 40000 16494
rect 26509 16418 26575 16421
rect 28901 16418 28967 16421
rect 26509 16416 28967 16418
rect 26509 16360 26514 16416
rect 26570 16360 28906 16416
rect 28962 16360 28967 16416
rect 26509 16358 28967 16360
rect 26509 16355 26575 16358
rect 28901 16355 28967 16358
rect 31477 16418 31543 16421
rect 35065 16418 35131 16421
rect 31477 16416 35131 16418
rect 31477 16360 31482 16416
rect 31538 16360 35070 16416
rect 35126 16360 35131 16416
rect 31477 16358 35131 16360
rect 31477 16355 31543 16358
rect 35065 16355 35131 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 26233 15330 26299 15333
rect 27838 15330 27844 15332
rect 26233 15328 27844 15330
rect 26233 15272 26238 15328
rect 26294 15272 27844 15328
rect 26233 15270 27844 15272
rect 26233 15267 26299 15270
rect 27838 15268 27844 15270
rect 27908 15268 27914 15332
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 8845 15196 8911 15197
rect 8845 15194 8892 15196
rect 8800 15192 8892 15194
rect 8800 15136 8850 15192
rect 8800 15134 8892 15136
rect 8845 15132 8892 15134
rect 8956 15132 8962 15196
rect 27153 15194 27219 15197
rect 27286 15194 27292 15196
rect 27153 15192 27292 15194
rect 27153 15136 27158 15192
rect 27214 15136 27292 15192
rect 27153 15134 27292 15136
rect 8845 15131 8911 15132
rect 27153 15131 27219 15134
rect 27286 15132 27292 15134
rect 27356 15132 27362 15196
rect 38101 15194 38167 15197
rect 39200 15194 40000 15224
rect 38101 15192 40000 15194
rect 38101 15136 38106 15192
rect 38162 15136 40000 15192
rect 38101 15134 40000 15136
rect 38101 15131 38167 15134
rect 39200 15104 40000 15134
rect 15193 15058 15259 15061
rect 17861 15058 17927 15061
rect 15193 15056 17927 15058
rect 15193 15000 15198 15056
rect 15254 15000 17866 15056
rect 17922 15000 17927 15056
rect 15193 14998 17927 15000
rect 15193 14995 15259 14998
rect 17861 14995 17927 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 21449 14514 21515 14517
rect 30925 14514 30991 14517
rect 21449 14512 30991 14514
rect 21449 14456 21454 14512
rect 21510 14456 30930 14512
rect 30986 14456 30991 14512
rect 21449 14454 30991 14456
rect 21449 14451 21515 14454
rect 30925 14451 30991 14454
rect 19517 14378 19583 14381
rect 19382 14376 19583 14378
rect 19382 14320 19522 14376
rect 19578 14320 19583 14376
rect 19382 14318 19583 14320
rect 19382 13973 19442 14318
rect 19517 14315 19583 14318
rect 33041 14378 33107 14381
rect 35157 14378 35223 14381
rect 33041 14376 35223 14378
rect 33041 14320 33046 14376
rect 33102 14320 35162 14376
rect 35218 14320 35223 14376
rect 33041 14318 35223 14320
rect 33041 14315 33107 14318
rect 35157 14315 35223 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 19382 13968 19491 13973
rect 19382 13912 19430 13968
rect 19486 13912 19491 13968
rect 19382 13910 19491 13912
rect 19425 13907 19491 13910
rect 38285 13834 38351 13837
rect 39200 13834 40000 13864
rect 38285 13832 40000 13834
rect 38285 13776 38290 13832
rect 38346 13776 40000 13832
rect 38285 13774 40000 13776
rect 38285 13771 38351 13774
rect 39200 13744 40000 13774
rect 25865 13698 25931 13701
rect 28349 13700 28415 13701
rect 25998 13698 26004 13700
rect 25865 13696 26004 13698
rect 25865 13640 25870 13696
rect 25926 13640 26004 13696
rect 25865 13638 26004 13640
rect 25865 13635 25931 13638
rect 25998 13636 26004 13638
rect 26068 13636 26074 13700
rect 28349 13696 28396 13700
rect 28460 13698 28466 13700
rect 28349 13640 28354 13696
rect 28349 13636 28396 13640
rect 28460 13638 28506 13698
rect 28460 13636 28466 13638
rect 28574 13636 28580 13700
rect 28644 13698 28650 13700
rect 29085 13698 29151 13701
rect 28644 13696 29151 13698
rect 28644 13640 29090 13696
rect 29146 13640 29151 13696
rect 28644 13638 29151 13640
rect 28644 13636 28650 13638
rect 28349 13635 28415 13636
rect 29085 13635 29151 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 19701 12882 19767 12885
rect 20253 12882 20319 12885
rect 25405 12882 25471 12885
rect 19701 12880 25471 12882
rect 19701 12824 19706 12880
rect 19762 12824 20258 12880
rect 20314 12824 25410 12880
rect 25466 12824 25471 12880
rect 19701 12822 25471 12824
rect 19701 12819 19767 12822
rect 20253 12819 20319 12822
rect 25405 12819 25471 12822
rect 21449 12610 21515 12613
rect 27797 12610 27863 12613
rect 21449 12608 27863 12610
rect 21449 12552 21454 12608
rect 21510 12552 27802 12608
rect 27858 12552 27863 12608
rect 21449 12550 27863 12552
rect 21449 12547 21515 12550
rect 27797 12547 27863 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 38285 12474 38351 12477
rect 39200 12474 40000 12504
rect 38285 12472 40000 12474
rect 38285 12416 38290 12472
rect 38346 12416 40000 12472
rect 38285 12414 40000 12416
rect 38285 12411 38351 12414
rect 39200 12384 40000 12414
rect 13997 12338 14063 12341
rect 17217 12338 17283 12341
rect 13997 12336 17283 12338
rect 13997 12280 14002 12336
rect 14058 12280 17222 12336
rect 17278 12280 17283 12336
rect 13997 12278 17283 12280
rect 13997 12275 14063 12278
rect 17217 12275 17283 12278
rect 27470 12276 27476 12340
rect 27540 12338 27546 12340
rect 27797 12338 27863 12341
rect 28257 12340 28323 12341
rect 28206 12338 28212 12340
rect 27540 12336 27863 12338
rect 27540 12280 27802 12336
rect 27858 12280 27863 12336
rect 27540 12278 27863 12280
rect 28166 12278 28212 12338
rect 28276 12336 28323 12340
rect 28318 12280 28323 12336
rect 27540 12276 27546 12278
rect 27797 12275 27863 12278
rect 28206 12276 28212 12278
rect 28276 12276 28323 12280
rect 28257 12275 28323 12276
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 38101 11114 38167 11117
rect 39200 11114 40000 11144
rect 38101 11112 40000 11114
rect 38101 11056 38106 11112
rect 38162 11056 40000 11112
rect 38101 11054 40000 11056
rect 38101 11051 38167 11054
rect 39200 11024 40000 11054
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 27102 10100 27108 10164
rect 27172 10162 27178 10164
rect 37825 10162 37891 10165
rect 27172 10160 37891 10162
rect 27172 10104 37830 10160
rect 37886 10104 37891 10160
rect 27172 10102 37891 10104
rect 27172 10100 27178 10102
rect 37825 10099 37891 10102
rect 30230 9828 30236 9892
rect 30300 9890 30306 9892
rect 37825 9890 37891 9893
rect 30300 9888 37891 9890
rect 30300 9832 37830 9888
rect 37886 9832 37891 9888
rect 30300 9830 37891 9832
rect 30300 9828 30306 9830
rect 37825 9827 37891 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 38101 9754 38167 9757
rect 39200 9754 40000 9784
rect 38101 9752 40000 9754
rect 38101 9696 38106 9752
rect 38162 9696 40000 9752
rect 38101 9694 40000 9696
rect 38101 9691 38167 9694
rect 39200 9664 40000 9694
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 38101 8394 38167 8397
rect 39200 8394 40000 8424
rect 38101 8392 40000 8394
rect 38101 8336 38106 8392
rect 38162 8336 40000 8392
rect 38101 8334 40000 8336
rect 38101 8331 38167 8334
rect 39200 8304 40000 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 38101 7034 38167 7037
rect 39200 7034 40000 7064
rect 38101 7032 40000 7034
rect 38101 6976 38106 7032
rect 38162 6976 40000 7032
rect 38101 6974 40000 6976
rect 38101 6971 38167 6974
rect 39200 6944 40000 6974
rect 14365 6762 14431 6765
rect 14733 6762 14799 6765
rect 18689 6762 18755 6765
rect 14365 6760 18755 6762
rect 14365 6704 14370 6760
rect 14426 6704 14738 6760
rect 14794 6704 18694 6760
rect 18750 6704 18755 6760
rect 14365 6702 18755 6704
rect 14365 6699 14431 6702
rect 14733 6699 14799 6702
rect 18689 6699 18755 6702
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 38101 5674 38167 5677
rect 39200 5674 40000 5704
rect 38101 5672 40000 5674
rect 38101 5616 38106 5672
rect 38162 5616 40000 5672
rect 38101 5614 40000 5616
rect 38101 5611 38167 5614
rect 39200 5584 40000 5614
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 38101 4314 38167 4317
rect 39200 4314 40000 4344
rect 38101 4312 40000 4314
rect 38101 4256 38106 4312
rect 38162 4256 40000 4312
rect 38101 4254 40000 4256
rect 38101 4251 38167 4254
rect 39200 4224 40000 4254
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 38101 2954 38167 2957
rect 39200 2954 40000 2984
rect 38101 2952 40000 2954
rect 38101 2896 38106 2952
rect 38162 2896 40000 2952
rect 38101 2894 40000 2896
rect 38101 2891 38167 2894
rect 39200 2864 40000 2894
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 38101 1594 38167 1597
rect 39200 1594 40000 1624
rect 38101 1592 40000 1594
rect 38101 1536 38106 1592
rect 38162 1536 40000 1592
rect 38101 1534 40000 1536
rect 38101 1531 38167 1534
rect 39200 1504 40000 1534
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 23980 35124 24044 35188
rect 30788 35048 30852 35052
rect 30788 34992 30802 35048
rect 30802 34992 30852 35048
rect 30788 34988 30852 34992
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 28028 34580 28092 34644
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 28764 34036 28828 34100
rect 20668 33900 20732 33964
rect 31340 33960 31404 33964
rect 31340 33904 31354 33960
rect 31354 33904 31404 33960
rect 31340 33900 31404 33904
rect 30052 33824 30116 33828
rect 30052 33768 30102 33824
rect 30102 33768 30116 33824
rect 30052 33764 30116 33768
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 27476 33356 27540 33420
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 32812 32812 32876 32876
rect 20484 32676 20548 32740
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 30604 32404 30668 32468
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 17172 31724 17236 31788
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 25820 31180 25884 31244
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 20484 30908 20548 30972
rect 20668 30908 20732 30972
rect 20116 30636 20180 30700
rect 35572 30696 35636 30700
rect 35572 30640 35586 30696
rect 35586 30640 35636 30696
rect 35572 30636 35636 30640
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 28028 30228 28092 30292
rect 30236 29956 30300 30020
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 31156 29684 31220 29748
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 20116 29004 20180 29068
rect 29500 29064 29564 29068
rect 29500 29008 29550 29064
rect 29550 29008 29564 29064
rect 29500 29004 29564 29008
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 22692 28052 22756 28116
rect 27292 27780 27356 27844
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 26004 27644 26068 27708
rect 28396 27644 28460 27708
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 8892 26692 8956 26756
rect 34652 26752 34716 26756
rect 34652 26696 34666 26752
rect 34666 26696 34716 26752
rect 34652 26692 34716 26696
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 29868 26284 29932 26348
rect 31156 26148 31220 26212
rect 34652 26284 34716 26348
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 27844 26012 27908 26076
rect 17172 25876 17236 25940
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 28580 24924 28644 24988
rect 27476 24848 27540 24852
rect 27476 24792 27490 24848
rect 27490 24792 27540 24848
rect 27476 24788 27540 24792
rect 32812 24788 32876 24852
rect 22692 24712 22756 24716
rect 22692 24656 22742 24712
rect 22742 24656 22756 24712
rect 22692 24652 22756 24656
rect 28028 24652 28092 24716
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 28764 23760 28828 23764
rect 28764 23704 28778 23760
rect 28778 23704 28828 23760
rect 28764 23700 28828 23704
rect 26924 23564 26988 23628
rect 30604 23428 30668 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 30052 23292 30116 23356
rect 30052 23020 30116 23084
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 29500 22612 29564 22676
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 28212 22204 28276 22268
rect 23980 21932 24044 21996
rect 30788 21932 30852 21996
rect 31340 21796 31404 21860
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 27108 20768 27172 20772
rect 27108 20712 27122 20768
rect 27122 20712 27172 20768
rect 27108 20708 27172 20712
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 25820 20572 25884 20636
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 26924 18804 26988 18868
rect 35572 18804 35636 18868
rect 30236 18668 30300 18732
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 26924 17988 26988 18052
rect 27476 17988 27540 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 30236 17716 30300 17780
rect 30052 17580 30116 17644
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 30236 16628 30300 16692
rect 29868 16492 29932 16556
rect 34652 16492 34716 16556
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 27844 15268 27908 15332
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 8892 15192 8956 15196
rect 8892 15136 8906 15192
rect 8906 15136 8956 15192
rect 8892 15132 8956 15136
rect 27292 15132 27356 15196
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 26004 13636 26068 13700
rect 28396 13696 28460 13700
rect 28396 13640 28410 13696
rect 28410 13640 28460 13696
rect 28396 13636 28460 13640
rect 28580 13636 28644 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 27476 12276 27540 12340
rect 28212 12336 28276 12340
rect 28212 12280 28262 12336
rect 28262 12280 28276 12336
rect 28212 12276 28276 12280
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 27108 10100 27172 10164
rect 30236 9828 30300 9892
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 23979 35188 24045 35189
rect 23979 35124 23980 35188
rect 24044 35124 24045 35188
rect 23979 35123 24045 35124
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 20667 33964 20733 33965
rect 20667 33900 20668 33964
rect 20732 33900 20733 33964
rect 20667 33899 20733 33900
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 20483 32740 20549 32741
rect 20483 32676 20484 32740
rect 20548 32676 20549 32740
rect 20483 32675 20549 32676
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 17171 31788 17237 31789
rect 17171 31724 17172 31788
rect 17236 31724 17237 31788
rect 17171 31723 17237 31724
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 8891 26756 8957 26757
rect 8891 26692 8892 26756
rect 8956 26692 8957 26756
rect 8891 26691 8957 26692
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 8894 15197 8954 26691
rect 17174 25941 17234 31723
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 20486 30973 20546 32675
rect 20670 30973 20730 33899
rect 20483 30972 20549 30973
rect 20483 30908 20484 30972
rect 20548 30908 20549 30972
rect 20483 30907 20549 30908
rect 20667 30972 20733 30973
rect 20667 30908 20668 30972
rect 20732 30908 20733 30972
rect 20667 30907 20733 30908
rect 20115 30700 20181 30701
rect 20115 30636 20116 30700
rect 20180 30636 20181 30700
rect 20115 30635 20181 30636
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 20118 29069 20178 30635
rect 20115 29068 20181 29069
rect 20115 29004 20116 29068
rect 20180 29004 20181 29068
rect 20115 29003 20181 29004
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 22691 28116 22757 28117
rect 22691 28052 22692 28116
rect 22756 28052 22757 28116
rect 22691 28051 22757 28052
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 17171 25940 17237 25941
rect 17171 25876 17172 25940
rect 17236 25876 17237 25940
rect 17171 25875 17237 25876
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 22694 24717 22754 28051
rect 22691 24716 22757 24717
rect 22691 24652 22692 24716
rect 22756 24652 22757 24716
rect 22691 24651 22757 24652
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 23982 21997 24042 35123
rect 30787 35052 30853 35053
rect 30787 34988 30788 35052
rect 30852 34988 30853 35052
rect 30787 34987 30853 34988
rect 28027 34644 28093 34645
rect 28027 34580 28028 34644
rect 28092 34580 28093 34644
rect 28027 34579 28093 34580
rect 27475 33420 27541 33421
rect 27475 33356 27476 33420
rect 27540 33356 27541 33420
rect 27475 33355 27541 33356
rect 25819 31244 25885 31245
rect 25819 31180 25820 31244
rect 25884 31180 25885 31244
rect 25819 31179 25885 31180
rect 23979 21996 24045 21997
rect 23979 21932 23980 21996
rect 24044 21932 24045 21996
rect 23979 21931 24045 21932
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 25822 20637 25882 31179
rect 27291 27844 27357 27845
rect 27291 27780 27292 27844
rect 27356 27780 27357 27844
rect 27291 27779 27357 27780
rect 26003 27708 26069 27709
rect 26003 27644 26004 27708
rect 26068 27644 26069 27708
rect 26003 27643 26069 27644
rect 25819 20636 25885 20637
rect 25819 20572 25820 20636
rect 25884 20572 25885 20636
rect 25819 20571 25885 20572
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 8891 15196 8957 15197
rect 8891 15132 8892 15196
rect 8956 15132 8957 15196
rect 8891 15131 8957 15132
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 26006 13701 26066 27643
rect 26923 23628 26989 23629
rect 26923 23564 26924 23628
rect 26988 23564 26989 23628
rect 26923 23563 26989 23564
rect 26926 18869 26986 23563
rect 27107 20772 27173 20773
rect 27107 20708 27108 20772
rect 27172 20708 27173 20772
rect 27107 20707 27173 20708
rect 26923 18868 26989 18869
rect 26923 18804 26924 18868
rect 26988 18804 26989 18868
rect 26923 18803 26989 18804
rect 26926 18053 26986 18803
rect 26923 18052 26989 18053
rect 26923 17988 26924 18052
rect 26988 17988 26989 18052
rect 26923 17987 26989 17988
rect 26003 13700 26069 13701
rect 26003 13636 26004 13700
rect 26068 13636 26069 13700
rect 26003 13635 26069 13636
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 27110 10165 27170 20707
rect 27294 15197 27354 27779
rect 27478 24853 27538 33355
rect 28030 30293 28090 34579
rect 28763 34100 28829 34101
rect 28763 34036 28764 34100
rect 28828 34036 28829 34100
rect 28763 34035 28829 34036
rect 28027 30292 28093 30293
rect 28027 30228 28028 30292
rect 28092 30228 28093 30292
rect 28027 30227 28093 30228
rect 27843 26076 27909 26077
rect 27843 26012 27844 26076
rect 27908 26012 27909 26076
rect 27843 26011 27909 26012
rect 27475 24852 27541 24853
rect 27475 24788 27476 24852
rect 27540 24788 27541 24852
rect 27475 24787 27541 24788
rect 27475 18052 27541 18053
rect 27475 17988 27476 18052
rect 27540 17988 27541 18052
rect 27475 17987 27541 17988
rect 27291 15196 27357 15197
rect 27291 15132 27292 15196
rect 27356 15132 27357 15196
rect 27291 15131 27357 15132
rect 27478 12341 27538 17987
rect 27846 15333 27906 26011
rect 28030 24717 28090 30227
rect 28395 27708 28461 27709
rect 28395 27644 28396 27708
rect 28460 27644 28461 27708
rect 28395 27643 28461 27644
rect 28027 24716 28093 24717
rect 28027 24652 28028 24716
rect 28092 24652 28093 24716
rect 28027 24651 28093 24652
rect 28211 22268 28277 22269
rect 28211 22204 28212 22268
rect 28276 22204 28277 22268
rect 28211 22203 28277 22204
rect 27843 15332 27909 15333
rect 27843 15268 27844 15332
rect 27908 15268 27909 15332
rect 27843 15267 27909 15268
rect 28214 12341 28274 22203
rect 28398 13701 28458 27643
rect 28579 24988 28645 24989
rect 28579 24924 28580 24988
rect 28644 24924 28645 24988
rect 28579 24923 28645 24924
rect 28582 13701 28642 24923
rect 28766 23765 28826 34035
rect 30051 33828 30117 33829
rect 30051 33764 30052 33828
rect 30116 33764 30117 33828
rect 30051 33763 30117 33764
rect 29499 29068 29565 29069
rect 29499 29004 29500 29068
rect 29564 29004 29565 29068
rect 29499 29003 29565 29004
rect 28763 23764 28829 23765
rect 28763 23700 28764 23764
rect 28828 23700 28829 23764
rect 28763 23699 28829 23700
rect 29502 22677 29562 29003
rect 29867 26348 29933 26349
rect 29867 26284 29868 26348
rect 29932 26284 29933 26348
rect 29867 26283 29933 26284
rect 29499 22676 29565 22677
rect 29499 22612 29500 22676
rect 29564 22612 29565 22676
rect 29499 22611 29565 22612
rect 29870 16557 29930 26283
rect 30054 23357 30114 33763
rect 30603 32468 30669 32469
rect 30603 32404 30604 32468
rect 30668 32404 30669 32468
rect 30603 32403 30669 32404
rect 30235 30020 30301 30021
rect 30235 29956 30236 30020
rect 30300 29956 30301 30020
rect 30235 29955 30301 29956
rect 30051 23356 30117 23357
rect 30051 23292 30052 23356
rect 30116 23292 30117 23356
rect 30051 23291 30117 23292
rect 30051 23084 30117 23085
rect 30051 23020 30052 23084
rect 30116 23020 30117 23084
rect 30051 23019 30117 23020
rect 30054 17645 30114 23019
rect 30238 18733 30298 29955
rect 30606 23493 30666 32403
rect 30603 23492 30669 23493
rect 30603 23428 30604 23492
rect 30668 23428 30669 23492
rect 30603 23427 30669 23428
rect 30790 21997 30850 34987
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 31339 33964 31405 33965
rect 31339 33900 31340 33964
rect 31404 33900 31405 33964
rect 31339 33899 31405 33900
rect 31155 29748 31221 29749
rect 31155 29684 31156 29748
rect 31220 29684 31221 29748
rect 31155 29683 31221 29684
rect 31158 26213 31218 29683
rect 31155 26212 31221 26213
rect 31155 26148 31156 26212
rect 31220 26148 31221 26212
rect 31155 26147 31221 26148
rect 30787 21996 30853 21997
rect 30787 21932 30788 21996
rect 30852 21932 30853 21996
rect 30787 21931 30853 21932
rect 31342 21861 31402 33899
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 32811 32876 32877 32877
rect 32811 32812 32812 32876
rect 32876 32812 32877 32876
rect 32811 32811 32877 32812
rect 32814 24853 32874 32811
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 35571 30700 35637 30701
rect 35571 30636 35572 30700
rect 35636 30636 35637 30700
rect 35571 30635 35637 30636
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34651 26756 34717 26757
rect 34651 26692 34652 26756
rect 34716 26692 34717 26756
rect 34651 26691 34717 26692
rect 34654 26349 34714 26691
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34651 26348 34717 26349
rect 34651 26284 34652 26348
rect 34716 26284 34717 26348
rect 34651 26283 34717 26284
rect 32811 24852 32877 24853
rect 32811 24788 32812 24852
rect 32876 24788 32877 24852
rect 32811 24787 32877 24788
rect 31339 21860 31405 21861
rect 31339 21796 31340 21860
rect 31404 21796 31405 21860
rect 31339 21795 31405 21796
rect 30235 18732 30301 18733
rect 30235 18668 30236 18732
rect 30300 18668 30301 18732
rect 30235 18667 30301 18668
rect 30238 17781 30298 18667
rect 30235 17780 30301 17781
rect 30235 17716 30236 17780
rect 30300 17716 30301 17780
rect 30235 17715 30301 17716
rect 30051 17644 30117 17645
rect 30051 17580 30052 17644
rect 30116 17580 30117 17644
rect 30051 17579 30117 17580
rect 30235 16692 30301 16693
rect 30235 16628 30236 16692
rect 30300 16628 30301 16692
rect 30235 16627 30301 16628
rect 29867 16556 29933 16557
rect 29867 16492 29868 16556
rect 29932 16492 29933 16556
rect 29867 16491 29933 16492
rect 28395 13700 28461 13701
rect 28395 13636 28396 13700
rect 28460 13636 28461 13700
rect 28395 13635 28461 13636
rect 28579 13700 28645 13701
rect 28579 13636 28580 13700
rect 28644 13636 28645 13700
rect 28579 13635 28645 13636
rect 27475 12340 27541 12341
rect 27475 12276 27476 12340
rect 27540 12276 27541 12340
rect 27475 12275 27541 12276
rect 28211 12340 28277 12341
rect 28211 12276 28212 12340
rect 28276 12276 28277 12340
rect 28211 12275 28277 12276
rect 27107 10164 27173 10165
rect 27107 10100 27108 10164
rect 27172 10100 27173 10164
rect 27107 10099 27173 10100
rect 30238 9893 30298 16627
rect 34654 16557 34714 26283
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 35574 18869 35634 30635
rect 35571 18868 35637 18869
rect 35571 18804 35572 18868
rect 35636 18804 35637 18868
rect 35571 18803 35637 18804
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34651 16556 34717 16557
rect 34651 16492 34652 16556
rect 34716 16492 34717 16556
rect 34651 16491 34717 16492
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 30235 9892 30301 9893
rect 30235 9828 30236 9892
rect 30300 9828 30301 9892
rect 30235 9827 30301 9828
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30728 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 13892 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1676037725
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1676037725
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1676037725
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1676037725
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1676037725
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1676037725
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1676037725
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1676037725
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1676037725
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1676037725
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_393 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1676037725
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_401
timestamp 1676037725
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_204
timestamp 1676037725
transform 1 0 19872 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_289
timestamp 1676037725
transform 1 0 27692 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_300
timestamp 1676037725
transform 1 0 28704 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_312
timestamp 1676037725
transform 1 0 29808 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_322
timestamp 1676037725
transform 1 0 30728 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1676037725
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_369
timestamp 1676037725
transform 1 0 35052 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_381
timestamp 1676037725
transform 1 0 36156 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_389
timestamp 1676037725
transform 1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_180
timestamp 1676037725
transform 1 0 17664 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1676037725
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_237
timestamp 1676037725
transform 1 0 22908 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_247
timestamp 1676037725
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_282
timestamp 1676037725
transform 1 0 27048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_302
timestamp 1676037725
transform 1 0 28888 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_327
timestamp 1676037725
transform 1 0 31188 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_339
timestamp 1676037725
transform 1 0 32292 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_351
timestamp 1676037725
transform 1 0 33396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_373
timestamp 1676037725
transform 1 0 35420 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_384
timestamp 1676037725
transform 1 0 36432 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_396
timestamp 1676037725
transform 1 0 37536 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1676037725
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_190
timestamp 1676037725
transform 1 0 18584 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_221
timestamp 1676037725
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_245
timestamp 1676037725
transform 1 0 23644 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_265
timestamp 1676037725
transform 1 0 25484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1676037725
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_328
timestamp 1676037725
transform 1 0 31280 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_355
timestamp 1676037725
transform 1 0 33764 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_367
timestamp 1676037725
transform 1 0 34868 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_387
timestamp 1676037725
transform 1 0 36708 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_404
timestamp 1676037725
transform 1 0 38272 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_175
timestamp 1676037725
transform 1 0 17204 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_183
timestamp 1676037725
transform 1 0 17940 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_234
timestamp 1676037725
transform 1 0 22632 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_246
timestamp 1676037725
transform 1 0 23736 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_264
timestamp 1676037725
transform 1 0 25392 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_272
timestamp 1676037725
transform 1 0 26128 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_284
timestamp 1676037725
transform 1 0 27232 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_292
timestamp 1676037725
transform 1 0 27968 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_302
timestamp 1676037725
transform 1 0 28888 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_317
timestamp 1676037725
transform 1 0 30268 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_335
timestamp 1676037725
transform 1 0 31924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_347
timestamp 1676037725
transform 1 0 33028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1676037725
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_372
timestamp 1676037725
transform 1 0 35328 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_384
timestamp 1676037725
transform 1 0 36432 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_388
timestamp 1676037725
transform 1 0 36800 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1676037725
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_155
timestamp 1676037725
transform 1 0 15364 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_163
timestamp 1676037725
transform 1 0 16100 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_214
timestamp 1676037725
transform 1 0 20792 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_221
timestamp 1676037725
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_250
timestamp 1676037725
transform 1 0 24104 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_258
timestamp 1676037725
transform 1 0 24840 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_266
timestamp 1676037725
transform 1 0 25576 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_275
timestamp 1676037725
transform 1 0 26404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_285
timestamp 1676037725
transform 1 0 27324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_302
timestamp 1676037725
transform 1 0 28888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_315
timestamp 1676037725
transform 1 0 30084 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_328
timestamp 1676037725
transform 1 0 31280 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_358
timestamp 1676037725
transform 1 0 34040 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_374
timestamp 1676037725
transform 1 0 35512 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_386
timestamp 1676037725
transform 1 0 36616 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_117
timestamp 1676037725
transform 1 0 11868 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_125
timestamp 1676037725
transform 1 0 12604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1676037725
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_150
timestamp 1676037725
transform 1 0 14904 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_169
timestamp 1676037725
transform 1 0 16652 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_190
timestamp 1676037725
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_218
timestamp 1676037725
transform 1 0 21160 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_225
timestamp 1676037725
transform 1 0 21804 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_231
timestamp 1676037725
transform 1 0 22356 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1676037725
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_259
timestamp 1676037725
transform 1 0 24932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_269
timestamp 1676037725
transform 1 0 25852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_284
timestamp 1676037725
transform 1 0 27232 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_295
timestamp 1676037725
transform 1 0 28244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_323
timestamp 1676037725
transform 1 0 30820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_335
timestamp 1676037725
transform 1 0 31924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_343
timestamp 1676037725
transform 1 0 32660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_355
timestamp 1676037725
transform 1 0 33764 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_375
timestamp 1676037725
transform 1 0 35604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_403
timestamp 1676037725
transform 1 0 38180 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_134
timestamp 1676037725
transform 1 0 13432 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_155
timestamp 1676037725
transform 1 0 15364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_179
timestamp 1676037725
transform 1 0 17572 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_200
timestamp 1676037725
transform 1 0 19504 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_204
timestamp 1676037725
transform 1 0 19872 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_213
timestamp 1676037725
transform 1 0 20700 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_254
timestamp 1676037725
transform 1 0 24472 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_266
timestamp 1676037725
transform 1 0 25576 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1676037725
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_316
timestamp 1676037725
transform 1 0 30176 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_328
timestamp 1676037725
transform 1 0 31280 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_356
timestamp 1676037725
transform 1 0 33856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_362
timestamp 1676037725
transform 1 0 34408 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_371
timestamp 1676037725
transform 1 0 35236 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_383
timestamp 1676037725
transform 1 0 36340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_404
timestamp 1676037725
transform 1 0 38272 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_115
timestamp 1676037725
transform 1 0 11684 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_122
timestamp 1676037725
transform 1 0 12328 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_130
timestamp 1676037725
transform 1 0 13064 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_158
timestamp 1676037725
transform 1 0 15640 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_162
timestamp 1676037725
transform 1 0 16008 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_171
timestamp 1676037725
transform 1 0 16836 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_181
timestamp 1676037725
transform 1 0 17756 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1676037725
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_203
timestamp 1676037725
transform 1 0 19780 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_219
timestamp 1676037725
transform 1 0 21252 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_239
timestamp 1676037725
transform 1 0 23092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_273
timestamp 1676037725
transform 1 0 26220 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_292
timestamp 1676037725
transform 1 0 27968 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1676037725
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_337
timestamp 1676037725
transform 1 0 32108 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_360
timestamp 1676037725
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_378
timestamp 1676037725
transform 1 0 35880 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_386
timestamp 1676037725
transform 1 0 36616 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1676037725
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_120
timestamp 1676037725
transform 1 0 12144 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_132
timestamp 1676037725
transform 1 0 13248 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_138
timestamp 1676037725
transform 1 0 13800 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_150
timestamp 1676037725
transform 1 0 14904 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_162
timestamp 1676037725
transform 1 0 16008 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_176
timestamp 1676037725
transform 1 0 17296 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_188
timestamp 1676037725
transform 1 0 18400 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_196
timestamp 1676037725
transform 1 0 19136 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_204
timestamp 1676037725
transform 1 0 19872 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_213
timestamp 1676037725
transform 1 0 20700 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_232
timestamp 1676037725
transform 1 0 22448 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_244
timestamp 1676037725
transform 1 0 23552 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_252
timestamp 1676037725
transform 1 0 24288 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_270
timestamp 1676037725
transform 1 0 25944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1676037725
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_292
timestamp 1676037725
transform 1 0 27968 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_313
timestamp 1676037725
transform 1 0 29900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp 1676037725
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_350
timestamp 1676037725
transform 1 0 33304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_354
timestamp 1676037725
transform 1 0 33672 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_360
timestamp 1676037725
transform 1 0 34224 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_382
timestamp 1676037725
transform 1 0 36248 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_390
timestamp 1676037725
transform 1 0 36984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_404
timestamp 1676037725
transform 1 0 38272 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_101
timestamp 1676037725
transform 1 0 10396 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_107
timestamp 1676037725
transform 1 0 10948 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_119
timestamp 1676037725
transform 1 0 12052 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_150
timestamp 1676037725
transform 1 0 14904 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_161
timestamp 1676037725
transform 1 0 15916 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_174
timestamp 1676037725
transform 1 0 17112 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_181
timestamp 1676037725
transform 1 0 17756 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_208
timestamp 1676037725
transform 1 0 20240 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_212
timestamp 1676037725
transform 1 0 20608 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_222
timestamp 1676037725
transform 1 0 21528 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_234
timestamp 1676037725
transform 1 0 22632 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_246
timestamp 1676037725
transform 1 0 23736 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_259
timestamp 1676037725
transform 1 0 24932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_269
timestamp 1676037725
transform 1 0 25852 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_279
timestamp 1676037725
transform 1 0 26772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_291
timestamp 1676037725
transform 1 0 27876 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1676037725
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1676037725
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_313
timestamp 1676037725
transform 1 0 29900 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_321
timestamp 1676037725
transform 1 0 30636 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_343
timestamp 1676037725
transform 1 0 32660 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_352
timestamp 1676037725
transform 1 0 33488 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_371
timestamp 1676037725
transform 1 0 35236 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_393
timestamp 1676037725
transform 1 0 37260 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1676037725
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_101
timestamp 1676037725
transform 1 0 10396 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1676037725
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_124
timestamp 1676037725
transform 1 0 12512 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_128
timestamp 1676037725
transform 1 0 12880 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_148
timestamp 1676037725
transform 1 0 14720 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_185
timestamp 1676037725
transform 1 0 18124 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_202
timestamp 1676037725
transform 1 0 19688 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_210
timestamp 1676037725
transform 1 0 20424 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_233
timestamp 1676037725
transform 1 0 22540 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_251
timestamp 1676037725
transform 1 0 24196 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_264
timestamp 1676037725
transform 1 0 25392 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1676037725
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_301
timestamp 1676037725
transform 1 0 28796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_313
timestamp 1676037725
transform 1 0 29900 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_324
timestamp 1676037725
transform 1 0 30912 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_348
timestamp 1676037725
transform 1 0 33120 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_368
timestamp 1676037725
transform 1 0 34960 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_380
timestamp 1676037725
transform 1 0 36064 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_106
timestamp 1676037725
transform 1 0 10856 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_114
timestamp 1676037725
transform 1 0 11592 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_126
timestamp 1676037725
transform 1 0 12696 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_130
timestamp 1676037725
transform 1 0 13064 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1676037725
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_149
timestamp 1676037725
transform 1 0 14812 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_160
timestamp 1676037725
transform 1 0 15824 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_171
timestamp 1676037725
transform 1 0 16836 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_182
timestamp 1676037725
transform 1 0 17848 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_190
timestamp 1676037725
transform 1 0 18584 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_221
timestamp 1676037725
transform 1 0 21436 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_228
timestamp 1676037725
transform 1 0 22080 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_235
timestamp 1676037725
transform 1 0 22724 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_247
timestamp 1676037725
transform 1 0 23828 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_261
timestamp 1676037725
transform 1 0 25116 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_269
timestamp 1676037725
transform 1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_283
timestamp 1676037725
transform 1 0 27140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_295
timestamp 1676037725
transform 1 0 28244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1676037725
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1676037725
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_333
timestamp 1676037725
transform 1 0 31740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_342
timestamp 1676037725
transform 1 0 32568 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_362
timestamp 1676037725
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_389
timestamp 1676037725
transform 1 0 36892 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_397
timestamp 1676037725
transform 1 0 37628 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_405
timestamp 1676037725
transform 1 0 38364 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_119
timestamp 1676037725
transform 1 0 12052 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_136
timestamp 1676037725
transform 1 0 13616 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_148
timestamp 1676037725
transform 1 0 14720 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_154
timestamp 1676037725
transform 1 0 15272 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_158
timestamp 1676037725
transform 1 0 15640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_175
timestamp 1676037725
transform 1 0 17204 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_185
timestamp 1676037725
transform 1 0 18124 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_197
timestamp 1676037725
transform 1 0 19228 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1676037725
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_234
timestamp 1676037725
transform 1 0 22632 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_246
timestamp 1676037725
transform 1 0 23736 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_254
timestamp 1676037725
transform 1 0 24472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_271
timestamp 1676037725
transform 1 0 26036 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1676037725
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_292
timestamp 1676037725
transform 1 0 27968 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_316
timestamp 1676037725
transform 1 0 30176 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_328
timestamp 1676037725
transform 1 0 31280 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_349
timestamp 1676037725
transform 1 0 33212 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_355
timestamp 1676037725
transform 1 0 33764 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_365
timestamp 1676037725
transform 1 0 34684 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_377
timestamp 1676037725
transform 1 0 35788 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_389
timestamp 1676037725
transform 1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_404
timestamp 1676037725
transform 1 0 38272 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_103
timestamp 1676037725
transform 1 0 10580 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_114
timestamp 1676037725
transform 1 0 11592 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_120
timestamp 1676037725
transform 1 0 12144 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_125
timestamp 1676037725
transform 1 0 12604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1676037725
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_149
timestamp 1676037725
transform 1 0 14812 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_155
timestamp 1676037725
transform 1 0 15364 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_170
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_177
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_187
timestamp 1676037725
transform 1 0 18308 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1676037725
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_204
timestamp 1676037725
transform 1 0 19872 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_216
timestamp 1676037725
transform 1 0 20976 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_229
timestamp 1676037725
transform 1 0 22172 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_241
timestamp 1676037725
transform 1 0 23276 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_249
timestamp 1676037725
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_268
timestamp 1676037725
transform 1 0 25760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_276
timestamp 1676037725
transform 1 0 26496 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_294
timestamp 1676037725
transform 1 0 28152 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1676037725
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_332
timestamp 1676037725
transform 1 0 31648 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_344
timestamp 1676037725
transform 1 0 32752 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_359
timestamp 1676037725
transform 1 0 34132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1676037725
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_383
timestamp 1676037725
transform 1 0 36340 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_403
timestamp 1676037725
transform 1 0 38180 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_73
timestamp 1676037725
transform 1 0 7820 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_90
timestamp 1676037725
transform 1 0 9384 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_98
timestamp 1676037725
transform 1 0 10120 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1676037725
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1676037725
transform 1 0 12236 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_127
timestamp 1676037725
transform 1 0 12788 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_139
timestamp 1676037725
transform 1 0 13892 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_147
timestamp 1676037725
transform 1 0 14628 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_157
timestamp 1676037725
transform 1 0 15548 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 1676037725
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_177
timestamp 1676037725
transform 1 0 17388 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_183
timestamp 1676037725
transform 1 0 17940 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_191
timestamp 1676037725
transform 1 0 18676 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_197
timestamp 1676037725
transform 1 0 19228 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_207
timestamp 1676037725
transform 1 0 20148 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_219
timestamp 1676037725
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1676037725
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_253
timestamp 1676037725
transform 1 0 24380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_266
timestamp 1676037725
transform 1 0 25576 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_275
timestamp 1676037725
transform 1 0 26404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1676037725
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_293
timestamp 1676037725
transform 1 0 28060 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_301
timestamp 1676037725
transform 1 0 28796 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_311
timestamp 1676037725
transform 1 0 29716 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_317
timestamp 1676037725
transform 1 0 30268 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1676037725
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_360
timestamp 1676037725
transform 1 0 34224 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_368
timestamp 1676037725
transform 1 0 34960 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1676037725
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_404
timestamp 1676037725
transform 1 0 38272 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_94
timestamp 1676037725
transform 1 0 9752 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_106
timestamp 1676037725
transform 1 0 10856 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_118
timestamp 1676037725
transform 1 0 11960 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_124
timestamp 1676037725
transform 1 0 12512 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_130
timestamp 1676037725
transform 1 0 13064 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_134
timestamp 1676037725
transform 1 0 13432 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_149
timestamp 1676037725
transform 1 0 14812 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_159
timestamp 1676037725
transform 1 0 15732 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_163
timestamp 1676037725
transform 1 0 16100 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_168
timestamp 1676037725
transform 1 0 16560 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_179
timestamp 1676037725
transform 1 0 17572 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_187
timestamp 1676037725
transform 1 0 18308 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_206
timestamp 1676037725
transform 1 0 20056 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_214
timestamp 1676037725
transform 1 0 20792 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_222
timestamp 1676037725
transform 1 0 21528 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_229
timestamp 1676037725
transform 1 0 22172 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_241
timestamp 1676037725
transform 1 0 23276 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_249
timestamp 1676037725
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_259
timestamp 1676037725
transform 1 0 24932 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_272
timestamp 1676037725
transform 1 0 26128 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_284
timestamp 1676037725
transform 1 0 27232 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_292
timestamp 1676037725
transform 1 0 27968 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_299
timestamp 1676037725
transform 1 0 28612 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1676037725
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_321
timestamp 1676037725
transform 1 0 30636 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_325
timestamp 1676037725
transform 1 0 31004 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_335
timestamp 1676037725
transform 1 0 31924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1676037725
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1676037725
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_377
timestamp 1676037725
transform 1 0 35788 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_385
timestamp 1676037725
transform 1 0 36524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_404
timestamp 1676037725
transform 1 0 38272 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_87
timestamp 1676037725
transform 1 0 9108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_121
timestamp 1676037725
transform 1 0 12236 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_128
timestamp 1676037725
transform 1 0 12880 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_138
timestamp 1676037725
transform 1 0 13800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_150
timestamp 1676037725
transform 1 0 14904 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp 1676037725
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_182
timestamp 1676037725
transform 1 0 17848 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_194
timestamp 1676037725
transform 1 0 18952 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_204
timestamp 1676037725
transform 1 0 19872 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_212
timestamp 1676037725
transform 1 0 20608 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_233
timestamp 1676037725
transform 1 0 22540 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_245
timestamp 1676037725
transform 1 0 23644 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_257
timestamp 1676037725
transform 1 0 24748 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_270
timestamp 1676037725
transform 1 0 25944 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1676037725
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_296
timestamp 1676037725
transform 1 0 28336 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_307
timestamp 1676037725
transform 1 0 29348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_319
timestamp 1676037725
transform 1 0 30452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_331
timestamp 1676037725
transform 1 0 31556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1676037725
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_341
timestamp 1676037725
transform 1 0 32476 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_351
timestamp 1676037725
transform 1 0 33396 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_363
timestamp 1676037725
transform 1 0 34500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_375
timestamp 1676037725
transform 1 0 35604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_387
timestamp 1676037725
transform 1 0 36708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1676037725
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_401
timestamp 1676037725
transform 1 0 37996 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1676037725
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_106
timestamp 1676037725
transform 1 0 10856 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_118
timestamp 1676037725
transform 1 0 11960 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_131
timestamp 1676037725
transform 1 0 13156 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_150
timestamp 1676037725
transform 1 0 14904 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_158
timestamp 1676037725
transform 1 0 15640 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_176
timestamp 1676037725
transform 1 0 17296 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_187
timestamp 1676037725
transform 1 0 18308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1676037725
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_209
timestamp 1676037725
transform 1 0 20332 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_218
timestamp 1676037725
transform 1 0 21160 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_226
timestamp 1676037725
transform 1 0 21896 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_238
timestamp 1676037725
transform 1 0 23000 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1676037725
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_265
timestamp 1676037725
transform 1 0 25484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_273
timestamp 1676037725
transform 1 0 26220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_277
timestamp 1676037725
transform 1 0 26588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_285
timestamp 1676037725
transform 1 0 27324 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1676037725
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1676037725
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_317
timestamp 1676037725
transform 1 0 30268 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_332
timestamp 1676037725
transform 1 0 31648 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_344
timestamp 1676037725
transform 1 0 32752 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_356
timestamp 1676037725
transform 1 0 33856 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_373
timestamp 1676037725
transform 1 0 35420 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_393
timestamp 1676037725
transform 1 0 37260 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_405
timestamp 1676037725
transform 1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_73
timestamp 1676037725
transform 1 0 7820 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_90
timestamp 1676037725
transform 1 0 9384 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_98
timestamp 1676037725
transform 1 0 10120 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1676037725
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_121
timestamp 1676037725
transform 1 0 12236 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_139
timestamp 1676037725
transform 1 0 13892 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1676037725
transform 1 0 15824 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_179
timestamp 1676037725
transform 1 0 17572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_191
timestamp 1676037725
transform 1 0 18676 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1676037725
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1676037725
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1676037725
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_233
timestamp 1676037725
transform 1 0 22540 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_242
timestamp 1676037725
transform 1 0 23368 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_254
timestamp 1676037725
transform 1 0 24472 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_261
timestamp 1676037725
transform 1 0 25116 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 1676037725
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_287
timestamp 1676037725
transform 1 0 27508 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_291
timestamp 1676037725
transform 1 0 27876 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_307
timestamp 1676037725
transform 1 0 29348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_315
timestamp 1676037725
transform 1 0 30084 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1676037725
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_343
timestamp 1676037725
transform 1 0 32660 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_352
timestamp 1676037725
transform 1 0 33488 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_373
timestamp 1676037725
transform 1 0 35420 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1676037725
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1676037725
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_401
timestamp 1676037725
transform 1 0 37996 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1676037725
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1676037725
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_109
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_122
timestamp 1676037725
transform 1 0 12328 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_130
timestamp 1676037725
transform 1 0 13064 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1676037725
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_159
timestamp 1676037725
transform 1 0 15732 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_171
timestamp 1676037725
transform 1 0 16836 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_183
timestamp 1676037725
transform 1 0 17940 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_229
timestamp 1676037725
transform 1 0 22172 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_260
timestamp 1676037725
transform 1 0 25024 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_267
timestamp 1676037725
transform 1 0 25668 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_279
timestamp 1676037725
transform 1 0 26772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_287
timestamp 1676037725
transform 1 0 27508 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_292
timestamp 1676037725
transform 1 0 27968 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_298
timestamp 1676037725
transform 1 0 28520 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1676037725
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_318
timestamp 1676037725
transform 1 0 30360 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_330
timestamp 1676037725
transform 1 0 31464 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_342
timestamp 1676037725
transform 1 0 32568 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_346
timestamp 1676037725
transform 1 0 32936 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_354
timestamp 1676037725
transform 1 0 33672 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1676037725
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_375
timestamp 1676037725
transform 1 0 35604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_387
timestamp 1676037725
transform 1 0 36708 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_405
timestamp 1676037725
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_77
timestamp 1676037725
transform 1 0 8188 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_88
timestamp 1676037725
transform 1 0 9200 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_96
timestamp 1676037725
transform 1 0 9936 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_103
timestamp 1676037725
transform 1 0 10580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_122
timestamp 1676037725
transform 1 0 12328 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_130
timestamp 1676037725
transform 1 0 13064 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_138
timestamp 1676037725
transform 1 0 13800 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_150
timestamp 1676037725
transform 1 0 14904 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_156
timestamp 1676037725
transform 1 0 15456 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_179
timestamp 1676037725
transform 1 0 17572 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_189
timestamp 1676037725
transform 1 0 18492 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_193
timestamp 1676037725
transform 1 0 18860 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_202
timestamp 1676037725
transform 1 0 19688 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1676037725
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_235
timestamp 1676037725
transform 1 0 22724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_247
timestamp 1676037725
transform 1 0 23828 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_255
timestamp 1676037725
transform 1 0 24564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_263
timestamp 1676037725
transform 1 0 25300 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_272
timestamp 1676037725
transform 1 0 26128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_287
timestamp 1676037725
transform 1 0 27508 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_295
timestamp 1676037725
transform 1 0 28244 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_307
timestamp 1676037725
transform 1 0 29348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_319
timestamp 1676037725
transform 1 0 30452 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_333
timestamp 1676037725
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_349
timestamp 1676037725
transform 1 0 33212 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_355
timestamp 1676037725
transform 1 0 33764 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_367
timestamp 1676037725
transform 1 0 34868 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_379
timestamp 1676037725
transform 1 0 35972 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1676037725
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1676037725
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_78
timestamp 1676037725
transform 1 0 8280 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_93
timestamp 1676037725
transform 1 0 9660 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_110
timestamp 1676037725
transform 1 0 11224 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_122
timestamp 1676037725
transform 1 0 12328 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_134
timestamp 1676037725
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_166
timestamp 1676037725
transform 1 0 16376 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_178
timestamp 1676037725
transform 1 0 17480 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1676037725
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_209
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_215
timestamp 1676037725
transform 1 0 20884 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_233
timestamp 1676037725
transform 1 0 22540 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_244
timestamp 1676037725
transform 1 0 23552 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_262
timestamp 1676037725
transform 1 0 25208 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_268
timestamp 1676037725
transform 1 0 25760 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_273
timestamp 1676037725
transform 1 0 26220 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_284
timestamp 1676037725
transform 1 0 27232 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_292
timestamp 1676037725
transform 1 0 27968 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_299
timestamp 1676037725
transform 1 0 28612 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1676037725
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_314
timestamp 1676037725
transform 1 0 29992 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_335
timestamp 1676037725
transform 1 0 31924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_343
timestamp 1676037725
transform 1 0 32660 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_352
timestamp 1676037725
transform 1 0 33488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1676037725
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_385
timestamp 1676037725
transform 1 0 36524 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_397
timestamp 1676037725
transform 1 0 37628 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_405
timestamp 1676037725
transform 1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_68
timestamp 1676037725
transform 1 0 7360 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_80
timestamp 1676037725
transform 1 0 8464 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_92
timestamp 1676037725
transform 1 0 9568 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_104
timestamp 1676037725
transform 1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1676037725
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_136
timestamp 1676037725
transform 1 0 13616 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1676037725
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1676037725
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_183
timestamp 1676037725
transform 1 0 17940 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_191
timestamp 1676037725
transform 1 0 18676 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1676037725
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1676037725
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_233
timestamp 1676037725
transform 1 0 22540 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_240
timestamp 1676037725
transform 1 0 23184 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_252
timestamp 1676037725
transform 1 0 24288 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_256
timestamp 1676037725
transform 1 0 24656 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_266
timestamp 1676037725
transform 1 0 25576 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1676037725
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_291
timestamp 1676037725
transform 1 0 27876 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_299
timestamp 1676037725
transform 1 0 28612 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_310
timestamp 1676037725
transform 1 0 29624 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_318
timestamp 1676037725
transform 1 0 30360 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_327
timestamp 1676037725
transform 1 0 31188 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1676037725
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_346
timestamp 1676037725
transform 1 0 32936 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_358
timestamp 1676037725
transform 1 0 34040 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_370
timestamp 1676037725
transform 1 0 35144 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_381
timestamp 1676037725
transform 1 0 36156 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_389
timestamp 1676037725
transform 1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_404
timestamp 1676037725
transform 1 0 38272 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_73
timestamp 1676037725
transform 1 0 7820 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_78
timestamp 1676037725
transform 1 0 8280 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_103
timestamp 1676037725
transform 1 0 10580 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_111
timestamp 1676037725
transform 1 0 11316 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_120
timestamp 1676037725
transform 1 0 12144 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_135
timestamp 1676037725
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_160
timestamp 1676037725
transform 1 0 15824 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_180
timestamp 1676037725
transform 1 0 17664 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1676037725
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_221
timestamp 1676037725
transform 1 0 21436 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_229
timestamp 1676037725
transform 1 0 22172 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_238
timestamp 1676037725
transform 1 0 23000 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_265
timestamp 1676037725
transform 1 0 25484 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_273
timestamp 1676037725
transform 1 0 26220 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_283
timestamp 1676037725
transform 1 0 27140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_295
timestamp 1676037725
transform 1 0 28244 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1676037725
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_321
timestamp 1676037725
transform 1 0 30636 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_330
timestamp 1676037725
transform 1 0 31464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_342
timestamp 1676037725
transform 1 0 32568 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_350
timestamp 1676037725
transform 1 0 33304 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_359
timestamp 1676037725
transform 1 0 34132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1676037725
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_377
timestamp 1676037725
transform 1 0 35788 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_385
timestamp 1676037725
transform 1 0 36524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_405
timestamp 1676037725
transform 1 0 38364 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_75
timestamp 1676037725
transform 1 0 8004 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_83
timestamp 1676037725
transform 1 0 8740 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_95
timestamp 1676037725
transform 1 0 9844 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1676037725
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_132
timestamp 1676037725
transform 1 0 13248 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_144
timestamp 1676037725
transform 1 0 14352 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_151
timestamp 1676037725
transform 1 0 14996 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_155
timestamp 1676037725
transform 1 0 15364 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_162
timestamp 1676037725
transform 1 0 16008 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_181
timestamp 1676037725
transform 1 0 17756 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_185
timestamp 1676037725
transform 1 0 18124 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_202
timestamp 1676037725
transform 1 0 19688 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_214
timestamp 1676037725
transform 1 0 20792 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_238
timestamp 1676037725
transform 1 0 23000 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_247
timestamp 1676037725
transform 1 0 23828 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_251
timestamp 1676037725
transform 1 0 24196 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_259
timestamp 1676037725
transform 1 0 24932 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1676037725
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_290
timestamp 1676037725
transform 1 0 27784 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_301
timestamp 1676037725
transform 1 0 28796 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_309
timestamp 1676037725
transform 1 0 29532 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_319
timestamp 1676037725
transform 1 0 30452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_331
timestamp 1676037725
transform 1 0 31556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1676037725
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_356
timestamp 1676037725
transform 1 0 33856 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_368
timestamp 1676037725
transform 1 0 34960 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_377
timestamp 1676037725
transform 1 0 35788 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_388
timestamp 1676037725
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_404
timestamp 1676037725
transform 1 0 38272 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_49
timestamp 1676037725
transform 1 0 5612 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_67
timestamp 1676037725
transform 1 0 7268 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_79
timestamp 1676037725
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_113
timestamp 1676037725
transform 1 0 11500 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_131
timestamp 1676037725
transform 1 0 13156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_155
timestamp 1676037725
transform 1 0 15364 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_172
timestamp 1676037725
transform 1 0 16928 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_184
timestamp 1676037725
transform 1 0 18032 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_204
timestamp 1676037725
transform 1 0 19872 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_216
timestamp 1676037725
transform 1 0 20976 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_227
timestamp 1676037725
transform 1 0 21988 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_235
timestamp 1676037725
transform 1 0 22724 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_241
timestamp 1676037725
transform 1 0 23276 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_271
timestamp 1676037725
transform 1 0 26036 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_279
timestamp 1676037725
transform 1 0 26772 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_290
timestamp 1676037725
transform 1 0 27784 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_302
timestamp 1676037725
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_319
timestamp 1676037725
transform 1 0 30452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_330
timestamp 1676037725
transform 1 0 31464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_341
timestamp 1676037725
transform 1 0 32476 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_347
timestamp 1676037725
transform 1 0 33028 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_355
timestamp 1676037725
transform 1 0 33764 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1676037725
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1676037725
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_389
timestamp 1676037725
transform 1 0 36892 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_397
timestamp 1676037725
transform 1 0 37628 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_405
timestamp 1676037725
transform 1 0 38364 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_61
timestamp 1676037725
transform 1 0 6716 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_65
timestamp 1676037725
transform 1 0 7084 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_73
timestamp 1676037725
transform 1 0 7820 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_90
timestamp 1676037725
transform 1 0 9384 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_96
timestamp 1676037725
transform 1 0 9936 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_104
timestamp 1676037725
transform 1 0 10672 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_135
timestamp 1676037725
transform 1 0 13524 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_148
timestamp 1676037725
transform 1 0 14720 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_158
timestamp 1676037725
transform 1 0 15640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1676037725
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1676037725
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_184
timestamp 1676037725
transform 1 0 18032 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_194
timestamp 1676037725
transform 1 0 18952 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_207
timestamp 1676037725
transform 1 0 20148 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1676037725
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1676037725
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_233
timestamp 1676037725
transform 1 0 22540 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_241
timestamp 1676037725
transform 1 0 23276 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_253
timestamp 1676037725
transform 1 0 24380 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_268
timestamp 1676037725
transform 1 0 25760 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_293
timestamp 1676037725
transform 1 0 28060 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_301
timestamp 1676037725
transform 1 0 28796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_310
timestamp 1676037725
transform 1 0 29624 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_318
timestamp 1676037725
transform 1 0 30360 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_327
timestamp 1676037725
transform 1 0 31188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1676037725
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_349
timestamp 1676037725
transform 1 0 33212 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_355
timestamp 1676037725
transform 1 0 33764 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_367
timestamp 1676037725
transform 1 0 34868 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_373
timestamp 1676037725
transform 1 0 35420 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_381
timestamp 1676037725
transform 1 0 36156 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_389
timestamp 1676037725
transform 1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_404
timestamp 1676037725
transform 1 0 38272 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_33
timestamp 1676037725
transform 1 0 4140 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_50
timestamp 1676037725
transform 1 0 5704 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_64
timestamp 1676037725
transform 1 0 6992 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 1676037725
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_89
timestamp 1676037725
transform 1 0 9292 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1676037725
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_135
timestamp 1676037725
transform 1 0 13524 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_146
timestamp 1676037725
transform 1 0 14536 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_157
timestamp 1676037725
transform 1 0 15548 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_169
timestamp 1676037725
transform 1 0 16652 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_179
timestamp 1676037725
transform 1 0 17572 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1676037725
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1676037725
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_212
timestamp 1676037725
transform 1 0 20608 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_220
timestamp 1676037725
transform 1 0 21344 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_228
timestamp 1676037725
transform 1 0 22080 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_235
timestamp 1676037725
transform 1 0 22724 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1676037725
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_260
timestamp 1676037725
transform 1 0 25024 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_268
timestamp 1676037725
transform 1 0 25760 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_286
timestamp 1676037725
transform 1 0 27416 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_298
timestamp 1676037725
transform 1 0 28520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1676037725
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_321
timestamp 1676037725
transform 1 0 30636 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_340
timestamp 1676037725
transform 1 0 32384 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_352
timestamp 1676037725
transform 1 0 33488 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_377
timestamp 1676037725
transform 1 0 35788 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_385
timestamp 1676037725
transform 1 0 36524 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_403
timestamp 1676037725
transform 1 0 38180 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1676037725
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_82
timestamp 1676037725
transform 1 0 8648 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_106
timestamp 1676037725
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_121
timestamp 1676037725
transform 1 0 12236 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_133
timestamp 1676037725
transform 1 0 13340 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_145
timestamp 1676037725
transform 1 0 14444 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_153
timestamp 1676037725
transform 1 0 15180 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1676037725
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1676037725
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_183
timestamp 1676037725
transform 1 0 17940 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_194
timestamp 1676037725
transform 1 0 18952 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_207
timestamp 1676037725
transform 1 0 20148 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_216
timestamp 1676037725
transform 1 0 20976 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_245
timestamp 1676037725
transform 1 0 23644 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_260
timestamp 1676037725
transform 1 0 25024 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_268
timestamp 1676037725
transform 1 0 25760 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1676037725
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_292
timestamp 1676037725
transform 1 0 27968 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_308
timestamp 1676037725
transform 1 0 29440 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_320
timestamp 1676037725
transform 1 0 30544 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1676037725
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1676037725
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_361
timestamp 1676037725
transform 1 0 34316 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_375
timestamp 1676037725
transform 1 0 35604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_387
timestamp 1676037725
transform 1 0 36708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1676037725
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1676037725
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_47
timestamp 1676037725
transform 1 0 5428 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_66
timestamp 1676037725
transform 1 0 7176 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1676037725
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_106
timestamp 1676037725
transform 1 0 10856 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_126
timestamp 1676037725
transform 1 0 12696 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_149
timestamp 1676037725
transform 1 0 14812 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_159
timestamp 1676037725
transform 1 0 15732 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_167
timestamp 1676037725
transform 1 0 16468 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_174
timestamp 1676037725
transform 1 0 17112 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_207
timestamp 1676037725
transform 1 0 20148 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_220
timestamp 1676037725
transform 1 0 21344 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_226
timestamp 1676037725
transform 1 0 21896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_235
timestamp 1676037725
transform 1 0 22724 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_247
timestamp 1676037725
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1676037725
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_260
timestamp 1676037725
transform 1 0 25024 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_272
timestamp 1676037725
transform 1 0 26128 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_280
timestamp 1676037725
transform 1 0 26864 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1676037725
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1676037725
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1676037725
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_317
timestamp 1676037725
transform 1 0 30268 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_332
timestamp 1676037725
transform 1 0 31648 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_344
timestamp 1676037725
transform 1 0 32752 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_353
timestamp 1676037725
transform 1 0 33580 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_361
timestamp 1676037725
transform 1 0 34316 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_384
timestamp 1676037725
transform 1 0 36432 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_396
timestamp 1676037725
transform 1 0 37536 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_405
timestamp 1676037725
transform 1 0 38364 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_27
timestamp 1676037725
transform 1 0 3588 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_76
timestamp 1676037725
transform 1 0 8096 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_88
timestamp 1676037725
transform 1 0 9200 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_97
timestamp 1676037725
transform 1 0 10028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp 1676037725
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_119
timestamp 1676037725
transform 1 0 12052 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_137
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_150
timestamp 1676037725
transform 1 0 14904 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_181
timestamp 1676037725
transform 1 0 17756 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_192
timestamp 1676037725
transform 1 0 18768 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_198
timestamp 1676037725
transform 1 0 19320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_215
timestamp 1676037725
transform 1 0 20884 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_243
timestamp 1676037725
transform 1 0 23460 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_254
timestamp 1676037725
transform 1 0 24472 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_264
timestamp 1676037725
transform 1 0 25392 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_268
timestamp 1676037725
transform 1 0 25760 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1676037725
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_289
timestamp 1676037725
transform 1 0 27692 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_298
timestamp 1676037725
transform 1 0 28520 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_312
timestamp 1676037725
transform 1 0 29808 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_328
timestamp 1676037725
transform 1 0 31280 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_349
timestamp 1676037725
transform 1 0 33212 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_358
timestamp 1676037725
transform 1 0 34040 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_370
timestamp 1676037725
transform 1 0 35144 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_379
timestamp 1676037725
transform 1 0 35972 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1676037725
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_404
timestamp 1676037725
transform 1 0 38272 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_59
timestamp 1676037725
transform 1 0 6532 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_66
timestamp 1676037725
transform 1 0 7176 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_78
timestamp 1676037725
transform 1 0 8280 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1676037725
transform 1 0 9476 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_108
timestamp 1676037725
transform 1 0 11040 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_120
timestamp 1676037725
transform 1 0 12144 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_132
timestamp 1676037725
transform 1 0 13248 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_152
timestamp 1676037725
transform 1 0 15088 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_162
timestamp 1676037725
transform 1 0 16008 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_170
timestamp 1676037725
transform 1 0 16744 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_191
timestamp 1676037725
transform 1 0 18676 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1676037725
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_209
timestamp 1676037725
transform 1 0 20332 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_231
timestamp 1676037725
transform 1 0 22356 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_243
timestamp 1676037725
transform 1 0 23460 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1676037725
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_273
timestamp 1676037725
transform 1 0 26220 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1676037725
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1676037725
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1676037725
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_314
timestamp 1676037725
transform 1 0 29992 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_326
timestamp 1676037725
transform 1 0 31096 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_337
timestamp 1676037725
transform 1 0 32108 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_341
timestamp 1676037725
transform 1 0 32476 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_346
timestamp 1676037725
transform 1 0 32936 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_358
timestamp 1676037725
transform 1 0 34040 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_377
timestamp 1676037725
transform 1 0 35788 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_385
timestamp 1676037725
transform 1 0 36524 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_403
timestamp 1676037725
transform 1 0 38180 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_35
timestamp 1676037725
transform 1 0 4324 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_47
timestamp 1676037725
transform 1 0 5428 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1676037725
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_66
timestamp 1676037725
transform 1 0 7176 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_70
timestamp 1676037725
transform 1 0 7544 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_78
timestamp 1676037725
transform 1 0 8280 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_91
timestamp 1676037725
transform 1 0 9476 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_99
timestamp 1676037725
transform 1 0 10212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1676037725
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_137
timestamp 1676037725
transform 1 0 13708 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_145
timestamp 1676037725
transform 1 0 14444 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_154
timestamp 1676037725
transform 1 0 15272 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_182
timestamp 1676037725
transform 1 0 17848 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_194
timestamp 1676037725
transform 1 0 18952 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_206
timestamp 1676037725
transform 1 0 20056 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_218
timestamp 1676037725
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_235
timestamp 1676037725
transform 1 0 22724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_247
timestamp 1676037725
transform 1 0 23828 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_255
timestamp 1676037725
transform 1 0 24564 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_262
timestamp 1676037725
transform 1 0 25208 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_270
timestamp 1676037725
transform 1 0 25944 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1676037725
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_290
timestamp 1676037725
transform 1 0 27784 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_304
timestamp 1676037725
transform 1 0 29072 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_316
timestamp 1676037725
transform 1 0 30176 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_334
timestamp 1676037725
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_347
timestamp 1676037725
transform 1 0 33028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_359
timestamp 1676037725
transform 1 0 34132 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_367
timestamp 1676037725
transform 1 0 34868 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_376
timestamp 1676037725
transform 1 0 35696 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_387
timestamp 1676037725
transform 1 0 36708 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1676037725
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_404
timestamp 1676037725
transform 1 0 38272 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_40
timestamp 1676037725
transform 1 0 4784 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_52
timestamp 1676037725
transform 1 0 5888 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_64
timestamp 1676037725
transform 1 0 6992 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_74
timestamp 1676037725
transform 1 0 7912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1676037725
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_92
timestamp 1676037725
transform 1 0 9568 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_100
timestamp 1676037725
transform 1 0 10304 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1676037725
transform 1 0 11960 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1676037725
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_148
timestamp 1676037725
transform 1 0 14720 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_160
timestamp 1676037725
transform 1 0 15824 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_169
timestamp 1676037725
transform 1 0 16652 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_181
timestamp 1676037725
transform 1 0 17756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1676037725
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1676037725
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_233
timestamp 1676037725
transform 1 0 22540 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_242
timestamp 1676037725
transform 1 0 23368 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_246
timestamp 1676037725
transform 1 0 23736 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_270
timestamp 1676037725
transform 1 0 25944 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_278
timestamp 1676037725
transform 1 0 26680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_286
timestamp 1676037725
transform 1 0 27416 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_290
timestamp 1676037725
transform 1 0 27784 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_294
timestamp 1676037725
transform 1 0 28152 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1676037725
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_329
timestamp 1676037725
transform 1 0 31372 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_341
timestamp 1676037725
transform 1 0 32476 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_350
timestamp 1676037725
transform 1 0 33304 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_361
timestamp 1676037725
transform 1 0 34316 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_384
timestamp 1676037725
transform 1 0 36432 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_388
timestamp 1676037725
transform 1 0 36800 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1676037725
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1676037725
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1676037725
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_42
timestamp 1676037725
transform 1 0 4968 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_65
timestamp 1676037725
transform 1 0 7084 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_73
timestamp 1676037725
transform 1 0 7820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_92
timestamp 1676037725
transform 1 0 9568 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1676037725
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_123
timestamp 1676037725
transform 1 0 12420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_135
timestamp 1676037725
transform 1 0 13524 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_143
timestamp 1676037725
transform 1 0 14260 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_147
timestamp 1676037725
transform 1 0 14628 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_154
timestamp 1676037725
transform 1 0 15272 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_178
timestamp 1676037725
transform 1 0 17480 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_197
timestamp 1676037725
transform 1 0 19228 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1676037725
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_247
timestamp 1676037725
transform 1 0 23828 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_251
timestamp 1676037725
transform 1 0 24196 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_265
timestamp 1676037725
transform 1 0 25484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_277
timestamp 1676037725
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_287
timestamp 1676037725
transform 1 0 27508 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_297
timestamp 1676037725
transform 1 0 28428 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_305
timestamp 1676037725
transform 1 0 29164 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_314
timestamp 1676037725
transform 1 0 29992 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_320
timestamp 1676037725
transform 1 0 30544 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1676037725
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_345
timestamp 1676037725
transform 1 0 32844 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_353
timestamp 1676037725
transform 1 0 33580 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_365
timestamp 1676037725
transform 1 0 34684 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_369
timestamp 1676037725
transform 1 0 35052 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_378
timestamp 1676037725
transform 1 0 35880 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_390
timestamp 1676037725
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1676037725
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1676037725
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_40
timestamp 1676037725
transform 1 0 4784 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_66
timestamp 1676037725
transform 1 0 7176 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_76
timestamp 1676037725
transform 1 0 8096 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_104
timestamp 1676037725
transform 1 0 10672 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_116
timestamp 1676037725
transform 1 0 11776 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_135
timestamp 1676037725
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1676037725
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_150
timestamp 1676037725
transform 1 0 14904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_158
timestamp 1676037725
transform 1 0 15640 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_165
timestamp 1676037725
transform 1 0 16284 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_171
timestamp 1676037725
transform 1 0 16836 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_188
timestamp 1676037725
transform 1 0 18400 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_205
timestamp 1676037725
transform 1 0 19964 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_215
timestamp 1676037725
transform 1 0 20884 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_228
timestamp 1676037725
transform 1 0 22080 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_240
timestamp 1676037725
transform 1 0 23184 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_265
timestamp 1676037725
transform 1 0 25484 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_269
timestamp 1676037725
transform 1 0 25852 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_285
timestamp 1676037725
transform 1 0 27324 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_289
timestamp 1676037725
transform 1 0 27692 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_293
timestamp 1676037725
transform 1 0 28060 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_306
timestamp 1676037725
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_325
timestamp 1676037725
transform 1 0 31004 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_337
timestamp 1676037725
transform 1 0 32108 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_349
timestamp 1676037725
transform 1 0 33212 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_361
timestamp 1676037725
transform 1 0 34316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_376
timestamp 1676037725
transform 1 0 35696 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_384
timestamp 1676037725
transform 1 0 36432 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_403
timestamp 1676037725
transform 1 0 38180 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_33
timestamp 1676037725
transform 1 0 4140 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_44
timestamp 1676037725
transform 1 0 5152 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1676037725
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_77
timestamp 1676037725
transform 1 0 8188 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_82
timestamp 1676037725
transform 1 0 8648 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_88
timestamp 1676037725
transform 1 0 9200 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_95
timestamp 1676037725
transform 1 0 9844 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_104
timestamp 1676037725
transform 1 0 10672 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1676037725
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1676037725
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1676037725
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1676037725
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1676037725
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1676037725
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_193
timestamp 1676037725
transform 1 0 18860 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_201
timestamp 1676037725
transform 1 0 19596 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_207
timestamp 1676037725
transform 1 0 20148 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_211
timestamp 1676037725
transform 1 0 20516 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1676037725
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_250
timestamp 1676037725
transform 1 0 24104 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_263
timestamp 1676037725
transform 1 0 25300 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1676037725
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_289
timestamp 1676037725
transform 1 0 27692 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_295
timestamp 1676037725
transform 1 0 28244 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_303
timestamp 1676037725
transform 1 0 28980 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_311
timestamp 1676037725
transform 1 0 29716 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_322
timestamp 1676037725
transform 1 0 30728 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1676037725
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_347
timestamp 1676037725
transform 1 0 33028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_359
timestamp 1676037725
transform 1 0 34132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_365
timestamp 1676037725
transform 1 0 34684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_374
timestamp 1676037725
transform 1 0 35512 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1676037725
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1676037725
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_404
timestamp 1676037725
transform 1 0 38272 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1676037725
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1676037725
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_53
timestamp 1676037725
transform 1 0 5980 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_66
timestamp 1676037725
transform 1 0 7176 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_81
timestamp 1676037725
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_95
timestamp 1676037725
transform 1 0 9844 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_103
timestamp 1676037725
transform 1 0 10580 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_120
timestamp 1676037725
transform 1 0 12144 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_132
timestamp 1676037725
transform 1 0 13248 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_159
timestamp 1676037725
transform 1 0 15732 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_167
timestamp 1676037725
transform 1 0 16468 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_187
timestamp 1676037725
transform 1 0 18308 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_210
timestamp 1676037725
transform 1 0 20424 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1676037725
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_243
timestamp 1676037725
transform 1 0 23460 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_260
timestamp 1676037725
transform 1 0 25024 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_268
timestamp 1676037725
transform 1 0 25760 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_277
timestamp 1676037725
transform 1 0 26588 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_283
timestamp 1676037725
transform 1 0 27140 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_292
timestamp 1676037725
transform 1 0 27968 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1676037725
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_322
timestamp 1676037725
transform 1 0 30728 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_342
timestamp 1676037725
transform 1 0 32568 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_354
timestamp 1676037725
transform 1 0 33672 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1676037725
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1676037725
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_389
timestamp 1676037725
transform 1 0 36892 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_397
timestamp 1676037725
transform 1 0 37628 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1676037725
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_15
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_33
timestamp 1676037725
transform 1 0 4140 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_46
timestamp 1676037725
transform 1 0 5336 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_50
timestamp 1676037725
transform 1 0 5704 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1676037725
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_64
timestamp 1676037725
transform 1 0 6992 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_75
timestamp 1676037725
transform 1 0 8004 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_87
timestamp 1676037725
transform 1 0 9108 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_91
timestamp 1676037725
transform 1 0 9476 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_98
timestamp 1676037725
transform 1 0 10120 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_109
timestamp 1676037725
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1676037725
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_137
timestamp 1676037725
transform 1 0 13708 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_160
timestamp 1676037725
transform 1 0 15824 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_190
timestamp 1676037725
transform 1 0 18584 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_202
timestamp 1676037725
transform 1 0 19688 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1676037725
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_239
timestamp 1676037725
transform 1 0 23092 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_243
timestamp 1676037725
transform 1 0 23460 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_253
timestamp 1676037725
transform 1 0 24380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1676037725
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1676037725
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_287
timestamp 1676037725
transform 1 0 27508 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_299
timestamp 1676037725
transform 1 0 28612 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_307
timestamp 1676037725
transform 1 0 29348 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_320
timestamp 1676037725
transform 1 0 30544 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_332
timestamp 1676037725
transform 1 0 31648 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_337
timestamp 1676037725
transform 1 0 32108 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_347
timestamp 1676037725
transform 1 0 33028 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_351
timestamp 1676037725
transform 1 0 33396 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_357
timestamp 1676037725
transform 1 0 33948 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_365
timestamp 1676037725
transform 1 0 34684 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_382
timestamp 1676037725
transform 1 0 36248 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_390
timestamp 1676037725
transform 1 0 36984 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_393
timestamp 1676037725
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_404
timestamp 1676037725
transform 1 0 38272 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_37
timestamp 1676037725
transform 1 0 4508 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_49
timestamp 1676037725
transform 1 0 5612 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_55
timestamp 1676037725
transform 1 0 6164 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_63
timestamp 1676037725
transform 1 0 6900 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_71
timestamp 1676037725
transform 1 0 7636 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1676037725
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_93
timestamp 1676037725
transform 1 0 9660 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_101
timestamp 1676037725
transform 1 0 10396 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_109
timestamp 1676037725
transform 1 0 11132 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_129
timestamp 1676037725
transform 1 0 12972 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_137
timestamp 1676037725
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_150
timestamp 1676037725
transform 1 0 14904 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_162
timestamp 1676037725
transform 1 0 16008 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_175
timestamp 1676037725
transform 1 0 17204 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1676037725
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_204
timestamp 1676037725
transform 1 0 19872 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_219
timestamp 1676037725
transform 1 0 21252 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_230
timestamp 1676037725
transform 1 0 22264 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_234
timestamp 1676037725
transform 1 0 22632 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_240
timestamp 1676037725
transform 1 0 23184 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_266
timestamp 1676037725
transform 1 0 25576 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_283
timestamp 1676037725
transform 1 0 27140 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_290
timestamp 1676037725
transform 1 0 27784 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_302
timestamp 1676037725
transform 1 0 28888 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_309
timestamp 1676037725
transform 1 0 29532 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_313
timestamp 1676037725
transform 1 0 29900 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_330
timestamp 1676037725
transform 1 0 31464 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_338
timestamp 1676037725
transform 1 0 32200 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_347
timestamp 1676037725
transform 1 0 33028 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1676037725
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_365
timestamp 1676037725
transform 1 0 34684 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_384
timestamp 1676037725
transform 1 0 36432 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_404
timestamp 1676037725
transform 1 0 38272 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1676037725
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_39
timestamp 1676037725
transform 1 0 4692 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_49
timestamp 1676037725
transform 1 0 5612 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_63
timestamp 1676037725
transform 1 0 6900 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_71
timestamp 1676037725
transform 1 0 7636 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_78
timestamp 1676037725
transform 1 0 8280 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_90
timestamp 1676037725
transform 1 0 9384 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_101
timestamp 1676037725
transform 1 0 10396 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_109
timestamp 1676037725
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_125
timestamp 1676037725
transform 1 0 12604 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_147
timestamp 1676037725
transform 1 0 14628 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_159
timestamp 1676037725
transform 1 0 15732 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1676037725
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_177
timestamp 1676037725
transform 1 0 17388 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_183
timestamp 1676037725
transform 1 0 17940 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_193
timestamp 1676037725
transform 1 0 18860 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_208
timestamp 1676037725
transform 1 0 20240 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_219
timestamp 1676037725
transform 1 0 21252 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1676037725
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_231
timestamp 1676037725
transform 1 0 22356 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_248
timestamp 1676037725
transform 1 0 23920 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_262
timestamp 1676037725
transform 1 0 25208 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_274
timestamp 1676037725
transform 1 0 26312 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_294
timestamp 1676037725
transform 1 0 28152 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_314
timestamp 1676037725
transform 1 0 29992 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_333
timestamp 1676037725
transform 1 0 31740 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_337
timestamp 1676037725
transform 1 0 32108 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_345
timestamp 1676037725
transform 1 0 32844 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_351
timestamp 1676037725
transform 1 0 33396 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_363
timestamp 1676037725
transform 1 0 34500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_375
timestamp 1676037725
transform 1 0 35604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_387
timestamp 1676037725
transform 1 0 36708 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1676037725
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_393
timestamp 1676037725
transform 1 0 37260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1676037725
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_33
timestamp 1676037725
transform 1 0 4140 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_37
timestamp 1676037725
transform 1 0 4508 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_48
timestamp 1676037725
transform 1 0 5520 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_52
timestamp 1676037725
transform 1 0 5888 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_57
timestamp 1676037725
transform 1 0 6348 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_64
timestamp 1676037725
transform 1 0 6992 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_76
timestamp 1676037725
transform 1 0 8096 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_95
timestamp 1676037725
transform 1 0 9844 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_119
timestamp 1676037725
transform 1 0 12052 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_131
timestamp 1676037725
transform 1 0 13156 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1676037725
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_149
timestamp 1676037725
transform 1 0 14812 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_164
timestamp 1676037725
transform 1 0 16192 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_185
timestamp 1676037725
transform 1 0 18124 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_193
timestamp 1676037725
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_209
timestamp 1676037725
transform 1 0 20332 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_215
timestamp 1676037725
transform 1 0 20884 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_225
timestamp 1676037725
transform 1 0 21804 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_229
timestamp 1676037725
transform 1 0 22172 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_236
timestamp 1676037725
transform 1 0 22816 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1676037725
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1676037725
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_264
timestamp 1676037725
transform 1 0 25392 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_273
timestamp 1676037725
transform 1 0 26220 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_281
timestamp 1676037725
transform 1 0 26956 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_288
timestamp 1676037725
transform 1 0 27600 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_299
timestamp 1676037725
transform 1 0 28612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1676037725
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_309
timestamp 1676037725
transform 1 0 29532 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_317
timestamp 1676037725
transform 1 0 30268 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_329
timestamp 1676037725
transform 1 0 31372 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_342
timestamp 1676037725
transform 1 0 32568 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_353
timestamp 1676037725
transform 1 0 33580 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1676037725
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_365
timestamp 1676037725
transform 1 0 34684 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_378
timestamp 1676037725
transform 1 0 35880 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_386
timestamp 1676037725
transform 1 0 36616 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_404
timestamp 1676037725
transform 1 0 38272 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_15
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_34
timestamp 1676037725
transform 1 0 4232 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_42
timestamp 1676037725
transform 1 0 4968 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1676037725
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_61
timestamp 1676037725
transform 1 0 6716 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_68
timestamp 1676037725
transform 1 0 7360 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_76
timestamp 1676037725
transform 1 0 8096 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_84
timestamp 1676037725
transform 1 0 8832 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_91
timestamp 1676037725
transform 1 0 9476 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_99
timestamp 1676037725
transform 1 0 10212 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1676037725
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_125
timestamp 1676037725
transform 1 0 12604 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_137
timestamp 1676037725
transform 1 0 13708 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_143
timestamp 1676037725
transform 1 0 14260 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_150
timestamp 1676037725
transform 1 0 14904 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_162
timestamp 1676037725
transform 1 0 16008 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_178
timestamp 1676037725
transform 1 0 17480 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_187
timestamp 1676037725
transform 1 0 18308 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_198
timestamp 1676037725
transform 1 0 19320 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_204
timestamp 1676037725
transform 1 0 19872 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_208
timestamp 1676037725
transform 1 0 20240 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_219
timestamp 1676037725
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1676037725
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_233
timestamp 1676037725
transform 1 0 22540 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_243
timestamp 1676037725
transform 1 0 23460 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_258
timestamp 1676037725
transform 1 0 24840 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_270
timestamp 1676037725
transform 1 0 25944 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1676037725
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_299
timestamp 1676037725
transform 1 0 28612 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_319
timestamp 1676037725
transform 1 0 30452 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_330
timestamp 1676037725
transform 1 0 31464 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_337
timestamp 1676037725
transform 1 0 32108 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_45_360
timestamp 1676037725
transform 1 0 34224 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_368
timestamp 1676037725
transform 1 0 34960 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_377
timestamp 1676037725
transform 1 0 35788 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_387
timestamp 1676037725
transform 1 0 36708 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1676037725
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1676037725
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_404
timestamp 1676037725
transform 1 0 38272 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1676037725
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_39
timestamp 1676037725
transform 1 0 4692 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_52
timestamp 1676037725
transform 1 0 5888 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_60
timestamp 1676037725
transform 1 0 6624 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_66
timestamp 1676037725
transform 1 0 7176 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_72
timestamp 1676037725
transform 1 0 7728 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1676037725
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_91
timestamp 1676037725
transform 1 0 9476 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_105
timestamp 1676037725
transform 1 0 10764 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_112
timestamp 1676037725
transform 1 0 11408 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_124
timestamp 1676037725
transform 1 0 12512 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_130
timestamp 1676037725
transform 1 0 13064 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1676037725
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_159
timestamp 1676037725
transform 1 0 15732 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_171
timestamp 1676037725
transform 1 0 16836 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_188
timestamp 1676037725
transform 1 0 18400 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_215
timestamp 1676037725
transform 1 0 20884 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_225
timestamp 1676037725
transform 1 0 21804 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_233
timestamp 1676037725
transform 1 0 22540 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1676037725
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_265
timestamp 1676037725
transform 1 0 25484 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_281
timestamp 1676037725
transform 1 0 26956 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_293
timestamp 1676037725
transform 1 0 28060 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_306
timestamp 1676037725
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1676037725
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_319
timestamp 1676037725
transform 1 0 30452 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_331
timestamp 1676037725
transform 1 0 31556 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_342
timestamp 1676037725
transform 1 0 32568 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_349
timestamp 1676037725
transform 1 0 33212 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_361
timestamp 1676037725
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1676037725
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1676037725
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_395
timestamp 1676037725
transform 1 0 37444 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1676037725
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1676037725
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_39
timestamp 1676037725
transform 1 0 4692 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_47
timestamp 1676037725
transform 1 0 5428 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_70
timestamp 1676037725
transform 1 0 7544 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_83
timestamp 1676037725
transform 1 0 8740 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_92
timestamp 1676037725
transform 1 0 9568 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_102
timestamp 1676037725
transform 1 0 10488 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_106
timestamp 1676037725
transform 1 0 10856 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1676037725
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_119
timestamp 1676037725
transform 1 0 12052 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_136
timestamp 1676037725
transform 1 0 13616 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_147
timestamp 1676037725
transform 1 0 14628 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_159
timestamp 1676037725
transform 1 0 15732 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1676037725
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_174
timestamp 1676037725
transform 1 0 17112 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_186
timestamp 1676037725
transform 1 0 18216 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_192
timestamp 1676037725
transform 1 0 18768 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_198
timestamp 1676037725
transform 1 0 19320 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_211
timestamp 1676037725
transform 1 0 20516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1676037725
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_235
timestamp 1676037725
transform 1 0 22724 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_243
timestamp 1676037725
transform 1 0 23460 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_251
timestamp 1676037725
transform 1 0 24196 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_261
timestamp 1676037725
transform 1 0 25116 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_270
timestamp 1676037725
transform 1 0 25944 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1676037725
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_291
timestamp 1676037725
transform 1 0 27876 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_303
timestamp 1676037725
transform 1 0 28980 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_323
timestamp 1676037725
transform 1 0 30820 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1676037725
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1676037725
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_349
timestamp 1676037725
transform 1 0 33212 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_355
timestamp 1676037725
transform 1 0 33764 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_373
timestamp 1676037725
transform 1 0 35420 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_379
timestamp 1676037725
transform 1 0 35972 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_384
timestamp 1676037725
transform 1 0 36432 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_393
timestamp 1676037725
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_404
timestamp 1676037725
transform 1 0 38272 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_40
timestamp 1676037725
transform 1 0 4784 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_51
timestamp 1676037725
transform 1 0 5796 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_59
timestamp 1676037725
transform 1 0 6532 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1676037725
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_96
timestamp 1676037725
transform 1 0 9936 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_104
timestamp 1676037725
transform 1 0 10672 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_112
timestamp 1676037725
transform 1 0 11408 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_122
timestamp 1676037725
transform 1 0 12328 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_129
timestamp 1676037725
transform 1 0 12972 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_137
timestamp 1676037725
transform 1 0 13708 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_150
timestamp 1676037725
transform 1 0 14904 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_162
timestamp 1676037725
transform 1 0 16008 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_171
timestamp 1676037725
transform 1 0 16836 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_179
timestamp 1676037725
transform 1 0 17572 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_184
timestamp 1676037725
transform 1 0 18032 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_207
timestamp 1676037725
transform 1 0 20148 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_215
timestamp 1676037725
transform 1 0 20884 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_224
timestamp 1676037725
transform 1 0 21712 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_232
timestamp 1676037725
transform 1 0 22448 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1676037725
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1676037725
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_266
timestamp 1676037725
transform 1 0 25576 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_278
timestamp 1676037725
transform 1 0 26680 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_288
timestamp 1676037725
transform 1 0 27600 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_299
timestamp 1676037725
transform 1 0 28612 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1676037725
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_309
timestamp 1676037725
transform 1 0 29532 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_324
timestamp 1676037725
transform 1 0 30912 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_337
timestamp 1676037725
transform 1 0 32108 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_341
timestamp 1676037725
transform 1 0 32476 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_349
timestamp 1676037725
transform 1 0 33212 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_361
timestamp 1676037725
transform 1 0 34316 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_365
timestamp 1676037725
transform 1 0 34684 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_378
timestamp 1676037725
transform 1 0 35880 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_386
timestamp 1676037725
transform 1 0 36616 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_405
timestamp 1676037725
transform 1 0 38364 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_31
timestamp 1676037725
transform 1 0 3956 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_48
timestamp 1676037725
transform 1 0 5520 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_65
timestamp 1676037725
transform 1 0 7084 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_75
timestamp 1676037725
transform 1 0 8004 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_83
timestamp 1676037725
transform 1 0 8740 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_91
timestamp 1676037725
transform 1 0 9476 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_104
timestamp 1676037725
transform 1 0 10672 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_118
timestamp 1676037725
transform 1 0 11960 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_126
timestamp 1676037725
transform 1 0 12696 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_132
timestamp 1676037725
transform 1 0 13248 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_147
timestamp 1676037725
transform 1 0 14628 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_159
timestamp 1676037725
transform 1 0 15732 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1676037725
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_178
timestamp 1676037725
transform 1 0 17480 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_182
timestamp 1676037725
transform 1 0 17848 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_194
timestamp 1676037725
transform 1 0 18952 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_203
timestamp 1676037725
transform 1 0 19780 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_216
timestamp 1676037725
transform 1 0 20976 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_238
timestamp 1676037725
transform 1 0 23000 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_249
timestamp 1676037725
transform 1 0 24012 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_257
timestamp 1676037725
transform 1 0 24748 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_266
timestamp 1676037725
transform 1 0 25576 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_275
timestamp 1676037725
transform 1 0 26404 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1676037725
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_290
timestamp 1676037725
transform 1 0 27784 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_301
timestamp 1676037725
transform 1 0 28796 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_314
timestamp 1676037725
transform 1 0 29992 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_327
timestamp 1676037725
transform 1 0 31188 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1676037725
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_337
timestamp 1676037725
transform 1 0 32108 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_345
timestamp 1676037725
transform 1 0 32844 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_349
timestamp 1676037725
transform 1 0 33212 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_367
timestamp 1676037725
transform 1 0 34868 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_375
timestamp 1676037725
transform 1 0 35604 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_384
timestamp 1676037725
transform 1 0 36432 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_393
timestamp 1676037725
transform 1 0 37260 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_401
timestamp 1676037725
transform 1 0 37996 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_15
timestamp 1676037725
transform 1 0 2484 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_26
timestamp 1676037725
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_40
timestamp 1676037725
transform 1 0 4784 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_50
timestamp 1676037725
transform 1 0 5704 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_57
timestamp 1676037725
transform 1 0 6348 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_63
timestamp 1676037725
transform 1 0 6900 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_74
timestamp 1676037725
transform 1 0 7912 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1676037725
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_107
timestamp 1676037725
transform 1 0 10948 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_111
timestamp 1676037725
transform 1 0 11316 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_119
timestamp 1676037725
transform 1 0 12052 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_128
timestamp 1676037725
transform 1 0 12880 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_135
timestamp 1676037725
transform 1 0 13524 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1676037725
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_154
timestamp 1676037725
transform 1 0 15272 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_163
timestamp 1676037725
transform 1 0 16100 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_167
timestamp 1676037725
transform 1 0 16468 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_171
timestamp 1676037725
transform 1 0 16836 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_175
timestamp 1676037725
transform 1 0 17204 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_182
timestamp 1676037725
transform 1 0 17848 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1676037725
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_205
timestamp 1676037725
transform 1 0 19964 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_214
timestamp 1676037725
transform 1 0 20792 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_222
timestamp 1676037725
transform 1 0 21528 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_228
timestamp 1676037725
transform 1 0 22080 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_237
timestamp 1676037725
transform 1 0 22908 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_244
timestamp 1676037725
transform 1 0 23552 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_258
timestamp 1676037725
transform 1 0 24840 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_266
timestamp 1676037725
transform 1 0 25576 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_273
timestamp 1676037725
transform 1 0 26220 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_279
timestamp 1676037725
transform 1 0 26772 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_287
timestamp 1676037725
transform 1 0 27508 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1676037725
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1676037725
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_309
timestamp 1676037725
transform 1 0 29532 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_320
timestamp 1676037725
transform 1 0 30544 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_324
timestamp 1676037725
transform 1 0 30912 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_336
timestamp 1676037725
transform 1 0 32016 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_344
timestamp 1676037725
transform 1 0 32752 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_351
timestamp 1676037725
transform 1 0 33396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1676037725
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_365
timestamp 1676037725
transform 1 0 34684 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_378
timestamp 1676037725
transform 1 0 35880 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_386
timestamp 1676037725
transform 1 0 36616 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_405
timestamp 1676037725
transform 1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_36
timestamp 1676037725
transform 1 0 4416 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_50
timestamp 1676037725
transform 1 0 5704 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_66
timestamp 1676037725
transform 1 0 7176 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_74
timestamp 1676037725
transform 1 0 7912 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_92
timestamp 1676037725
transform 1 0 9568 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_103
timestamp 1676037725
transform 1 0 10580 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1676037725
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_124
timestamp 1676037725
transform 1 0 12512 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_134
timestamp 1676037725
transform 1 0 13432 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_144
timestamp 1676037725
transform 1 0 14352 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_154
timestamp 1676037725
transform 1 0 15272 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_163
timestamp 1676037725
transform 1 0 16100 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1676037725
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_182
timestamp 1676037725
transform 1 0 17848 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_189
timestamp 1676037725
transform 1 0 18492 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_201
timestamp 1676037725
transform 1 0 19596 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_207
timestamp 1676037725
transform 1 0 20148 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_213
timestamp 1676037725
transform 1 0 20700 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_221
timestamp 1676037725
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_233
timestamp 1676037725
transform 1 0 22540 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_243
timestamp 1676037725
transform 1 0 23460 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_251
timestamp 1676037725
transform 1 0 24196 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_257
timestamp 1676037725
transform 1 0 24748 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_263
timestamp 1676037725
transform 1 0 25300 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 1676037725
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_281
timestamp 1676037725
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_292
timestamp 1676037725
transform 1 0 27968 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_305
timestamp 1676037725
transform 1 0 29164 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_51_319
timestamp 1676037725
transform 1 0 30452 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_324
timestamp 1676037725
transform 1 0 30912 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1676037725
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1676037725
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_349
timestamp 1676037725
transform 1 0 33212 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_372
timestamp 1676037725
transform 1 0 35328 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_376
timestamp 1676037725
transform 1 0 35696 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1676037725
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1676037725
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_393
timestamp 1676037725
transform 1 0 37260 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_404
timestamp 1676037725
transform 1 0 38272 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_46
timestamp 1676037725
transform 1 0 5336 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_55
timestamp 1676037725
transform 1 0 6164 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_65
timestamp 1676037725
transform 1 0 7084 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_73
timestamp 1676037725
transform 1 0 7820 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_80
timestamp 1676037725
transform 1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_93
timestamp 1676037725
transform 1 0 9660 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_101
timestamp 1676037725
transform 1 0 10396 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_109
timestamp 1676037725
transform 1 0 11132 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_121
timestamp 1676037725
transform 1 0 12236 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_125
timestamp 1676037725
transform 1 0 12604 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_129
timestamp 1676037725
transform 1 0 12972 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_137
timestamp 1676037725
transform 1 0 13708 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_149
timestamp 1676037725
transform 1 0 14812 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_161
timestamp 1676037725
transform 1 0 15916 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_165
timestamp 1676037725
transform 1 0 16284 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_171
timestamp 1676037725
transform 1 0 16836 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_185
timestamp 1676037725
transform 1 0 18124 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_193
timestamp 1676037725
transform 1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_205
timestamp 1676037725
transform 1 0 19964 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_213
timestamp 1676037725
transform 1 0 20700 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_225
timestamp 1676037725
transform 1 0 21804 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_237
timestamp 1676037725
transform 1 0 22908 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 1676037725
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_265
timestamp 1676037725
transform 1 0 25484 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_274
timestamp 1676037725
transform 1 0 26312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_281
timestamp 1676037725
transform 1 0 26956 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_288
timestamp 1676037725
transform 1 0 27600 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_292
timestamp 1676037725
transform 1 0 27968 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_298
timestamp 1676037725
transform 1 0 28520 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_305
timestamp 1676037725
transform 1 0 29164 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1676037725
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_316
timestamp 1676037725
transform 1 0 30176 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_331
timestamp 1676037725
transform 1 0 31556 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_344
timestamp 1676037725
transform 1 0 32752 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_356
timestamp 1676037725
transform 1 0 33856 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_365
timestamp 1676037725
transform 1 0 34684 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_376
timestamp 1676037725
transform 1 0 35696 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_384
timestamp 1676037725
transform 1 0 36432 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_393
timestamp 1676037725
transform 1 0 37260 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_403
timestamp 1676037725
transform 1 0 38180 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1676037725
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1676037725
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_39
timestamp 1676037725
transform 1 0 4692 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_45
timestamp 1676037725
transform 1 0 5244 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1676037725
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1676037725
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_65
timestamp 1676037725
transform 1 0 7084 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_73
timestamp 1676037725
transform 1 0 7820 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_88
timestamp 1676037725
transform 1 0 9200 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_96
timestamp 1676037725
transform 1 0 9936 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_104
timestamp 1676037725
transform 1 0 10672 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_121
timestamp 1676037725
transform 1 0 12236 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_129
timestamp 1676037725
transform 1 0 12972 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_137
timestamp 1676037725
transform 1 0 13708 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_141
timestamp 1676037725
transform 1 0 14076 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_149
timestamp 1676037725
transform 1 0 14812 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_153
timestamp 1676037725
transform 1 0 15180 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_160
timestamp 1676037725
transform 1 0 15824 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_179
timestamp 1676037725
transform 1 0 17572 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_185
timestamp 1676037725
transform 1 0 18124 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_194
timestamp 1676037725
transform 1 0 18952 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_198
timestamp 1676037725
transform 1 0 19320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_206
timestamp 1676037725
transform 1 0 20056 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_214
timestamp 1676037725
transform 1 0 20792 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_218
timestamp 1676037725
transform 1 0 21160 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1676037725
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_236
timestamp 1676037725
transform 1 0 22816 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_244
timestamp 1676037725
transform 1 0 23552 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_254
timestamp 1676037725
transform 1 0 24472 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_262
timestamp 1676037725
transform 1 0 25208 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_272
timestamp 1676037725
transform 1 0 26128 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_281
timestamp 1676037725
transform 1 0 26956 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_294
timestamp 1676037725
transform 1 0 28152 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_303
timestamp 1676037725
transform 1 0 28980 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_312
timestamp 1676037725
transform 1 0 29808 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_320
timestamp 1676037725
transform 1 0 30544 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1676037725
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1676037725
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_337
timestamp 1676037725
transform 1 0 32108 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_345
timestamp 1676037725
transform 1 0 32844 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_357
timestamp 1676037725
transform 1 0 33948 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_370
timestamp 1676037725
transform 1 0 35144 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_382
timestamp 1676037725
transform 1 0 36248 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_390
timestamp 1676037725
transform 1 0 36984 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_393
timestamp 1676037725
transform 1 0 37260 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_404
timestamp 1676037725
transform 1 0 38272 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_36
timestamp 1676037725
transform 1 0 4416 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_47
timestamp 1676037725
transform 1 0 5428 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_55
timestamp 1676037725
transform 1 0 6164 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_65
timestamp 1676037725
transform 1 0 7084 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_71
timestamp 1676037725
transform 1 0 7636 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_79
timestamp 1676037725
transform 1 0 8372 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1676037725
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_94
timestamp 1676037725
transform 1 0 9752 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_104
timestamp 1676037725
transform 1 0 10672 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_112
timestamp 1676037725
transform 1 0 11408 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_120
timestamp 1676037725
transform 1 0 12144 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_129
timestamp 1676037725
transform 1 0 12972 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_137
timestamp 1676037725
transform 1 0 13708 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_153
timestamp 1676037725
transform 1 0 15180 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_162
timestamp 1676037725
transform 1 0 16008 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_170
timestamp 1676037725
transform 1 0 16744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_179
timestamp 1676037725
transform 1 0 17572 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_187
timestamp 1676037725
transform 1 0 18308 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1676037725
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_204
timestamp 1676037725
transform 1 0 19872 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_216
timestamp 1676037725
transform 1 0 20976 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_226
timestamp 1676037725
transform 1 0 21896 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_234
timestamp 1676037725
transform 1 0 22632 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1676037725
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1676037725
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_262
timestamp 1676037725
transform 1 0 25208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_271
timestamp 1676037725
transform 1 0 26036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_277
timestamp 1676037725
transform 1 0 26588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_284
timestamp 1676037725
transform 1 0 27232 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1676037725
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_309
timestamp 1676037725
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_314
timestamp 1676037725
transform 1 0 29992 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_326
timestamp 1676037725
transform 1 0 31096 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_334
timestamp 1676037725
transform 1 0 31832 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_340
timestamp 1676037725
transform 1 0 32384 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_347
timestamp 1676037725
transform 1 0 33028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_359
timestamp 1676037725
transform 1 0 34132 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1676037725
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_365
timestamp 1676037725
transform 1 0 34684 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_379
timestamp 1676037725
transform 1 0 35972 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_400
timestamp 1676037725
transform 1 0 37904 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_406
timestamp 1676037725
transform 1 0 38456 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1676037725
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_27
timestamp 1676037725
transform 1 0 3588 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_35
timestamp 1676037725
transform 1 0 4324 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_41
timestamp 1676037725
transform 1 0 4876 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_54
timestamp 1676037725
transform 1 0 6072 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_64
timestamp 1676037725
transform 1 0 6992 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_76
timestamp 1676037725
transform 1 0 8096 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_82
timestamp 1676037725
transform 1 0 8648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_86
timestamp 1676037725
transform 1 0 9016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_96
timestamp 1676037725
transform 1 0 9936 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_106
timestamp 1676037725
transform 1 0 10856 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_123
timestamp 1676037725
transform 1 0 12420 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_132
timestamp 1676037725
transform 1 0 13248 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_140
timestamp 1676037725
transform 1 0 13984 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_148
timestamp 1676037725
transform 1 0 14720 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_158
timestamp 1676037725
transform 1 0 15640 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1676037725
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_179
timestamp 1676037725
transform 1 0 17572 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_186
timestamp 1676037725
transform 1 0 18216 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_198
timestamp 1676037725
transform 1 0 19320 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_206
timestamp 1676037725
transform 1 0 20056 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_214
timestamp 1676037725
transform 1 0 20792 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_218
timestamp 1676037725
transform 1 0 21160 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1676037725
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_232
timestamp 1676037725
transform 1 0 22448 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_238
timestamp 1676037725
transform 1 0 23000 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_246
timestamp 1676037725
transform 1 0 23736 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_259
timestamp 1676037725
transform 1 0 24932 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_267
timestamp 1676037725
transform 1 0 25668 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1676037725
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1676037725
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_286
timestamp 1676037725
transform 1 0 27416 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_304
timestamp 1676037725
transform 1 0 29072 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_324
timestamp 1676037725
transform 1 0 30912 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_337
timestamp 1676037725
transform 1 0 32108 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_343
timestamp 1676037725
transform 1 0 32660 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_361
timestamp 1676037725
transform 1 0 34316 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_374
timestamp 1676037725
transform 1 0 35512 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_386
timestamp 1676037725
transform 1 0 36616 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_55_393
timestamp 1676037725
transform 1 0 37260 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1676037725
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1676037725
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_40
timestamp 1676037725
transform 1 0 4784 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_51
timestamp 1676037725
transform 1 0 5796 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_59
timestamp 1676037725
transform 1 0 6532 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_64
timestamp 1676037725
transform 1 0 6992 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_73
timestamp 1676037725
transform 1 0 7820 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_81
timestamp 1676037725
transform 1 0 8556 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_102
timestamp 1676037725
transform 1 0 10488 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_113
timestamp 1676037725
transform 1 0 11500 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_56_126
timestamp 1676037725
transform 1 0 12696 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_134
timestamp 1676037725
transform 1 0 13432 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1676037725
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_154
timestamp 1676037725
transform 1 0 15272 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_163
timestamp 1676037725
transform 1 0 16100 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_175
timestamp 1676037725
transform 1 0 17204 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_182
timestamp 1676037725
transform 1 0 17848 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_190
timestamp 1676037725
transform 1 0 18584 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_201
timestamp 1676037725
transform 1 0 19596 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_205
timestamp 1676037725
transform 1 0 19964 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_217
timestamp 1676037725
transform 1 0 21068 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_225
timestamp 1676037725
transform 1 0 21804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_230
timestamp 1676037725
transform 1 0 22264 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_243
timestamp 1676037725
transform 1 0 23460 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1676037725
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_266
timestamp 1676037725
transform 1 0 25576 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_270
timestamp 1676037725
transform 1 0 25944 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_287
timestamp 1676037725
transform 1 0 27508 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_304
timestamp 1676037725
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_309
timestamp 1676037725
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_319
timestamp 1676037725
transform 1 0 30452 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_331
timestamp 1676037725
transform 1 0 31556 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_342
timestamp 1676037725
transform 1 0 32568 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_354
timestamp 1676037725
transform 1 0 33672 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_362
timestamp 1676037725
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_365
timestamp 1676037725
transform 1 0 34684 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_373
timestamp 1676037725
transform 1 0 35420 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_384
timestamp 1676037725
transform 1 0 36432 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_405
timestamp 1676037725
transform 1 0 38364 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1676037725
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1676037725
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_39
timestamp 1676037725
transform 1 0 4692 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_45
timestamp 1676037725
transform 1 0 5244 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_53
timestamp 1676037725
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_63
timestamp 1676037725
transform 1 0 6900 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_70
timestamp 1676037725
transform 1 0 7544 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_83
timestamp 1676037725
transform 1 0 8740 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_95
timestamp 1676037725
transform 1 0 9844 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_122
timestamp 1676037725
transform 1 0 12328 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_136
timestamp 1676037725
transform 1 0 13616 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_148
timestamp 1676037725
transform 1 0 14720 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_154
timestamp 1676037725
transform 1 0 15272 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_163
timestamp 1676037725
transform 1 0 16100 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1676037725
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_187
timestamp 1676037725
transform 1 0 18308 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_202
timestamp 1676037725
transform 1 0 19688 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_212
timestamp 1676037725
transform 1 0 20608 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_218
timestamp 1676037725
transform 1 0 21160 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 1676037725
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_231
timestamp 1676037725
transform 1 0 22356 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_241
timestamp 1676037725
transform 1 0 23276 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_254
timestamp 1676037725
transform 1 0 24472 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_267
timestamp 1676037725
transform 1 0 25668 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1676037725
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_281
timestamp 1676037725
transform 1 0 26956 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_285
timestamp 1676037725
transform 1 0 27324 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_295
timestamp 1676037725
transform 1 0 28244 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_306
timestamp 1676037725
transform 1 0 29256 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_319
timestamp 1676037725
transform 1 0 30452 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_334
timestamp 1676037725
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_337
timestamp 1676037725
transform 1 0 32108 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_353
timestamp 1676037725
transform 1 0 33580 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_361
timestamp 1676037725
transform 1 0 34316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_369
timestamp 1676037725
transform 1 0 35052 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_381
timestamp 1676037725
transform 1 0 36156 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_389
timestamp 1676037725
transform 1 0 36892 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_393
timestamp 1676037725
transform 1 0 37260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_404
timestamp 1676037725
transform 1 0 38272 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1676037725
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_45
timestamp 1676037725
transform 1 0 5244 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_55
timestamp 1676037725
transform 1 0 6164 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_63
timestamp 1676037725
transform 1 0 6900 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 1676037725
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_98
timestamp 1676037725
transform 1 0 10120 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_58_111
timestamp 1676037725
transform 1 0 11316 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_120
timestamp 1676037725
transform 1 0 12144 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_132
timestamp 1676037725
transform 1 0 13248 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_153
timestamp 1676037725
transform 1 0 15180 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_157
timestamp 1676037725
transform 1 0 15548 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_169
timestamp 1676037725
transform 1 0 16652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_173
timestamp 1676037725
transform 1 0 17020 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_188
timestamp 1676037725
transform 1 0 18400 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_202
timestamp 1676037725
transform 1 0 19688 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_209
timestamp 1676037725
transform 1 0 20332 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_215
timestamp 1676037725
transform 1 0 20884 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_224
timestamp 1676037725
transform 1 0 21712 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_236
timestamp 1676037725
transform 1 0 22816 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1676037725
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_264
timestamp 1676037725
transform 1 0 25392 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_274
timestamp 1676037725
transform 1 0 26312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_282
timestamp 1676037725
transform 1 0 27048 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_295
timestamp 1676037725
transform 1 0 28244 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_306
timestamp 1676037725
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 1676037725
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_319
timestamp 1676037725
transform 1 0 30452 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_335
timestamp 1676037725
transform 1 0 31924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_347
timestamp 1676037725
transform 1 0 33028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_359
timestamp 1676037725
transform 1 0 34132 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1676037725
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1676037725
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1676037725
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_389
timestamp 1676037725
transform 1 0 36892 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_397
timestamp 1676037725
transform 1 0 37628 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_405
timestamp 1676037725
transform 1 0 38364 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1676037725
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_27
timestamp 1676037725
transform 1 0 3588 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1676037725
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1676037725
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_65
timestamp 1676037725
transform 1 0 7084 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_79
timestamp 1676037725
transform 1 0 8372 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_91
timestamp 1676037725
transform 1 0 9476 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_101
timestamp 1676037725
transform 1 0 10396 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_109
timestamp 1676037725
transform 1 0 11132 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1676037725
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1676037725
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1676037725
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1676037725
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1676037725
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_177
timestamp 1676037725
transform 1 0 17388 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_199
timestamp 1676037725
transform 1 0 19412 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_205
timestamp 1676037725
transform 1 0 19964 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_211
timestamp 1676037725
transform 1 0 20516 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1676037725
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_238
timestamp 1676037725
transform 1 0 23000 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_242
timestamp 1676037725
transform 1 0 23368 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_249
timestamp 1676037725
transform 1 0 24012 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_257
timestamp 1676037725
transform 1 0 24748 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_272
timestamp 1676037725
transform 1 0 26128 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1676037725
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_290
timestamp 1676037725
transform 1 0 27784 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_299
timestamp 1676037725
transform 1 0 28612 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_309
timestamp 1676037725
transform 1 0 29532 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_321
timestamp 1676037725
transform 1 0 30636 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_333
timestamp 1676037725
transform 1 0 31740 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_337
timestamp 1676037725
transform 1 0 32108 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_352
timestamp 1676037725
transform 1 0 33488 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_358
timestamp 1676037725
transform 1 0 34040 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_376
timestamp 1676037725
transform 1 0 35696 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_380
timestamp 1676037725
transform 1 0 36064 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_390
timestamp 1676037725
transform 1 0 36984 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_393
timestamp 1676037725
transform 1 0 37260 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1676037725
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1676037725
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_52
timestamp 1676037725
transform 1 0 5888 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_64
timestamp 1676037725
transform 1 0 6992 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_76
timestamp 1676037725
transform 1 0 8096 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_103
timestamp 1676037725
transform 1 0 10580 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_109
timestamp 1676037725
transform 1 0 11132 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_119
timestamp 1676037725
transform 1 0 12052 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_135
timestamp 1676037725
transform 1 0 13524 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1676037725
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_147
timestamp 1676037725
transform 1 0 14628 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_151
timestamp 1676037725
transform 1 0 14996 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_176
timestamp 1676037725
transform 1 0 17296 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_184
timestamp 1676037725
transform 1 0 18032 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1676037725
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_209
timestamp 1676037725
transform 1 0 20332 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_219
timestamp 1676037725
transform 1 0 21252 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_227
timestamp 1676037725
transform 1 0 21988 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_234
timestamp 1676037725
transform 1 0 22632 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1676037725
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_281
timestamp 1676037725
transform 1 0 26956 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_290
timestamp 1676037725
transform 1 0 27784 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_298
timestamp 1676037725
transform 1 0 28520 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_305
timestamp 1676037725
transform 1 0 29164 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1676037725
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_329
timestamp 1676037725
transform 1 0 31372 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_341
timestamp 1676037725
transform 1 0 32476 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_350
timestamp 1676037725
transform 1 0 33304 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1676037725
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1676037725
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_377
timestamp 1676037725
transform 1 0 35788 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_381
timestamp 1676037725
transform 1 0 36156 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_399
timestamp 1676037725
transform 1 0 37812 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1676037725
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1676037725
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1676037725
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_74
timestamp 1676037725
transform 1 0 7912 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_86
timestamp 1676037725
transform 1 0 9016 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_101
timestamp 1676037725
transform 1 0 10396 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_109
timestamp 1676037725
transform 1 0 11132 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_124
timestamp 1676037725
transform 1 0 12512 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_132
timestamp 1676037725
transform 1 0 13248 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_154
timestamp 1676037725
transform 1 0 15272 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_166
timestamp 1676037725
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_174
timestamp 1676037725
transform 1 0 17112 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_186
timestamp 1676037725
transform 1 0 18216 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_198
timestamp 1676037725
transform 1 0 19320 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_202
timestamp 1676037725
transform 1 0 19688 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_206
timestamp 1676037725
transform 1 0 20056 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_216
timestamp 1676037725
transform 1 0 20976 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_236
timestamp 1676037725
transform 1 0 22816 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_247
timestamp 1676037725
transform 1 0 23828 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_255
timestamp 1676037725
transform 1 0 24564 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_269
timestamp 1676037725
transform 1 0 25852 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_273
timestamp 1676037725
transform 1 0 26220 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 1676037725
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1676037725
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_292
timestamp 1676037725
transform 1 0 27968 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_298
timestamp 1676037725
transform 1 0 28520 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_316
timestamp 1676037725
transform 1 0 30176 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_328
timestamp 1676037725
transform 1 0 31280 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_337
timestamp 1676037725
transform 1 0 32108 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_343
timestamp 1676037725
transform 1 0 32660 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_348
timestamp 1676037725
transform 1 0 33120 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_352
timestamp 1676037725
transform 1 0 33488 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_356
timestamp 1676037725
transform 1 0 33856 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_368
timestamp 1676037725
transform 1 0 34960 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_380
timestamp 1676037725
transform 1 0 36064 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_386
timestamp 1676037725
transform 1 0 36616 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1676037725
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_393
timestamp 1676037725
transform 1 0 37260 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_404
timestamp 1676037725
transform 1 0 38272 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_53
timestamp 1676037725
transform 1 0 5980 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_73
timestamp 1676037725
transform 1 0 7820 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_81
timestamp 1676037725
transform 1 0 8556 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_96
timestamp 1676037725
transform 1 0 9936 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_118
timestamp 1676037725
transform 1 0 11960 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_124
timestamp 1676037725
transform 1 0 12512 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_134
timestamp 1676037725
transform 1 0 13432 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_156
timestamp 1676037725
transform 1 0 15456 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_181
timestamp 1676037725
transform 1 0 17756 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_187
timestamp 1676037725
transform 1 0 18308 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1676037725
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_202
timestamp 1676037725
transform 1 0 19688 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_214
timestamp 1676037725
transform 1 0 20792 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_241
timestamp 1676037725
transform 1 0 23276 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_249
timestamp 1676037725
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_267
timestamp 1676037725
transform 1 0 25668 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_290
timestamp 1676037725
transform 1 0 27784 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_300
timestamp 1676037725
transform 1 0 28704 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_309
timestamp 1676037725
transform 1 0 29532 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_318
timestamp 1676037725
transform 1 0 30360 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_333
timestamp 1676037725
transform 1 0 31740 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_341
timestamp 1676037725
transform 1 0 32476 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_345
timestamp 1676037725
transform 1 0 32844 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_354
timestamp 1676037725
transform 1 0 33672 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_362
timestamp 1676037725
transform 1 0 34408 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_365
timestamp 1676037725
transform 1 0 34684 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_384
timestamp 1676037725
transform 1 0 36432 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1676037725
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1676037725
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_27
timestamp 1676037725
transform 1 0 3588 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_35
timestamp 1676037725
transform 1 0 4324 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1676037725
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_68
timestamp 1676037725
transform 1 0 7360 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_90
timestamp 1676037725
transform 1 0 9384 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_102
timestamp 1676037725
transform 1 0 10488 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1676037725
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_135
timestamp 1676037725
transform 1 0 13524 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_163
timestamp 1676037725
transform 1 0 16100 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_174
timestamp 1676037725
transform 1 0 17112 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_180
timestamp 1676037725
transform 1 0 17664 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_201
timestamp 1676037725
transform 1 0 19596 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_218
timestamp 1676037725
transform 1 0 21160 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_243
timestamp 1676037725
transform 1 0 23460 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_247
timestamp 1676037725
transform 1 0 23828 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_269
timestamp 1676037725
transform 1 0 25852 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1676037725
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_281
timestamp 1676037725
transform 1 0 26956 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_303
timestamp 1676037725
transform 1 0 28980 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_307
timestamp 1676037725
transform 1 0 29348 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_324
timestamp 1676037725
transform 1 0 30912 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1676037725
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_356
timestamp 1676037725
transform 1 0 33856 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_377
timestamp 1676037725
transform 1 0 35788 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_383
timestamp 1676037725
transform 1 0 36340 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1676037725
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_393
timestamp 1676037725
transform 1 0 37260 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1676037725
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_7
timestamp 1676037725
transform 1 0 1748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_20
timestamp 1676037725
transform 1 0 2944 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_54
timestamp 1676037725
transform 1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_57
timestamp 1676037725
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_69
timestamp 1676037725
transform 1 0 7452 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1676037725
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_96
timestamp 1676037725
transform 1 0 9936 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_108
timestamp 1676037725
transform 1 0 11040 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_113
timestamp 1676037725
transform 1 0 11500 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_128
timestamp 1676037725
transform 1 0 12880 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_149
timestamp 1676037725
transform 1 0 14812 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_161
timestamp 1676037725
transform 1 0 15916 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1676037725
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_169
timestamp 1676037725
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_181
timestamp 1676037725
transform 1 0 17756 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1676037725
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1676037725
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_221
timestamp 1676037725
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1676037725
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_239
timestamp 1676037725
transform 1 0 23092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1676037725
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_259
timestamp 1676037725
transform 1 0 24932 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_269
timestamp 1676037725
transform 1 0 25852 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_278
timestamp 1676037725
transform 1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_281
timestamp 1676037725
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_293
timestamp 1676037725
transform 1 0 28060 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_300
timestamp 1676037725
transform 1 0 28704 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1676037725
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1676037725
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_333
timestamp 1676037725
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1676037725
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_343
timestamp 1676037725
transform 1 0 32660 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_351
timestamp 1676037725
transform 1 0 33396 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_358
timestamp 1676037725
transform 1 0 34040 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1676037725
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_377
timestamp 1676037725
transform 1 0 35788 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_383
timestamp 1676037725
transform 1 0 36340 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_390
timestamp 1676037725
transform 1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_393
timestamp 1676037725
transform 1 0 37260 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1676037725
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0828_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28336 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1676037725
transform 1 0 27508 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0830_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20424 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1676037725
transform 1 0 18676 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1676037725
transform 1 0 14996 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1676037725
transform 1 0 16008 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1676037725
transform 1 0 14628 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1676037725
transform 1 0 15180 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1676037725
transform 1 0 15272 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0838_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27968 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_8  _0839_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21344 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_8  _0840_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8096 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__clkinv_4  _0841_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _0842_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0843_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8280 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_4  _0844_
timestamp 1676037725
transform 1 0 5336 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_4  _0845_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12420 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_8  _0846_
timestamp 1676037725
transform 1 0 12144 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1676037725
transform 1 0 8372 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0848_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27324 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0849_
timestamp 1676037725
transform 1 0 21068 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0850_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18216 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0851_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23276 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0852_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19780 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0853_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0855_
timestamp 1676037725
transform 1 0 23644 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0856_
timestamp 1676037725
transform 1 0 26864 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _0857_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_4  _0858_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24748 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _0859_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26220 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0860_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0861_
timestamp 1676037725
transform 1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _0862_
timestamp 1676037725
transform 1 0 28612 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_4  _0863_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_8  _0864_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24748 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_4  _0865_
timestamp 1676037725
transform 1 0 24932 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0866_
timestamp 1676037725
transform 1 0 20056 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _0867_
timestamp 1676037725
transform 1 0 21988 0 -1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__or3b_4  _0868_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0869_
timestamp 1676037725
transform 1 0 23184 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0870_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24840 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0871_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25852 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0872_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20056 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _0873_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0874_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25576 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand4b_4  _0875_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17664 0 -1 34816
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_2  _0876_
timestamp 1676037725
transform 1 0 19412 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _0877_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0878_
timestamp 1676037725
transform 1 0 27048 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_4  _0879_
timestamp 1676037725
transform 1 0 17940 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_2  _0880_
timestamp 1676037725
transform 1 0 25484 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0881_
timestamp 1676037725
transform 1 0 24104 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _0882_
timestamp 1676037725
transform 1 0 22080 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0883_
timestamp 1676037725
transform 1 0 20332 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0884_
timestamp 1676037725
transform 1 0 21988 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0885_
timestamp 1676037725
transform 1 0 21252 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _0886_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21896 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0887_
timestamp 1676037725
transform 1 0 22632 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1676037725
transform 1 0 15824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0889_
timestamp 1676037725
transform 1 0 24288 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0890_
timestamp 1676037725
transform 1 0 26680 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0891_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24932 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0892_
timestamp 1676037725
transform 1 0 29348 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1676037725
transform 1 0 36708 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0894_
timestamp 1676037725
transform 1 0 23092 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0895_
timestamp 1676037725
transform 1 0 17848 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0896_
timestamp 1676037725
transform 1 0 25760 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_4  _0897_
timestamp 1676037725
transform 1 0 17204 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _0898_
timestamp 1676037725
transform 1 0 18860 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0899_
timestamp 1676037725
transform 1 0 22724 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _0900_
timestamp 1676037725
transform 1 0 20792 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0901_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0902_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0903_
timestamp 1676037725
transform 1 0 11868 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0904_
timestamp 1676037725
transform 1 0 20240 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_4  _0905_
timestamp 1676037725
transform 1 0 24564 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _0906_
timestamp 1676037725
transform 1 0 20608 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _0907_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25944 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _0908_
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _0909_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21160 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_4  _0910_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_2  _0911_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22540 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0912_
timestamp 1676037725
transform 1 0 19320 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _0913_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20148 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0914_
timestamp 1676037725
transform 1 0 19964 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0915_
timestamp 1676037725
transform 1 0 19412 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_4  _0916_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16928 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__or4_4  _0917_
timestamp 1676037725
transform 1 0 24840 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1676037725
transform 1 0 21252 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0919_
timestamp 1676037725
transform 1 0 21988 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _0920_
timestamp 1676037725
transform 1 0 16928 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0921_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0922_
timestamp 1676037725
transform 1 0 23828 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _0923_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23552 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1676037725
transform 1 0 27692 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0925_
timestamp 1676037725
transform 1 0 18032 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _0926_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20700 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0927_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25760 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_4  _0928_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16560 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__o22ai_1  _0929_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18860 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0930_
timestamp 1676037725
transform 1 0 22632 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _0931_
timestamp 1676037725
transform 1 0 27140 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _0932_
timestamp 1676037725
transform 1 0 26680 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _0933_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19964 0 -1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__a32o_1  _0934_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19596 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_2  _0935_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nand4b_4  _0936_
timestamp 1676037725
transform 1 0 16836 0 -1 25024
box -38 -48 1786 592
use sky130_fd_sc_hd__o31a_1  _0937_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _0938_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14904 0 1 26112
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_4  _0939_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27600 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_8  _0940_
timestamp 1676037725
transform 1 0 18216 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__and4_1  _0941_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16560 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_4  _0942_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16744 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__or2_1  _0943_
timestamp 1676037725
transform 1 0 33764 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0944_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_8  _0945_
timestamp 1676037725
transform 1 0 30268 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_8  _0946_
timestamp 1676037725
transform 1 0 33488 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__a221oi_4  _0947_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34960 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _0948_
timestamp 1676037725
transform 1 0 27784 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_8  _0949_
timestamp 1676037725
transform 1 0 22448 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_4  _0950_
timestamp 1676037725
transform 1 0 21620 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_4  _0951_
timestamp 1676037725
transform 1 0 23000 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _0952_
timestamp 1676037725
transform 1 0 24564 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _0953_
timestamp 1676037725
transform 1 0 22448 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_4  _0954_
timestamp 1676037725
transform 1 0 23644 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0955_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23368 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0956_
timestamp 1676037725
transform 1 0 22540 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _0957_
timestamp 1676037725
transform 1 0 25668 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _0958_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28428 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _0959_
timestamp 1676037725
transform 1 0 24288 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0960_
timestamp 1676037725
transform 1 0 18676 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0961_
timestamp 1676037725
transform 1 0 34868 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0962_
timestamp 1676037725
transform 1 0 34776 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _0963_
timestamp 1676037725
transform 1 0 35052 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _0964_
timestamp 1676037725
transform 1 0 27876 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _0965_
timestamp 1676037725
transform 1 0 27600 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _0966_
timestamp 1676037725
transform 1 0 24748 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _0967_
timestamp 1676037725
transform 1 0 20424 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0968_
timestamp 1676037725
transform 1 0 20608 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0969_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21160 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0970_
timestamp 1676037725
transform 1 0 19688 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0971_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20056 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _0972_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20148 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _0973_
timestamp 1676037725
transform 1 0 20976 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_4  _0974_
timestamp 1676037725
transform 1 0 21988 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0975_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0976_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17756 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _0977_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18768 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _0978_
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_1  _0979_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18492 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _0980_
timestamp 1676037725
transform 1 0 17572 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _0981_
timestamp 1676037725
transform 1 0 17388 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0982_
timestamp 1676037725
transform 1 0 17480 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0983_
timestamp 1676037725
transform 1 0 17388 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1676037725
transform 1 0 17112 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0985_
timestamp 1676037725
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0986_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17296 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_2  _0987_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17204 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _0988_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22080 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1676037725
transform 1 0 15640 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _0990_
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1676037725
transform 1 0 16100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0992_
timestamp 1676037725
transform 1 0 15364 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0993_
timestamp 1676037725
transform 1 0 15088 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0994_
timestamp 1676037725
transform 1 0 16836 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0995_
timestamp 1676037725
transform 1 0 14444 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_4  _0996_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13892 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__or2_1  _0997_
timestamp 1676037725
transform 1 0 33028 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0998_
timestamp 1676037725
transform 1 0 31832 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _0999_
timestamp 1676037725
transform 1 0 32292 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_1  _1000_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28336 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1001_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28244 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _1002_
timestamp 1676037725
transform 1 0 27692 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1003_
timestamp 1676037725
transform 1 0 23092 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1004_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22448 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1005_
timestamp 1676037725
transform 1 0 21712 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1006_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21528 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1007_
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1008_
timestamp 1676037725
transform 1 0 20700 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1009_
timestamp 1676037725
transform 1 0 16192 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1676037725
transform 1 0 17480 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1011_
timestamp 1676037725
transform 1 0 20700 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1012_
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1013_
timestamp 1676037725
transform 1 0 20148 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1014_
timestamp 1676037725
transform 1 0 21988 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1015_
timestamp 1676037725
transform 1 0 33580 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1016_
timestamp 1676037725
transform 1 0 34868 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _1017_
timestamp 1676037725
transform 1 0 35328 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_1  _1018_
timestamp 1676037725
transform 1 0 28152 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1019_
timestamp 1676037725
transform 1 0 27140 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _1020_
timestamp 1676037725
transform 1 0 26680 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1021_
timestamp 1676037725
transform 1 0 21436 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1022_
timestamp 1676037725
transform 1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1023_
timestamp 1676037725
transform 1 0 21528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1024_
timestamp 1676037725
transform 1 0 20884 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1025_
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1026_
timestamp 1676037725
transform 1 0 20976 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1027_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20884 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _1028_
timestamp 1676037725
transform 1 0 20700 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1676037725
transform 1 0 19504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1030_
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _1031_
timestamp 1676037725
transform 1 0 20148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_1  _1032_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1033_
timestamp 1676037725
transform 1 0 24472 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1034_
timestamp 1676037725
transform 1 0 25852 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1035_
timestamp 1676037725
transform 1 0 25760 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1036_
timestamp 1676037725
transform 1 0 25024 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1037_
timestamp 1676037725
transform 1 0 27968 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1038_
timestamp 1676037725
transform 1 0 25852 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _1039_
timestamp 1676037725
transform 1 0 25300 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1040_
timestamp 1676037725
transform 1 0 20792 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1041_
timestamp 1676037725
transform 1 0 19596 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1042_
timestamp 1676037725
transform 1 0 19596 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1043_
timestamp 1676037725
transform 1 0 18952 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1044_
timestamp 1676037725
transform 1 0 18584 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1045_
timestamp 1676037725
transform 1 0 19320 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1046_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1047_
timestamp 1676037725
transform 1 0 19412 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1048_
timestamp 1676037725
transform 1 0 18492 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1049_
timestamp 1676037725
transform 1 0 16468 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1050_
timestamp 1676037725
transform 1 0 29256 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1051_
timestamp 1676037725
transform 1 0 30452 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _1052_
timestamp 1676037725
transform 1 0 29716 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1053_
timestamp 1676037725
transform 1 0 27508 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1054_
timestamp 1676037725
transform 1 0 28060 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1055_
timestamp 1676037725
transform 1 0 27600 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1056_
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1057_
timestamp 1676037725
transform 1 0 17940 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1058_
timestamp 1676037725
transform 1 0 17112 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1059_
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1060_
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1061_
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1062_
timestamp 1676037725
transform 1 0 17204 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1063_
timestamp 1676037725
transform 1 0 14996 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_4  _1064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20976 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__and3_1  _1065_
timestamp 1676037725
transform 1 0 25944 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1066_
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1067_
timestamp 1676037725
transform 1 0 26220 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1068_
timestamp 1676037725
transform 1 0 24748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1069_
timestamp 1676037725
transform 1 0 25300 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1070_
timestamp 1676037725
transform 1 0 25944 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1071_
timestamp 1676037725
transform 1 0 25852 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1072_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _1073_
timestamp 1676037725
transform 1 0 15640 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17664 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _1075_
timestamp 1676037725
transform 1 0 15732 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_2  _1076_
timestamp 1676037725
transform 1 0 14904 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _1077_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _1078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__and2b_1  _1079_
timestamp 1676037725
transform 1 0 13248 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1080_
timestamp 1676037725
transform 1 0 15088 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1081_
timestamp 1676037725
transform 1 0 14352 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1082_
timestamp 1676037725
transform 1 0 15640 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1083_
timestamp 1676037725
transform 1 0 16560 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1084_
timestamp 1676037725
transform 1 0 16836 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1085_
timestamp 1676037725
transform 1 0 16836 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1086_
timestamp 1676037725
transform 1 0 22540 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1087_
timestamp 1676037725
transform 1 0 18308 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1088_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22448 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1089_
timestamp 1676037725
transform 1 0 15272 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1090_
timestamp 1676037725
transform 1 0 14260 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1091_
timestamp 1676037725
transform 1 0 13156 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1092_
timestamp 1676037725
transform 1 0 13340 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_4  _1093_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_2  _1094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16100 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_2  _1095_
timestamp 1676037725
transform 1 0 15456 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _1096_
timestamp 1676037725
transform 1 0 15456 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_2  _1097_
timestamp 1676037725
transform 1 0 18308 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1098_
timestamp 1676037725
transform 1 0 18124 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1099_
timestamp 1676037725
transform 1 0 17020 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1100_
timestamp 1676037725
transform 1 0 18216 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _1101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_4  _1102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17940 0 -1 6528
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _1103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 2062 592
use sky130_fd_sc_hd__o211ai_4  _1104_
timestamp 1676037725
transform 1 0 17940 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_2  _1105_
timestamp 1676037725
transform 1 0 15272 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_4  _1106_
timestamp 1676037725
transform 1 0 17020 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _1107_
timestamp 1676037725
transform 1 0 21528 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1108_
timestamp 1676037725
transform 1 0 19964 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__o21bai_4  _1109_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__o211ai_4  _1110_
timestamp 1676037725
transform 1 0 13800 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__or2_1  _1111_
timestamp 1676037725
transform 1 0 28336 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1112_
timestamp 1676037725
transform 1 0 29164 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _1113_
timestamp 1676037725
transform 1 0 29716 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _1114_
timestamp 1676037725
transform 1 0 28980 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1115_
timestamp 1676037725
transform 1 0 28244 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _1116_
timestamp 1676037725
transform 1 0 27692 0 1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_2  _1117_
timestamp 1676037725
transform 1 0 21252 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1118_
timestamp 1676037725
transform 1 0 19780 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1119_
timestamp 1676037725
transform 1 0 19504 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1120_
timestamp 1676037725
transform 1 0 19228 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1121_
timestamp 1676037725
transform 1 0 18952 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1122_
timestamp 1676037725
transform 1 0 12512 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1123_
timestamp 1676037725
transform 1 0 14996 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _1124_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13156 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1125_
timestamp 1676037725
transform 1 0 13156 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1126_
timestamp 1676037725
transform 1 0 12604 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1127_
timestamp 1676037725
transform 1 0 11776 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1128_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12696 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1129_
timestamp 1676037725
transform 1 0 11684 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _1130_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1131_
timestamp 1676037725
transform 1 0 14996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1132_
timestamp 1676037725
transform 1 0 16192 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1133_
timestamp 1676037725
transform 1 0 16928 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1134_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14168 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1135_
timestamp 1676037725
transform 1 0 14720 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1136_
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1137_
timestamp 1676037725
transform 1 0 12328 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1138_
timestamp 1676037725
transform 1 0 12144 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1139_
timestamp 1676037725
transform 1 0 11776 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1140_
timestamp 1676037725
transform 1 0 10672 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1141_
timestamp 1676037725
transform 1 0 11224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1142_
timestamp 1676037725
transform 1 0 10488 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1143_
timestamp 1676037725
transform 1 0 14260 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1144_
timestamp 1676037725
transform 1 0 12144 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1145_
timestamp 1676037725
transform 1 0 10948 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _1146_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _1147_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1148_
timestamp 1676037725
transform 1 0 10396 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1149_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1150_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13156 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1151_
timestamp 1676037725
transform 1 0 29716 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1152_
timestamp 1676037725
transform 1 0 25852 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1153_
timestamp 1676037725
transform 1 0 28520 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _1154_
timestamp 1676037725
transform 1 0 25852 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _1155_
timestamp 1676037725
transform 1 0 27784 0 -1 32640
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_2  _1156_
timestamp 1676037725
transform 1 0 29716 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_8  _1157_
timestamp 1676037725
transform 1 0 27140 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__o31ai_4  _1158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30268 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_8  _1159_
timestamp 1676037725
transform 1 0 28980 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__a22o_1  _1160_
timestamp 1676037725
transform 1 0 30820 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1161_
timestamp 1676037725
transform 1 0 30544 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1162_
timestamp 1676037725
transform 1 0 25944 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1163_
timestamp 1676037725
transform 1 0 27140 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1164_
timestamp 1676037725
transform 1 0 22724 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1165_
timestamp 1676037725
transform 1 0 24564 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1166_
timestamp 1676037725
transform 1 0 25760 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1167_
timestamp 1676037725
transform 1 0 26220 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1168_
timestamp 1676037725
transform 1 0 27324 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1169_
timestamp 1676037725
transform 1 0 29164 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28152 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_8  _1172_
timestamp 1676037725
transform 1 0 26036 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__or4_2  _1173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29348 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1174_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31832 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1175_
timestamp 1676037725
transform 1 0 32936 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1176_
timestamp 1676037725
transform 1 0 33856 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1177_
timestamp 1676037725
transform 1 0 33488 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _1178_
timestamp 1676037725
transform 1 0 28612 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1179_
timestamp 1676037725
transform 1 0 31832 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_4  _1180_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32384 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__or3b_2  _1181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33120 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1182_
timestamp 1676037725
transform 1 0 33028 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _1183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30636 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__a221o_1  _1184_
timestamp 1676037725
transform 1 0 32752 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1185_
timestamp 1676037725
transform 1 0 32844 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1186_
timestamp 1676037725
transform 1 0 33304 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1187_
timestamp 1676037725
transform 1 0 33488 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1188_
timestamp 1676037725
transform 1 0 32476 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1189_
timestamp 1676037725
transform 1 0 32568 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1190_
timestamp 1676037725
transform 1 0 33580 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1191_
timestamp 1676037725
transform 1 0 32936 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1192_
timestamp 1676037725
transform 1 0 32568 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1193_
timestamp 1676037725
transform 1 0 32660 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1194_
timestamp 1676037725
transform 1 0 33120 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1195_
timestamp 1676037725
transform 1 0 33672 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1196_
timestamp 1676037725
transform 1 0 32936 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1197_
timestamp 1676037725
transform 1 0 34316 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1198_
timestamp 1676037725
transform 1 0 33488 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1199_
timestamp 1676037725
transform 1 0 33764 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1200_
timestamp 1676037725
transform 1 0 32292 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _1201_
timestamp 1676037725
transform 1 0 32384 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1202_
timestamp 1676037725
transform 1 0 33948 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1203_
timestamp 1676037725
transform 1 0 32936 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1204_
timestamp 1676037725
transform 1 0 32936 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1205_
timestamp 1676037725
transform 1 0 30360 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1206_
timestamp 1676037725
transform 1 0 28612 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1207_
timestamp 1676037725
transform 1 0 30820 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1208_
timestamp 1676037725
transform 1 0 31280 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1209_
timestamp 1676037725
transform 1 0 32568 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1210_
timestamp 1676037725
transform 1 0 30084 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1211_
timestamp 1676037725
transform 1 0 31096 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1212_
timestamp 1676037725
transform 1 0 32292 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1213_
timestamp 1676037725
transform 1 0 32384 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1214_
timestamp 1676037725
transform 1 0 33120 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1215_
timestamp 1676037725
transform 1 0 29808 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1216_
timestamp 1676037725
transform 1 0 30728 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1217_
timestamp 1676037725
transform 1 0 32108 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1218_
timestamp 1676037725
transform 1 0 29716 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1219_
timestamp 1676037725
transform 1 0 30636 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1220_
timestamp 1676037725
transform 1 0 32292 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1221_
timestamp 1676037725
transform 1 0 32016 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1222_
timestamp 1676037725
transform 1 0 32752 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1223_
timestamp 1676037725
transform 1 0 30176 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1224_
timestamp 1676037725
transform 1 0 31004 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1225_
timestamp 1676037725
transform 1 0 32844 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1226_
timestamp 1676037725
transform 1 0 30820 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1227_
timestamp 1676037725
transform 1 0 31188 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1228_
timestamp 1676037725
transform 1 0 32844 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1229_
timestamp 1676037725
transform 1 0 32752 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1230_
timestamp 1676037725
transform 1 0 33580 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1231_
timestamp 1676037725
transform 1 0 29716 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1232_
timestamp 1676037725
transform 1 0 31740 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1233_
timestamp 1676037725
transform 1 0 32568 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1234_
timestamp 1676037725
transform 1 0 33212 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1235_
timestamp 1676037725
transform 1 0 33580 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1236_
timestamp 1676037725
transform 1 0 29716 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1237_
timestamp 1676037725
transform 1 0 30636 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1238_
timestamp 1676037725
transform 1 0 31096 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1239_
timestamp 1676037725
transform 1 0 20332 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1240_
timestamp 1676037725
transform 1 0 21160 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1241_
timestamp 1676037725
transform 1 0 18032 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1242_
timestamp 1676037725
transform 1 0 9568 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1243_
timestamp 1676037725
transform 1 0 5336 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1244_
timestamp 1676037725
transform 1 0 6716 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1245_
timestamp 1676037725
transform 1 0 11224 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1246_
timestamp 1676037725
transform 1 0 9936 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _1247_
timestamp 1676037725
transform 1 0 7268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1248_
timestamp 1676037725
transform 1 0 5336 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1249_
timestamp 1676037725
transform 1 0 5152 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1250_
timestamp 1676037725
transform 1 0 5152 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1251_
timestamp 1676037725
transform 1 0 4416 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1252_
timestamp 1676037725
transform 1 0 4324 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and2_4  _1253_
timestamp 1676037725
transform 1 0 4784 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1254_
timestamp 1676037725
transform 1 0 5244 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1255_
timestamp 1676037725
transform 1 0 7360 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_8  _1256_
timestamp 1676037725
transform 1 0 7176 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_4  _1257_
timestamp 1676037725
transform 1 0 8096 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1258_
timestamp 1676037725
transform 1 0 9108 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1259_
timestamp 1676037725
transform 1 0 6532 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_2  _1260_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6348 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1261_
timestamp 1676037725
transform 1 0 12788 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16100 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1263_
timestamp 1676037725
transform 1 0 25392 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1264_
timestamp 1676037725
transform 1 0 15088 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o31ai_1  _1265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14720 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1266_
timestamp 1676037725
transform 1 0 15824 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1267_
timestamp 1676037725
transform 1 0 5336 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _1268_
timestamp 1676037725
transform 1 0 9752 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1269_
timestamp 1676037725
transform 1 0 5704 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1270_
timestamp 1676037725
transform 1 0 9568 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1271_
timestamp 1676037725
transform 1 0 12420 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1272_
timestamp 1676037725
transform 1 0 13248 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1273_
timestamp 1676037725
transform 1 0 15640 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1274_
timestamp 1676037725
transform 1 0 6716 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1275_
timestamp 1676037725
transform 1 0 10948 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1276_
timestamp 1676037725
transform 1 0 6072 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1277_
timestamp 1676037725
transform 1 0 9108 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1278_
timestamp 1676037725
transform 1 0 6808 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _1279_
timestamp 1676037725
transform 1 0 10856 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1280_
timestamp 1676037725
transform 1 0 10856 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1281_
timestamp 1676037725
transform 1 0 18216 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1282_
timestamp 1676037725
transform 1 0 21252 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1283_
timestamp 1676037725
transform 1 0 23644 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1284_
timestamp 1676037725
transform 1 0 16376 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1285_
timestamp 1676037725
transform 1 0 18492 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1286_
timestamp 1676037725
transform 1 0 17572 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1287_
timestamp 1676037725
transform 1 0 17388 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1288_
timestamp 1676037725
transform 1 0 12788 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1289_
timestamp 1676037725
transform 1 0 20332 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1290_
timestamp 1676037725
transform 1 0 16836 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1291_
timestamp 1676037725
transform 1 0 11684 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1292_
timestamp 1676037725
transform 1 0 15548 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1293_
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1294_
timestamp 1676037725
transform 1 0 8832 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1295_
timestamp 1676037725
transform 1 0 12696 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1296_
timestamp 1676037725
transform 1 0 9936 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1297_
timestamp 1676037725
transform 1 0 13156 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1298_
timestamp 1676037725
transform 1 0 18216 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1299_
timestamp 1676037725
transform 1 0 5060 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1300_
timestamp 1676037725
transform 1 0 4508 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1301_
timestamp 1676037725
transform 1 0 8188 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1302_
timestamp 1676037725
transform 1 0 10120 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1303_
timestamp 1676037725
transform 1 0 12696 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1304_
timestamp 1676037725
transform 1 0 14260 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1305_
timestamp 1676037725
transform 1 0 9108 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _1306_
timestamp 1676037725
transform 1 0 9936 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1307_
timestamp 1676037725
transform 1 0 12052 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1308_
timestamp 1676037725
transform 1 0 11776 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1309_
timestamp 1676037725
transform 1 0 11500 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1310_
timestamp 1676037725
transform 1 0 10120 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _1311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17020 0 1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__xnor2_2  _1312_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18032 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _1313_
timestamp 1676037725
transform 1 0 21252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1314_
timestamp 1676037725
transform 1 0 10028 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1315_
timestamp 1676037725
transform 1 0 19412 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _1316_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15088 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1317_
timestamp 1676037725
transform 1 0 12052 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _1318_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13064 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1319_
timestamp 1676037725
transform 1 0 8188 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1320_
timestamp 1676037725
transform 1 0 12512 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1321_
timestamp 1676037725
transform 1 0 7912 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1322_
timestamp 1676037725
transform 1 0 3956 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1323_
timestamp 1676037725
transform 1 0 6532 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1324_
timestamp 1676037725
transform 1 0 7728 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1325_
timestamp 1676037725
transform 1 0 7176 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1326_
timestamp 1676037725
transform 1 0 6624 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1327_
timestamp 1676037725
transform 1 0 6532 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1328_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11408 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _1329_
timestamp 1676037725
transform 1 0 11408 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1330_
timestamp 1676037725
transform 1 0 9200 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _1331_
timestamp 1676037725
transform 1 0 9108 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1332_
timestamp 1676037725
transform 1 0 9660 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _1333_
timestamp 1676037725
transform 1 0 11776 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1334_
timestamp 1676037725
transform 1 0 24932 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1335_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24472 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_2  _1336_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24656 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _1337_
timestamp 1676037725
transform 1 0 19044 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1338_
timestamp 1676037725
transform 1 0 14260 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1339_
timestamp 1676037725
transform 1 0 16836 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1340_
timestamp 1676037725
transform 1 0 14628 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1341_
timestamp 1676037725
transform 1 0 15640 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1342_
timestamp 1676037725
transform 1 0 11868 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1343_
timestamp 1676037725
transform 1 0 13340 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _1344_
timestamp 1676037725
transform 1 0 10672 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1345_
timestamp 1676037725
transform 1 0 16744 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1346_
timestamp 1676037725
transform 1 0 13524 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1347_
timestamp 1676037725
transform 1 0 14168 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1348_
timestamp 1676037725
transform 1 0 13984 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1349_
timestamp 1676037725
transform 1 0 15272 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1350_
timestamp 1676037725
transform 1 0 20332 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1351_
timestamp 1676037725
transform 1 0 19412 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1352_
timestamp 1676037725
transform 1 0 13800 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1353_
timestamp 1676037725
transform 1 0 15364 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1354_
timestamp 1676037725
transform 1 0 22080 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1355_
timestamp 1676037725
transform 1 0 20976 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_4  _1356_
timestamp 1676037725
transform 1 0 22908 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1357_
timestamp 1676037725
transform 1 0 17756 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1358_
timestamp 1676037725
transform 1 0 17296 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1359_
timestamp 1676037725
transform 1 0 12052 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1360_
timestamp 1676037725
transform 1 0 17296 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1361_
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_2  _1362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22724 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1363_
timestamp 1676037725
transform 1 0 23276 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1364_
timestamp 1676037725
transform 1 0 17940 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1365_
timestamp 1676037725
transform 1 0 19412 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1366_
timestamp 1676037725
transform 1 0 18216 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1367_
timestamp 1676037725
transform 1 0 19412 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_4  _1368_
timestamp 1676037725
transform 1 0 29808 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_4  _1369_
timestamp 1676037725
transform 1 0 29900 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_4  _1370_
timestamp 1676037725
transform 1 0 27600 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__o21ai_4  _1371_
timestamp 1676037725
transform 1 0 27876 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_1  _1372_
timestamp 1676037725
transform 1 0 28060 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1373_
timestamp 1676037725
transform 1 0 28888 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1374_
timestamp 1676037725
transform 1 0 22172 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _1375_
timestamp 1676037725
transform 1 0 28336 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _1376_
timestamp 1676037725
transform 1 0 25392 0 -1 30464
box -38 -48 1326 592
use sky130_fd_sc_hd__or3_4  _1377_
timestamp 1676037725
transform 1 0 29900 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_4  _1378_
timestamp 1676037725
transform 1 0 22724 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__a22o_1  _1379_
timestamp 1676037725
transform 1 0 32292 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_4  _1380_
timestamp 1676037725
transform 1 0 30820 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__or4_4  _1381_
timestamp 1676037725
transform 1 0 31280 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _1382_
timestamp 1676037725
transform 1 0 30452 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1383_
timestamp 1676037725
transform 1 0 30820 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1384_
timestamp 1676037725
transform 1 0 35052 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1385_
timestamp 1676037725
transform 1 0 29808 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1386_
timestamp 1676037725
transform 1 0 35512 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1387_
timestamp 1676037725
transform 1 0 35052 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1388_
timestamp 1676037725
transform 1 0 34868 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1389_
timestamp 1676037725
transform 1 0 36156 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1390_
timestamp 1676037725
transform 1 0 35052 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1391_
timestamp 1676037725
transform 1 0 35788 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1392_
timestamp 1676037725
transform 1 0 35512 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1393_
timestamp 1676037725
transform 1 0 34868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1394_
timestamp 1676037725
transform 1 0 32752 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1395_
timestamp 1676037725
transform 1 0 35328 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1396_
timestamp 1676037725
transform 1 0 34960 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1397_
timestamp 1676037725
transform 1 0 35144 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1398_
timestamp 1676037725
transform 1 0 36064 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1399_
timestamp 1676037725
transform 1 0 34776 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1400_
timestamp 1676037725
transform 1 0 34960 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1401_
timestamp 1676037725
transform 1 0 35880 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1402_
timestamp 1676037725
transform 1 0 31832 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1403_
timestamp 1676037725
transform 1 0 30636 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1404_
timestamp 1676037725
transform 1 0 32384 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1405_
timestamp 1676037725
transform 1 0 30820 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _1406_
timestamp 1676037725
transform 1 0 29716 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1407_
timestamp 1676037725
transform 1 0 31924 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1408_
timestamp 1676037725
transform 1 0 32936 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1409_
timestamp 1676037725
transform 1 0 35144 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1410_
timestamp 1676037725
transform 1 0 35236 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1411_
timestamp 1676037725
transform 1 0 36156 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1412_
timestamp 1676037725
transform 1 0 35236 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1413_
timestamp 1676037725
transform 1 0 35696 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1414_
timestamp 1676037725
transform 1 0 35052 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1415_
timestamp 1676037725
transform 1 0 35788 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1416_
timestamp 1676037725
transform 1 0 34500 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1417_
timestamp 1676037725
transform 1 0 35236 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1418_
timestamp 1676037725
transform 1 0 34868 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1419_
timestamp 1676037725
transform 1 0 35696 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1420_
timestamp 1676037725
transform 1 0 34408 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1421_
timestamp 1676037725
transform 1 0 35420 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1422_
timestamp 1676037725
transform 1 0 31924 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1423_
timestamp 1676037725
transform 1 0 32844 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _1424_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26036 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_4  _1425_
timestamp 1676037725
transform 1 0 25944 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__a22o_1  _1426_
timestamp 1676037725
transform 1 0 27140 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1427_
timestamp 1676037725
transform 1 0 26496 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1428_
timestamp 1676037725
transform 1 0 26956 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _1429_
timestamp 1676037725
transform 1 0 27140 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1430_
timestamp 1676037725
transform 1 0 27140 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1431_
timestamp 1676037725
transform 1 0 28704 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _1432_
timestamp 1676037725
transform 1 0 28520 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1433_
timestamp 1676037725
transform 1 0 28152 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1434_
timestamp 1676037725
transform 1 0 29348 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1435_
timestamp 1676037725
transform 1 0 29716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _1436_
timestamp 1676037725
transform 1 0 28888 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1437_
timestamp 1676037725
transform 1 0 26036 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1438_
timestamp 1676037725
transform 1 0 27048 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_4  _1439_
timestamp 1676037725
transform 1 0 27968 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__o21a_1  _1440_
timestamp 1676037725
transform 1 0 27140 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1441_
timestamp 1676037725
transform 1 0 27232 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1442_
timestamp 1676037725
transform 1 0 28980 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_2  _1443_
timestamp 1676037725
transform 1 0 28152 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _1444_
timestamp 1676037725
transform 1 0 28704 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1445_
timestamp 1676037725
transform 1 0 29716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1446_
timestamp 1676037725
transform 1 0 29256 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1447_
timestamp 1676037725
transform 1 0 28336 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1448_
timestamp 1676037725
transform 1 0 29716 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1449_
timestamp 1676037725
transform 1 0 26036 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1450_
timestamp 1676037725
transform 1 0 29808 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1451_
timestamp 1676037725
transform 1 0 29716 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1452_
timestamp 1676037725
transform 1 0 26772 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1453_
timestamp 1676037725
transform 1 0 27784 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _1454_
timestamp 1676037725
transform 1 0 26956 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_4  _1455_
timestamp 1676037725
transform 1 0 17940 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_4  _1456_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22540 0 -1 22848
box -38 -48 1326 592
use sky130_fd_sc_hd__and3_4  _1457_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29348 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1458_
timestamp 1676037725
transform 1 0 24748 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1459_
timestamp 1676037725
transform 1 0 25024 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1460_
timestamp 1676037725
transform 1 0 22724 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _1461_
timestamp 1676037725
transform 1 0 22356 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1462_
timestamp 1676037725
transform 1 0 23092 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1463_
timestamp 1676037725
transform 1 0 24748 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1464_
timestamp 1676037725
transform 1 0 24012 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1465_
timestamp 1676037725
transform 1 0 25392 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1466_
timestamp 1676037725
transform 1 0 25392 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1467_
timestamp 1676037725
transform 1 0 29900 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1468_
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1469_
timestamp 1676037725
transform 1 0 24840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1470_
timestamp 1676037725
transform 1 0 23552 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1471_
timestamp 1676037725
transform 1 0 22724 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_2  _1472_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23276 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1473_
timestamp 1676037725
transform 1 0 25852 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1474_
timestamp 1676037725
transform 1 0 23736 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1475_
timestamp 1676037725
transform 1 0 28612 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1476_
timestamp 1676037725
transform 1 0 29716 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_4  _1477_
timestamp 1676037725
transform 1 0 30544 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _1478_
timestamp 1676037725
transform 1 0 32568 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1479_
timestamp 1676037725
transform 1 0 30820 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1480_
timestamp 1676037725
transform 1 0 32476 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1481_
timestamp 1676037725
transform 1 0 22540 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1482_
timestamp 1676037725
transform 1 0 23368 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1483_
timestamp 1676037725
transform 1 0 23460 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1484_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1485_
timestamp 1676037725
transform 1 0 24380 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _1486_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30544 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1487_
timestamp 1676037725
transform 1 0 33580 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1488_
timestamp 1676037725
transform 1 0 23644 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1489_
timestamp 1676037725
transform 1 0 23000 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1490_
timestamp 1676037725
transform 1 0 22908 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1491_
timestamp 1676037725
transform 1 0 24288 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _1492_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _1493_
timestamp 1676037725
transform 1 0 32936 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1494_
timestamp 1676037725
transform 1 0 23644 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1495_
timestamp 1676037725
transform 1 0 23828 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1496_
timestamp 1676037725
transform 1 0 24748 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1497_
timestamp 1676037725
transform 1 0 24840 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_4  _1498_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _1499_
timestamp 1676037725
transform 1 0 27140 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1500_
timestamp 1676037725
transform 1 0 30268 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1501_
timestamp 1676037725
transform 1 0 24932 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1502_
timestamp 1676037725
transform 1 0 28060 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1503_
timestamp 1676037725
transform 1 0 23276 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1504_
timestamp 1676037725
transform 1 0 35052 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1505_
timestamp 1676037725
transform 1 0 31096 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1506_
timestamp 1676037725
transform 1 0 34960 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1507_
timestamp 1676037725
transform 1 0 33856 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1508_
timestamp 1676037725
transform 1 0 27140 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1509_
timestamp 1676037725
transform 1 0 26680 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1510_
timestamp 1676037725
transform 1 0 20516 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1511_
timestamp 1676037725
transform 1 0 27324 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1512_
timestamp 1676037725
transform 1 0 22264 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1513_
timestamp 1676037725
transform 1 0 22908 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1514_
timestamp 1676037725
transform 1 0 20792 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1515_
timestamp 1676037725
transform 1 0 20056 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1516_
timestamp 1676037725
transform 1 0 21988 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1517_
timestamp 1676037725
transform 1 0 27140 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1518_
timestamp 1676037725
transform 1 0 26128 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1519_
timestamp 1676037725
transform 1 0 31096 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1520_
timestamp 1676037725
transform 1 0 37444 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1521_
timestamp 1676037725
transform 1 0 37444 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1522_
timestamp 1676037725
transform 1 0 37444 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1523_
timestamp 1676037725
transform 1 0 37444 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1524_
timestamp 1676037725
transform 1 0 37444 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1525_
timestamp 1676037725
transform 1 0 37444 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1526_
timestamp 1676037725
transform 1 0 37444 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1527_
timestamp 1676037725
transform 1 0 16192 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1528_
timestamp 1676037725
transform 1 0 14720 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1529_
timestamp 1676037725
transform 1 0 15640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1530_
timestamp 1676037725
transform 1 0 15272 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1531_
timestamp 1676037725
transform 1 0 15272 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1532_
timestamp 1676037725
transform 1 0 14904 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1533_
timestamp 1676037725
transform 1 0 14076 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1534_
timestamp 1676037725
transform 1 0 14260 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1535_
timestamp 1676037725
transform 1 0 17388 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1536_
timestamp 1676037725
transform 1 0 16560 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1537_
timestamp 1676037725
transform 1 0 18308 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1538_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1539_
timestamp 1676037725
transform 1 0 21528 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1540_
timestamp 1676037725
transform 1 0 21988 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1541_
timestamp 1676037725
transform 1 0 22448 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1542_
timestamp 1676037725
transform 1 0 19780 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1543_
timestamp 1676037725
transform 1 0 19320 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1544_
timestamp 1676037725
transform 1 0 18124 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1545_
timestamp 1676037725
transform 1 0 16928 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1546_
timestamp 1676037725
transform 1 0 17940 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1547_
timestamp 1676037725
transform 1 0 20516 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1548_
timestamp 1676037725
transform 1 0 19320 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1549_
timestamp 1676037725
transform 1 0 12972 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1550_
timestamp 1676037725
transform 1 0 15088 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1551_
timestamp 1676037725
transform 1 0 13892 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1552_
timestamp 1676037725
transform 1 0 12696 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1553_
timestamp 1676037725
transform 1 0 12328 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1554_
timestamp 1676037725
transform 1 0 20608 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _1555_
timestamp 1676037725
transform 1 0 18952 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1556_
timestamp 1676037725
transform 1 0 19780 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1557_
timestamp 1676037725
transform 1 0 20056 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1558_
timestamp 1676037725
transform 1 0 21252 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1559_
timestamp 1676037725
transform 1 0 19688 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1560_
timestamp 1676037725
transform 1 0 14720 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1561_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1562_
timestamp 1676037725
transform 1 0 9108 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1563_
timestamp 1676037725
transform 1 0 10212 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1564_
timestamp 1676037725
transform 1 0 10396 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1565_
timestamp 1676037725
transform 1 0 14628 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1566_
timestamp 1676037725
transform 1 0 15456 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1567_
timestamp 1676037725
transform 1 0 16100 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1568_
timestamp 1676037725
transform 1 0 23184 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1569_
timestamp 1676037725
transform 1 0 6532 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1570_
timestamp 1676037725
transform 1 0 5060 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1571_
timestamp 1676037725
transform 1 0 7084 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1572_
timestamp 1676037725
transform 1 0 11684 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1573_
timestamp 1676037725
transform 1 0 9568 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1574_
timestamp 1676037725
transform 1 0 9108 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1575_
timestamp 1676037725
transform 1 0 12604 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1576_
timestamp 1676037725
transform 1 0 21988 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1577_
timestamp 1676037725
transform 1 0 26404 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1578_
timestamp 1676037725
transform 1 0 26312 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _1579_
timestamp 1676037725
transform 1 0 11776 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1580_
timestamp 1676037725
transform 1 0 6716 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _1581_
timestamp 1676037725
transform 1 0 7820 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1582_
timestamp 1676037725
transform 1 0 5796 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1583_
timestamp 1676037725
transform 1 0 8188 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1584_
timestamp 1676037725
transform 1 0 5152 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1585_
timestamp 1676037725
transform 1 0 4692 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1586_
timestamp 1676037725
transform 1 0 4876 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1587_
timestamp 1676037725
transform 1 0 7820 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1588_
timestamp 1676037725
transform 1 0 7544 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1589_
timestamp 1676037725
transform 1 0 4232 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1590_
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _1591_
timestamp 1676037725
transform 1 0 6808 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1592_
timestamp 1676037725
transform 1 0 5060 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1593_
timestamp 1676037725
transform 1 0 5060 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1594_
timestamp 1676037725
transform 1 0 3864 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1595_
timestamp 1676037725
transform 1 0 28152 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1596_
timestamp 1676037725
transform 1 0 3220 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _1597_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4784 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1598_
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1599_
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1600_
timestamp 1676037725
transform 1 0 13248 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1601_
timestamp 1676037725
transform 1 0 13156 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1602_
timestamp 1676037725
transform 1 0 5520 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1603_
timestamp 1676037725
transform 1 0 5520 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1604_
timestamp 1676037725
transform 1 0 4508 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1605_
timestamp 1676037725
transform 1 0 3956 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1606_
timestamp 1676037725
transform 1 0 6532 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1607_
timestamp 1676037725
transform 1 0 6532 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1608_
timestamp 1676037725
transform 1 0 6256 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1609_
timestamp 1676037725
transform 1 0 4692 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1610_
timestamp 1676037725
transform 1 0 3956 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1611_
timestamp 1676037725
transform 1 0 4048 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1612_
timestamp 1676037725
transform 1 0 3956 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1613_
timestamp 1676037725
transform 1 0 8372 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1614_
timestamp 1676037725
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1615_
timestamp 1676037725
transform 1 0 9108 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1616_
timestamp 1676037725
transform 1 0 10396 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1617_
timestamp 1676037725
transform 1 0 5152 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1618_
timestamp 1676037725
transform 1 0 3956 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1619_
timestamp 1676037725
transform 1 0 10212 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1620_
timestamp 1676037725
transform 1 0 8924 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1621_
timestamp 1676037725
transform 1 0 3956 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1622_
timestamp 1676037725
transform 1 0 7544 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1623_
timestamp 1676037725
transform 1 0 6532 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1624_
timestamp 1676037725
transform 1 0 9844 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1625_
timestamp 1676037725
transform 1 0 9384 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1626_
timestamp 1676037725
transform 1 0 7912 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1627_
timestamp 1676037725
transform 1 0 10672 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1628_
timestamp 1676037725
transform 1 0 9016 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1629_
timestamp 1676037725
transform 1 0 11500 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1630_
timestamp 1676037725
transform 1 0 6900 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1631_
timestamp 1676037725
transform 1 0 6624 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1632_
timestamp 1676037725
transform 1 0 6532 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1633_
timestamp 1676037725
transform 1 0 9200 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1634_
timestamp 1676037725
transform 1 0 8372 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1635_
timestamp 1676037725
transform 1 0 11776 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1636_
timestamp 1676037725
transform 1 0 9568 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1637_
timestamp 1676037725
transform 1 0 7176 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1638_
timestamp 1676037725
transform 1 0 10028 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1639_
timestamp 1676037725
transform 1 0 6900 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1640_
timestamp 1676037725
transform 1 0 6532 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_2  _1641_
timestamp 1676037725
transform 1 0 6992 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1642_
timestamp 1676037725
transform 1 0 7820 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _1643_
timestamp 1676037725
transform 1 0 7176 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1644_
timestamp 1676037725
transform 1 0 8280 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1645_
timestamp 1676037725
transform 1 0 7636 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1646_
timestamp 1676037725
transform 1 0 7728 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1647_
timestamp 1676037725
transform 1 0 6532 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1648_
timestamp 1676037725
transform 1 0 8004 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1649_
timestamp 1676037725
transform 1 0 8096 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1650_
timestamp 1676037725
transform 1 0 5060 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _1651_
timestamp 1676037725
transform 1 0 6256 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1652_
timestamp 1676037725
transform 1 0 9292 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1653_
timestamp 1676037725
transform 1 0 10120 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1654_
timestamp 1676037725
transform 1 0 10488 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _1655_
timestamp 1676037725
transform 1 0 9108 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1656_
timestamp 1676037725
transform 1 0 10488 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1657_
timestamp 1676037725
transform 1 0 10028 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1658_
timestamp 1676037725
transform 1 0 8004 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1659_
timestamp 1676037725
transform 1 0 10212 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1660_
timestamp 1676037725
transform 1 0 9384 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1661_
timestamp 1676037725
transform 1 0 14260 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1662_
timestamp 1676037725
transform 1 0 13984 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1663_
timestamp 1676037725
transform 1 0 29716 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1664_
timestamp 1676037725
transform 1 0 28796 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1665_
timestamp 1676037725
transform 1 0 30544 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1666_
timestamp 1676037725
transform 1 0 37444 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1667_
timestamp 1676037725
transform 1 0 37444 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1668_
timestamp 1676037725
transform 1 0 37444 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1669_
timestamp 1676037725
transform 1 0 37444 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1670_
timestamp 1676037725
transform 1 0 37444 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1671_
timestamp 1676037725
transform 1 0 36156 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1672_
timestamp 1676037725
transform 1 0 37444 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1673_
timestamp 1676037725
transform 1 0 29072 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1674_
timestamp 1676037725
transform 1 0 24564 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1675_
timestamp 1676037725
transform 1 0 30452 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1676_
timestamp 1676037725
transform 1 0 24564 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1677_
timestamp 1676037725
transform 1 0 35604 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1678_
timestamp 1676037725
transform 1 0 32292 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1679_
timestamp 1676037725
transform 1 0 37444 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1680_
timestamp 1676037725
transform 1 0 37444 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1681_
timestamp 1676037725
transform 1 0 27968 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1682_
timestamp 1676037725
transform 1 0 29992 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1683_
timestamp 1676037725
transform 1 0 24748 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1684_
timestamp 1676037725
transform 1 0 27876 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1685_
timestamp 1676037725
transform 1 0 23000 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1686_
timestamp 1676037725
transform 1 0 37444 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1687_
timestamp 1676037725
transform 1 0 32568 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1688_
timestamp 1676037725
transform 1 0 37444 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1689_
timestamp 1676037725
transform 1 0 37444 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1690_
timestamp 1676037725
transform 1 0 28888 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1691_
timestamp 1676037725
transform 1 0 14720 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1692_
timestamp 1676037725
transform 1 0 16836 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1693_
timestamp 1676037725
transform 1 0 16836 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1694_
timestamp 1676037725
transform 1 0 19412 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1695_
timestamp 1676037725
transform 1 0 26220 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1696_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1697_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13340 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1698_
timestamp 1676037725
transform 1 0 15364 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1699_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15824 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1700_
timestamp 1676037725
transform 1 0 17756 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1701_
timestamp 1676037725
transform 1 0 23920 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _1702_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24472 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1703_
timestamp 1676037725
transform 1 0 29716 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1704_
timestamp 1676037725
transform 1 0 25576 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1705_
timestamp 1676037725
transform 1 0 32292 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1706_
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1707_
timestamp 1676037725
transform 1 0 33580 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1708_
timestamp 1676037725
transform 1 0 32384 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1709_
timestamp 1676037725
transform 1 0 26496 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1710_
timestamp 1676037725
transform 1 0 24564 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1711_
timestamp 1676037725
transform 1 0 27416 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1712_
timestamp 1676037725
transform 1 0 22448 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1713_
timestamp 1676037725
transform 1 0 34776 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 1676037725
transform 1 0 30360 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 1676037725
transform 1 0 34868 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1716_
timestamp 1676037725
transform 1 0 32936 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1717_
timestamp 1676037725
transform 1 0 26680 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1718_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9476 0 -1 13056
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1719_
timestamp 1676037725
transform 1 0 9108 0 1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 1676037725
transform 1 0 21620 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1721_
timestamp 1676037725
transform 1 0 14168 0 -1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1722_
timestamp 1676037725
transform 1 0 15916 0 1 4352
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1723_
timestamp 1676037725
transform 1 0 19688 0 -1 5440
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1724_
timestamp 1676037725
transform 1 0 18124 0 -1 4352
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1725_
timestamp 1676037725
transform 1 0 20884 0 1 5440
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1726_
timestamp 1676037725
transform 1 0 11684 0 -1 7616
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1727_
timestamp 1676037725
transform 1 0 12972 0 -1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1728_
timestamp 1676037725
transform 1 0 7636 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1729_
timestamp 1676037725
transform 1 0 7912 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1730_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25852 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1731_
timestamp 1676037725
transform 1 0 33856 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1732_
timestamp 1676037725
transform 1 0 35696 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1733_
timestamp 1676037725
transform 1 0 34960 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1734_
timestamp 1676037725
transform 1 0 34868 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1735_
timestamp 1676037725
transform 1 0 34868 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1736_
timestamp 1676037725
transform 1 0 34868 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1737_
timestamp 1676037725
transform 1 0 32660 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1738_
timestamp 1676037725
transform 1 0 33856 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1739_
timestamp 1676037725
transform 1 0 33304 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1740_
timestamp 1676037725
transform 1 0 33764 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1741_
timestamp 1676037725
transform 1 0 32752 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1742_
timestamp 1676037725
transform 1 0 34132 0 -1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1743_
timestamp 1676037725
transform 1 0 34868 0 1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1744_
timestamp 1676037725
transform 1 0 34224 0 -1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1745_
timestamp 1676037725
transform 1 0 32292 0 -1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1746_
timestamp 1676037725
transform 1 0 30360 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1747_
timestamp 1676037725
transform 1 0 36892 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1748_
timestamp 1676037725
transform 1 0 36800 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1749_
timestamp 1676037725
transform 1 0 36708 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1750_
timestamp 1676037725
transform 1 0 36708 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1751_
timestamp 1676037725
transform 1 0 36892 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1752_
timestamp 1676037725
transform 1 0 36708 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1753_
timestamp 1676037725
transform 1 0 36800 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1754_
timestamp 1676037725
transform 1 0 12144 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1755_
timestamp 1676037725
transform 1 0 19964 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1756_
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1757_
timestamp 1676037725
transform 1 0 18216 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1758_
timestamp 1676037725
transform 1 0 19412 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1759_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1760_
timestamp 1676037725
transform 1 0 19780 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1761_
timestamp 1676037725
transform 1 0 16192 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1762_
timestamp 1676037725
transform 1 0 4416 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1763_
timestamp 1676037725
transform 1 0 4324 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1764_
timestamp 1676037725
transform 1 0 6348 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1765_
timestamp 1676037725
transform 1 0 10488 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1766_
timestamp 1676037725
transform 1 0 9108 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1767_
timestamp 1676037725
transform 1 0 7912 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1768_
timestamp 1676037725
transform 1 0 12052 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1769_
timestamp 1676037725
transform 1 0 21988 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1770_
timestamp 1676037725
transform 1 0 26036 0 1 35904
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1771_
timestamp 1676037725
transform 1 0 3956 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1772_
timestamp 1676037725
transform 1 0 27508 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1773_
timestamp 1676037725
transform 1 0 13156 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1774_
timestamp 1676037725
transform 1 0 2668 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1775_
timestamp 1676037725
transform 1 0 2668 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1776_
timestamp 1676037725
transform 1 0 2760 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1777_
timestamp 1676037725
transform 1 0 10580 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1778_
timestamp 1676037725
transform 1 0 2852 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1779_
timestamp 1676037725
transform 1 0 9108 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1780_
timestamp 1676037725
transform 1 0 2760 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1781_
timestamp 1676037725
transform 1 0 4508 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1782_
timestamp 1676037725
transform 1 0 9568 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1783_
timestamp 1676037725
transform 1 0 10488 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1784_
timestamp 1676037725
transform 1 0 12144 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1785_
timestamp 1676037725
transform 1 0 6532 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1786_
timestamp 1676037725
transform 1 0 7912 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1787_
timestamp 1676037725
transform 1 0 12052 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1788_
timestamp 1676037725
transform 1 0 9752 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1789_
timestamp 1676037725
transform 1 0 6716 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1790_
timestamp 1676037725
transform 1 0 5612 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1791_
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1792_
timestamp 1676037725
transform 1 0 4232 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1793_
timestamp 1676037725
transform 1 0 5796 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1794_
timestamp 1676037725
transform 1 0 10672 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1795_
timestamp 1676037725
transform 1 0 11500 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1796_
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1797_
timestamp 1676037725
transform 1 0 7912 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1798_
timestamp 1676037725
transform 1 0 11224 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1799_
timestamp 1676037725
transform 1 0 9384 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1800_
timestamp 1676037725
transform 1 0 14076 0 -1 25024
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1801_
timestamp 1676037725
transform 1 0 14260 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1802_
timestamp 1676037725
transform 1 0 16928 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1803_
timestamp 1676037725
transform 1 0 12328 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1804_
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1805_
timestamp 1676037725
transform 1 0 29440 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1806_
timestamp 1676037725
transform 1 0 28612 0 -1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1807_
timestamp 1676037725
transform 1 0 29992 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1808_
timestamp 1676037725
transform 1 0 36708 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1809_
timestamp 1676037725
transform 1 0 36800 0 1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1810_
timestamp 1676037725
transform 1 0 36800 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1811_
timestamp 1676037725
transform 1 0 36340 0 1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1812_
timestamp 1676037725
transform 1 0 36800 0 1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1813_
timestamp 1676037725
transform 1 0 36248 0 1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1814_
timestamp 1676037725
transform 1 0 36800 0 1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1815_
timestamp 1676037725
transform 1 0 22724 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1816_
timestamp 1676037725
transform 1 0 30452 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1817_
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1818_
timestamp 1676037725
transform 1 0 35236 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1819_
timestamp 1676037725
transform 1 0 31188 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1820_
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1821_
timestamp 1676037725
transform 1 0 36708 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1822_
timestamp 1676037725
transform 1 0 27324 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1823_
timestamp 1676037725
transform 1 0 22908 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1676037725
transform 1 0 27416 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1676037725
transform 1 0 22172 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1676037725
transform 1 0 32476 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1828_
timestamp 1676037725
transform 1 0 36800 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1676037725
transform 1 0 36708 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1676037725
transform 1 0 28704 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20516 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7636 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1676037725
transform 1 0 7360 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1676037725
transform 1 0 12144 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1676037725
transform 1 0 12512 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1676037725
transform 1 0 8188 0 -1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1676037725
transform 1 0 9108 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1676037725
transform 1 0 13616 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1676037725
transform 1 0 14260 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1676037725
transform 1 0 26220 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1676037725
transform 1 0 26128 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1676037725
transform 1 0 33212 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1676037725
transform 1 0 33120 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1676037725
transform 1 0 30728 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1676037725
transform 1 0 31004 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1676037725
transform 1 0 35236 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1676037725
transform 1 0 34868 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31740 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout39 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37628 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31188 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36064 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 1676037725
transform 1 0 15824 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout43
timestamp 1676037725
transform 1 0 30084 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  fanout44 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17480 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  fanout45
timestamp 1676037725
transform 1 0 25760 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout46
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout47
timestamp 1676037725
transform 1 0 5152 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout48
timestamp 1676037725
transform 1 0 28244 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout49
timestamp 1676037725
transform 1 0 20976 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout50
timestamp 1676037725
transform 1 0 10304 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout51
timestamp 1676037725
transform 1 0 27600 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout52
timestamp 1676037725
transform 1 0 7176 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout53
timestamp 1676037725
transform 1 0 24564 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout54
timestamp 1676037725
transform 1 0 27232 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout55
timestamp 1676037725
transform 1 0 11684 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout56
timestamp 1676037725
transform 1 0 10396 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout57
timestamp 1676037725
transform 1 0 14352 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout58
timestamp 1676037725
transform 1 0 15272 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout59
timestamp 1676037725
transform 1 0 16008 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout60
timestamp 1676037725
transform 1 0 27140 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout61
timestamp 1676037725
transform 1 0 9292 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout62
timestamp 1676037725
transform 1 0 14260 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout63
timestamp 1676037725
transform 1 0 12880 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  fanout64
timestamp 1676037725
transform 1 0 20056 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_8  fanout65
timestamp 1676037725
transform 1 0 16836 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout66
timestamp 1676037725
transform 1 0 24748 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout67
timestamp 1676037725
transform 1 0 24656 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout68
timestamp 1676037725
transform 1 0 28980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout69
timestamp 1676037725
transform 1 0 29624 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  fanout70
timestamp 1676037725
transform 1 0 9108 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_12  fanout71
timestamp 1676037725
transform 1 0 28520 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  fanout72
timestamp 1676037725
transform 1 0 6992 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout73
timestamp 1676037725
transform 1 0 22816 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout74
timestamp 1676037725
transform 1 0 27416 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout75 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25024 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  fanout76
timestamp 1676037725
transform 1 0 25116 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_6  fanout77
timestamp 1676037725
transform 1 0 27324 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout78
timestamp 1676037725
transform 1 0 27416 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout79
timestamp 1676037725
transform 1 0 15456 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout80
timestamp 1676037725
transform 1 0 20424 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout81
timestamp 1676037725
transform 1 0 20240 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout82
timestamp 1676037725
transform 1 0 22080 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout83
timestamp 1676037725
transform 1 0 18768 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout84
timestamp 1676037725
transform 1 0 23460 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout85
timestamp 1676037725
transform 1 0 18400 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout86
timestamp 1676037725
transform 1 0 17388 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_2  fanout87 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23644 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout88
timestamp 1676037725
transform 1 0 23552 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout89
timestamp 1676037725
transform 1 0 17664 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  input1
timestamp 1676037725
transform 1 0 1840 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input2
timestamp 1676037725
transform 1 0 4968 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  input3
timestamp 1676037725
transform 1 0 7820 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  input4
timestamp 1676037725
transform 1 0 11776 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  input5
timestamp 1676037725
transform 1 0 15088 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input6
timestamp 1676037725
transform 1 0 18124 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  input7
timestamp 1676037725
transform 1 0 21988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  input8
timestamp 1676037725
transform 1 0 25024 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1676037725
transform 1 0 28336 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1676037725
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input11
timestamp 1676037725
transform 1 0 37536 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  output12
timestamp 1676037725
transform 1 0 36432 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output13
timestamp 1676037725
transform 1 0 37812 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output14
timestamp 1676037725
transform 1 0 37812 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output15
timestamp 1676037725
transform 1 0 37812 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output16
timestamp 1676037725
transform 1 0 37812 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output17
timestamp 1676037725
transform 1 0 37812 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output18
timestamp 1676037725
transform 1 0 37812 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output19
timestamp 1676037725
transform 1 0 37812 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output20
timestamp 1676037725
transform 1 0 37812 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output21
timestamp 1676037725
transform 1 0 37812 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output22
timestamp 1676037725
transform 1 0 37812 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output23
timestamp 1676037725
transform 1 0 36892 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output24
timestamp 1676037725
transform 1 0 37812 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output25
timestamp 1676037725
transform 1 0 37444 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output26
timestamp 1676037725
transform 1 0 36708 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output27
timestamp 1676037725
transform 1 0 37812 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output28
timestamp 1676037725
transform 1 0 37812 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output29
timestamp 1676037725
transform 1 0 37812 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output30
timestamp 1676037725
transform 1 0 37812 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output31
timestamp 1676037725
transform 1 0 36432 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output32
timestamp 1676037725
transform 1 0 37812 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output33
timestamp 1676037725
transform 1 0 37812 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output34
timestamp 1676037725
transform 1 0 37812 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output35
timestamp 1676037725
transform 1 0 37812 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output36
timestamp 1676037725
transform 1 0 37812 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output37
timestamp 1676037725
transform 1 0 37812 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  wrapped_6502_90 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38088 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wrapped_6502_91
timestamp 1676037725
transform 1 0 38088 0 -1 14144
box -38 -48 314 592
<< labels >>
flabel metal2 s 34886 39200 34942 40000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 1766 39200 1822 40000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 5078 39200 5134 40000 0 FreeSans 224 90 0 0 io_in[1]
port 2 nsew signal input
flabel metal2 s 8390 39200 8446 40000 0 FreeSans 224 90 0 0 io_in[2]
port 3 nsew signal input
flabel metal2 s 11702 39200 11758 40000 0 FreeSans 224 90 0 0 io_in[3]
port 4 nsew signal input
flabel metal2 s 15014 39200 15070 40000 0 FreeSans 224 90 0 0 io_in[4]
port 5 nsew signal input
flabel metal2 s 18326 39200 18382 40000 0 FreeSans 224 90 0 0 io_in[5]
port 6 nsew signal input
flabel metal2 s 21638 39200 21694 40000 0 FreeSans 224 90 0 0 io_in[6]
port 7 nsew signal input
flabel metal2 s 24950 39200 25006 40000 0 FreeSans 224 90 0 0 io_in[7]
port 8 nsew signal input
flabel metal2 s 28262 39200 28318 40000 0 FreeSans 224 90 0 0 io_in[8]
port 9 nsew signal input
flabel metal2 s 31574 39200 31630 40000 0 FreeSans 224 90 0 0 io_in[9]
port 10 nsew signal input
flabel metal3 s 39200 38224 40000 38344 0 FreeSans 480 0 0 0 io_oeb
port 11 nsew signal tristate
flabel metal3 s 39200 1504 40000 1624 0 FreeSans 480 0 0 0 io_out[0]
port 12 nsew signal tristate
flabel metal3 s 39200 15104 40000 15224 0 FreeSans 480 0 0 0 io_out[10]
port 13 nsew signal tristate
flabel metal3 s 39200 16464 40000 16584 0 FreeSans 480 0 0 0 io_out[11]
port 14 nsew signal tristate
flabel metal3 s 39200 17824 40000 17944 0 FreeSans 480 0 0 0 io_out[12]
port 15 nsew signal tristate
flabel metal3 s 39200 19184 40000 19304 0 FreeSans 480 0 0 0 io_out[13]
port 16 nsew signal tristate
flabel metal3 s 39200 20544 40000 20664 0 FreeSans 480 0 0 0 io_out[14]
port 17 nsew signal tristate
flabel metal3 s 39200 21904 40000 22024 0 FreeSans 480 0 0 0 io_out[15]
port 18 nsew signal tristate
flabel metal3 s 39200 23264 40000 23384 0 FreeSans 480 0 0 0 io_out[16]
port 19 nsew signal tristate
flabel metal3 s 39200 24624 40000 24744 0 FreeSans 480 0 0 0 io_out[17]
port 20 nsew signal tristate
flabel metal3 s 39200 25984 40000 26104 0 FreeSans 480 0 0 0 io_out[18]
port 21 nsew signal tristate
flabel metal3 s 39200 27344 40000 27464 0 FreeSans 480 0 0 0 io_out[19]
port 22 nsew signal tristate
flabel metal3 s 39200 2864 40000 2984 0 FreeSans 480 0 0 0 io_out[1]
port 23 nsew signal tristate
flabel metal3 s 39200 28704 40000 28824 0 FreeSans 480 0 0 0 io_out[20]
port 24 nsew signal tristate
flabel metal3 s 39200 30064 40000 30184 0 FreeSans 480 0 0 0 io_out[21]
port 25 nsew signal tristate
flabel metal3 s 39200 31424 40000 31544 0 FreeSans 480 0 0 0 io_out[22]
port 26 nsew signal tristate
flabel metal3 s 39200 32784 40000 32904 0 FreeSans 480 0 0 0 io_out[23]
port 27 nsew signal tristate
flabel metal3 s 39200 34144 40000 34264 0 FreeSans 480 0 0 0 io_out[24]
port 28 nsew signal tristate
flabel metal3 s 39200 35504 40000 35624 0 FreeSans 480 0 0 0 io_out[25]
port 29 nsew signal tristate
flabel metal3 s 39200 36864 40000 36984 0 FreeSans 480 0 0 0 io_out[26]
port 30 nsew signal tristate
flabel metal3 s 39200 4224 40000 4344 0 FreeSans 480 0 0 0 io_out[2]
port 31 nsew signal tristate
flabel metal3 s 39200 5584 40000 5704 0 FreeSans 480 0 0 0 io_out[3]
port 32 nsew signal tristate
flabel metal3 s 39200 6944 40000 7064 0 FreeSans 480 0 0 0 io_out[4]
port 33 nsew signal tristate
flabel metal3 s 39200 8304 40000 8424 0 FreeSans 480 0 0 0 io_out[5]
port 34 nsew signal tristate
flabel metal3 s 39200 9664 40000 9784 0 FreeSans 480 0 0 0 io_out[6]
port 35 nsew signal tristate
flabel metal3 s 39200 11024 40000 11144 0 FreeSans 480 0 0 0 io_out[7]
port 36 nsew signal tristate
flabel metal3 s 39200 12384 40000 12504 0 FreeSans 480 0 0 0 io_out[8]
port 37 nsew signal tristate
flabel metal3 s 39200 13744 40000 13864 0 FreeSans 480 0 0 0 io_out[9]
port 38 nsew signal tristate
flabel metal2 s 38198 39200 38254 40000 0 FreeSans 224 90 0 0 rst
port 39 nsew signal input
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
