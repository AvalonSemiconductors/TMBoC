magic
tech sky130B
magscale 1 2
timestamp 1683541606
<< obsli1 >>
rect 1104 2159 16836 15793
<< obsm1 >>
rect 842 892 17098 17332
<< metal2 >>
rect 4434 17200 4490 18000
rect 13450 17200 13506 18000
rect 846 0 902 800
rect 2318 0 2374 800
rect 3790 0 3846 800
rect 5262 0 5318 800
rect 6734 0 6790 800
rect 8206 0 8262 800
rect 9678 0 9734 800
rect 11150 0 11206 800
rect 12622 0 12678 800
rect 14094 0 14150 800
rect 15566 0 15622 800
rect 17038 0 17094 800
<< obsm2 >>
rect 848 17144 4378 17354
rect 4546 17144 13394 17354
rect 13562 17144 17092 17354
rect 848 856 17092 17144
rect 958 734 2262 856
rect 2430 734 3734 856
rect 3902 734 5206 856
rect 5374 734 6678 856
rect 6846 734 8150 856
rect 8318 734 9622 856
rect 9790 734 11094 856
rect 11262 734 12566 856
rect 12734 734 14038 856
rect 14206 734 15510 856
rect 15678 734 16982 856
<< obsm3 >>
rect 2912 2143 16993 15809
<< metal4 >>
rect 2910 2128 3230 15824
rect 4876 2128 5196 15824
rect 6843 2128 7163 15824
rect 8809 2128 9129 15824
rect 10776 2128 11096 15824
rect 12742 2128 13062 15824
rect 14709 2128 15029 15824
rect 16675 2128 16995 15824
<< labels >>
rlabel metal2 s 4434 17200 4490 18000 6 clk
port 1 nsew signal input
rlabel metal2 s 846 0 902 800 6 io_out[0]
port 2 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 io_out[10]
port 3 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 io_out[11]
port 4 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 io_out[1]
port 5 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 io_out[2]
port 6 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 io_out[3]
port 7 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 io_out[4]
port 8 nsew signal output
rlabel metal2 s 8206 0 8262 800 6 io_out[5]
port 9 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 io_out[6]
port 10 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 io_out[7]
port 11 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 io_out[8]
port 12 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 io_out[9]
port 13 nsew signal output
rlabel metal2 s 13450 17200 13506 18000 6 rst
port 14 nsew signal input
rlabel metal4 s 2910 2128 3230 15824 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 6843 2128 7163 15824 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 10776 2128 11096 15824 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 14709 2128 15029 15824 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 4876 2128 5196 15824 6 vssd1
port 16 nsew ground bidirectional
rlabel metal4 s 8809 2128 9129 15824 6 vssd1
port 16 nsew ground bidirectional
rlabel metal4 s 12742 2128 13062 15824 6 vssd1
port 16 nsew ground bidirectional
rlabel metal4 s 16675 2128 16995 15824 6 vssd1
port 16 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 18000 18000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 726936
string GDS_FILE /media/lucah/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/MultiplexedCounter/runs/23_05_08_12_25/results/signoff/tt2_tholin_multiplexed_counter.magic.gds
string GDS_START 270124
<< end >>

