// This is the unpowered netlist.
module posit_unit (clk,
    rst,
    io_in,
    io_out);
 input clk;
 input rst;
 input [2:0] io_in;
 output [3:0] io_out;

 wire net243;
 wire net244;
 wire net245;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire \cmd[0] ;
 wire \cmd[6] ;
 wire \cmd[7] ;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \in_reg[0] ;
 wire \in_reg[10] ;
 wire \in_reg[11] ;
 wire \in_reg[12] ;
 wire \in_reg[13] ;
 wire \in_reg[14] ;
 wire \in_reg[15] ;
 wire \in_reg[1] ;
 wire \in_reg[2] ;
 wire \in_reg[3] ;
 wire \in_reg[4] ;
 wire \in_reg[5] ;
 wire \in_reg[6] ;
 wire \in_reg[7] ;
 wire \in_reg[8] ;
 wire \in_reg[9] ;
 wire last_SCLK;
 wire mode;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \out_reg[0] ;
 wire \out_reg[10] ;
 wire \out_reg[11] ;
 wire \out_reg[12] ;
 wire \out_reg[13] ;
 wire \out_reg[14] ;
 wire \out_reg[15] ;
 wire \out_reg[1] ;
 wire \out_reg[2] ;
 wire \out_reg[3] ;
 wire \out_reg[4] ;
 wire \out_reg[5] ;
 wire \out_reg[6] ;
 wire \out_reg[7] ;
 wire \out_reg[8] ;
 wire \out_reg[9] ;
 wire \posit_add.in1[0] ;
 wire \posit_add.in1[10] ;
 wire \posit_add.in1[11] ;
 wire \posit_add.in1[12] ;
 wire \posit_add.in1[13] ;
 wire \posit_add.in1[14] ;
 wire \posit_add.in1[15] ;
 wire \posit_add.in1[1] ;
 wire \posit_add.in1[2] ;
 wire \posit_add.in1[3] ;
 wire \posit_add.in1[4] ;
 wire \posit_add.in1[5] ;
 wire \posit_add.in1[6] ;
 wire \posit_add.in1[7] ;
 wire \posit_add.in1[8] ;
 wire \posit_add.in1[9] ;
 wire \posit_add.in2[0] ;
 wire \posit_add.in2[10] ;
 wire \posit_add.in2[11] ;
 wire \posit_add.in2[12] ;
 wire \posit_add.in2[13] ;
 wire \posit_add.in2[14] ;
 wire \posit_add.in2[15] ;
 wire \posit_add.in2[1] ;
 wire \posit_add.in2[2] ;
 wire \posit_add.in2[3] ;
 wire \posit_add.in2[4] ;
 wire \posit_add.in2[5] ;
 wire \posit_add.in2[6] ;
 wire \posit_add.in2[7] ;
 wire \posit_add.in2[8] ;
 wire \posit_add.in2[9] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_1230_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_1471_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_1645_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_3476_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_3476_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_3496_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net83));
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_96 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _4004_ (.A(mode),
    .Y(_0635_));
 sky130_fd_sc_hd__inv_2 _4005_ (.A(net234),
    .Y(_0646_));
 sky130_fd_sc_hd__inv_2 _4006_ (.A(\posit_add.in2[0] ),
    .Y(_0657_));
 sky130_fd_sc_hd__inv_2 _4007_ (.A(net231),
    .Y(_0668_));
 sky130_fd_sc_hd__or4_1 _4008_ (.A(\in_reg[5] ),
    .B(\in_reg[4] ),
    .C(\in_reg[7] ),
    .D(\in_reg[6] ),
    .X(_0679_));
 sky130_fd_sc_hd__or4_1 _4009_ (.A(\in_reg[1] ),
    .B(\in_reg[0] ),
    .C(\in_reg[3] ),
    .D(\in_reg[2] ),
    .X(_0690_));
 sky130_fd_sc_hd__or3_2 _4010_ (.A(\counter[2] ),
    .B(\counter[1] ),
    .C(\counter[0] ),
    .X(_0701_));
 sky130_fd_sc_hd__nor4b_4 _4011_ (.A(\counter[4] ),
    .B(mode),
    .C(_0701_),
    .D_N(\counter[3] ),
    .Y(_0712_));
 sky130_fd_sc_hd__o21ai_1 _4012_ (.A1(_0679_),
    .A2(_0690_),
    .B1(_0712_),
    .Y(_0723_));
 sky130_fd_sc_hd__or3b_4 _4013_ (.A(net238),
    .B(_0723_),
    .C_N(net240),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _4014_ (.A0(\in_reg[0] ),
    .A1(\cmd[0] ),
    .S(_0734_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _4015_ (.A0(\in_reg[6] ),
    .A1(\cmd[6] ),
    .S(_0734_),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _4016_ (.A0(\in_reg[7] ),
    .A1(\cmd[7] ),
    .S(_0734_),
    .X(_0002_));
 sky130_fd_sc_hd__and2b_4 _4017_ (.A_N(last_SCLK),
    .B(net2),
    .X(_0775_));
 sky130_fd_sc_hd__and2_2 _4018_ (.A(net239),
    .B(net228),
    .X(_0786_));
 sky130_fd_sc_hd__nand2_1 _4019_ (.A(net239),
    .B(_0775_),
    .Y(_0797_));
 sky130_fd_sc_hd__or2_2 _4020_ (.A(net238),
    .B(_0797_),
    .X(_0808_));
 sky130_fd_sc_hd__mux2_1 _4021_ (.A0(net3),
    .A1(\in_reg[0] ),
    .S(net217),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _4022_ (.A0(\in_reg[0] ),
    .A1(\in_reg[1] ),
    .S(net218),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _4023_ (.A0(\in_reg[1] ),
    .A1(\in_reg[2] ),
    .S(net217),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _4024_ (.A0(\in_reg[2] ),
    .A1(\in_reg[3] ),
    .S(net217),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _4025_ (.A0(\in_reg[3] ),
    .A1(\in_reg[4] ),
    .S(net217),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _4026_ (.A0(\in_reg[4] ),
    .A1(\in_reg[5] ),
    .S(net218),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _4027_ (.A0(\in_reg[5] ),
    .A1(\in_reg[6] ),
    .S(net218),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _4028_ (.A0(\in_reg[6] ),
    .A1(\in_reg[7] ),
    .S(net218),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _4029_ (.A0(\in_reg[7] ),
    .A1(\in_reg[8] ),
    .S(net217),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _4030_ (.A0(\in_reg[8] ),
    .A1(\in_reg[9] ),
    .S(net217),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _4031_ (.A0(\in_reg[9] ),
    .A1(\in_reg[10] ),
    .S(net217),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _4032_ (.A0(\in_reg[10] ),
    .A1(\in_reg[11] ),
    .S(net217),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _4033_ (.A0(\in_reg[11] ),
    .A1(\in_reg[12] ),
    .S(net217),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _4034_ (.A0(\in_reg[12] ),
    .A1(\in_reg[13] ),
    .S(net218),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _4035_ (.A0(\in_reg[13] ),
    .A1(\in_reg[14] ),
    .S(net218),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _4036_ (.A0(\in_reg[14] ),
    .A1(\in_reg[15] ),
    .S(net218),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _4037_ (.A0(last_SCLK),
    .A1(net2),
    .S(net240),
    .X(_0979_));
 sky130_fd_sc_hd__and2b_1 _4038_ (.A_N(net238),
    .B(_0979_),
    .X(_0019_));
 sky130_fd_sc_hd__or4_4 _4039_ (.A(net235),
    .B(\posit_add.in1[3] ),
    .C(\posit_add.in1[2] ),
    .D(\posit_add.in1[1] ),
    .X(_1000_));
 sky130_fd_sc_hd__or4_2 _4040_ (.A(\posit_add.in1[6] ),
    .B(\posit_add.in1[5] ),
    .C(\posit_add.in1[4] ),
    .D(_1000_),
    .X(_1011_));
 sky130_fd_sc_hd__or2_4 _4041_ (.A(\posit_add.in1[7] ),
    .B(_1011_),
    .X(_1022_));
 sky130_fd_sc_hd__or4_4 _4042_ (.A(\posit_add.in1[9] ),
    .B(\posit_add.in1[8] ),
    .C(\posit_add.in1[7] ),
    .D(_1011_),
    .X(_1033_));
 sky130_fd_sc_hd__or3_4 _4043_ (.A(\posit_add.in1[11] ),
    .B(\posit_add.in1[10] ),
    .C(_1033_),
    .X(_1044_));
 sky130_fd_sc_hd__or2_2 _4044_ (.A(\posit_add.in1[13] ),
    .B(\posit_add.in1[12] ),
    .X(_1055_));
 sky130_fd_sc_hd__o41a_1 _4045_ (.A1(\posit_add.in1[11] ),
    .A2(\posit_add.in1[10] ),
    .A3(_1033_),
    .A4(_1055_),
    .B1(net232),
    .X(_1066_));
 sky130_fd_sc_hd__xnor2_1 _4046_ (.A(\posit_add.in1[14] ),
    .B(_1066_),
    .Y(_1077_));
 sky130_fd_sc_hd__clkinv_8 _4047_ (.A(net204),
    .Y(_1088_));
 sky130_fd_sc_hd__nand2_8 _4048_ (.A(net233),
    .B(_1022_),
    .Y(_1099_));
 sky130_fd_sc_hd__xor2_4 _4049_ (.A(\posit_add.in1[8] ),
    .B(_1099_),
    .X(_1110_));
 sky130_fd_sc_hd__xnor2_4 _4050_ (.A(\posit_add.in1[8] ),
    .B(_1099_),
    .Y(_1121_));
 sky130_fd_sc_hd__and2_2 _4051_ (.A(net203),
    .B(_1110_),
    .X(_1132_));
 sky130_fd_sc_hd__and2_2 _4052_ (.A(net232),
    .B(_1011_),
    .X(_1143_));
 sky130_fd_sc_hd__xnor2_1 _4053_ (.A(\posit_add.in1[7] ),
    .B(_1143_),
    .Y(_1154_));
 sky130_fd_sc_hd__xor2_4 _4054_ (.A(\posit_add.in1[7] ),
    .B(_1143_),
    .X(_1165_));
 sky130_fd_sc_hd__nor2_2 _4055_ (.A(net203),
    .B(_1110_),
    .Y(_1176_));
 sky130_fd_sc_hd__mux2_4 _4056_ (.A0(_1132_),
    .A1(_1176_),
    .S(_1165_),
    .X(_1187_));
 sky130_fd_sc_hd__nand2_2 _4057_ (.A(net232),
    .B(_1033_),
    .Y(_1198_));
 sky130_fd_sc_hd__xnor2_4 _4058_ (.A(\posit_add.in1[10] ),
    .B(_1198_),
    .Y(_1209_));
 sky130_fd_sc_hd__xnor2_4 _4059_ (.A(net203),
    .B(_1209_),
    .Y(_1220_));
 sky130_fd_sc_hd__o21a_2 _4060_ (.A1(\posit_add.in1[8] ),
    .A2(_1022_),
    .B1(net233),
    .X(_1231_));
 sky130_fd_sc_hd__xor2_4 _4061_ (.A(\posit_add.in1[9] ),
    .B(_1231_),
    .X(_1242_));
 sky130_fd_sc_hd__xnor2_4 _4062_ (.A(net203),
    .B(_1242_),
    .Y(_1253_));
 sky130_fd_sc_hd__nor2_4 _4063_ (.A(_1220_),
    .B(_1253_),
    .Y(_1264_));
 sky130_fd_sc_hd__nand2_4 _4064_ (.A(_1187_),
    .B(_1264_),
    .Y(_1275_));
 sky130_fd_sc_hd__clkinv_2 _4065_ (.A(_1275_),
    .Y(_1286_));
 sky130_fd_sc_hd__nand2_2 _4066_ (.A(net232),
    .B(_1044_),
    .Y(_1297_));
 sky130_fd_sc_hd__o21a_2 _4067_ (.A1(\posit_add.in1[12] ),
    .A2(_1044_),
    .B1(net233),
    .X(_1308_));
 sky130_fd_sc_hd__xnor2_4 _4068_ (.A(\posit_add.in1[13] ),
    .B(_1308_),
    .Y(_1319_));
 sky130_fd_sc_hd__inv_2 _4069_ (.A(_1319_),
    .Y(_1330_));
 sky130_fd_sc_hd__xnor2_4 _4070_ (.A(_1088_),
    .B(_1319_),
    .Y(_1341_));
 sky130_fd_sc_hd__xnor2_4 _4071_ (.A(net203),
    .B(_1319_),
    .Y(_1352_));
 sky130_fd_sc_hd__xnor2_4 _4072_ (.A(\posit_add.in1[12] ),
    .B(_1297_),
    .Y(_1363_));
 sky130_fd_sc_hd__xnor2_4 _4073_ (.A(_1088_),
    .B(_1363_),
    .Y(_1374_));
 sky130_fd_sc_hd__xnor2_4 _4074_ (.A(net203),
    .B(_1363_),
    .Y(_1385_));
 sky130_fd_sc_hd__o21ai_4 _4075_ (.A1(\posit_add.in1[10] ),
    .A2(_1033_),
    .B1(net232),
    .Y(_1396_));
 sky130_fd_sc_hd__xnor2_4 _4076_ (.A(\posit_add.in1[11] ),
    .B(_1396_),
    .Y(_1407_));
 sky130_fd_sc_hd__xor2_4 _4077_ (.A(net203),
    .B(_1407_),
    .X(_1418_));
 sky130_fd_sc_hd__nand2_2 _4078_ (.A(_1374_),
    .B(_1418_),
    .Y(_1429_));
 sky130_fd_sc_hd__or2_4 _4079_ (.A(_1341_),
    .B(_1429_),
    .X(_1440_));
 sky130_fd_sc_hd__and3b_4 _4080_ (.A_N(_1440_),
    .B(_1022_),
    .C(_1286_),
    .X(_1451_));
 sky130_fd_sc_hd__or3b_4 _4081_ (.A(_1275_),
    .B(_1440_),
    .C_N(_1022_),
    .X(_1462_));
 sky130_fd_sc_hd__o21ai_4 _4082_ (.A1(net235),
    .A2(\posit_add.in1[1] ),
    .B1(net233),
    .Y(_1473_));
 sky130_fd_sc_hd__xnor2_4 _4083_ (.A(\posit_add.in1[2] ),
    .B(_1473_),
    .Y(_1484_));
 sky130_fd_sc_hd__xor2_1 _4084_ (.A(net204),
    .B(_1484_),
    .X(_1495_));
 sky130_fd_sc_hd__nand2_2 _4085_ (.A(\posit_add.in1[0] ),
    .B(net232),
    .Y(_1506_));
 sky130_fd_sc_hd__xnor2_4 _4086_ (.A(\posit_add.in1[1] ),
    .B(_1506_),
    .Y(_1517_));
 sky130_fd_sc_hd__xor2_1 _4087_ (.A(net204),
    .B(_1517_),
    .X(_1528_));
 sky130_fd_sc_hd__or4_1 _4088_ (.A(net235),
    .B(\posit_add.in1[2] ),
    .C(\posit_add.in1[1] ),
    .D(_1088_),
    .X(_1539_));
 sky130_fd_sc_hd__o31a_2 _4089_ (.A1(\posit_add.in1[5] ),
    .A2(\posit_add.in1[4] ),
    .A3(_1000_),
    .B1(net232),
    .X(_1550_));
 sky130_fd_sc_hd__xor2_4 _4090_ (.A(\posit_add.in1[6] ),
    .B(_1550_),
    .X(_1561_));
 sky130_fd_sc_hd__xor2_4 _4091_ (.A(net204),
    .B(_1561_),
    .X(_1572_));
 sky130_fd_sc_hd__o21ai_4 _4092_ (.A1(\posit_add.in1[4] ),
    .A2(_1000_),
    .B1(net232),
    .Y(_1583_));
 sky130_fd_sc_hd__xnor2_4 _4093_ (.A(\posit_add.in1[5] ),
    .B(_1583_),
    .Y(_1594_));
 sky130_fd_sc_hd__xor2_2 _4094_ (.A(net205),
    .B(_1594_),
    .X(_1605_));
 sky130_fd_sc_hd__nand2_1 _4095_ (.A(_1572_),
    .B(_1605_),
    .Y(_1616_));
 sky130_fd_sc_hd__nand2_2 _4096_ (.A(net232),
    .B(_1000_),
    .Y(_1627_));
 sky130_fd_sc_hd__xnor2_4 _4097_ (.A(\posit_add.in1[4] ),
    .B(_1627_),
    .Y(_1638_));
 sky130_fd_sc_hd__xnor2_2 _4098_ (.A(net204),
    .B(_1638_),
    .Y(_1649_));
 sky130_fd_sc_hd__o31a_2 _4099_ (.A1(net235),
    .A2(\posit_add.in1[2] ),
    .A3(\posit_add.in1[1] ),
    .B1(net232),
    .X(_1660_));
 sky130_fd_sc_hd__xor2_4 _4100_ (.A(\posit_add.in1[3] ),
    .B(_1660_),
    .X(_1671_));
 sky130_fd_sc_hd__xnor2_1 _4101_ (.A(net204),
    .B(_1671_),
    .Y(_1682_));
 sky130_fd_sc_hd__or2_1 _4102_ (.A(_1649_),
    .B(_1682_),
    .X(_1693_));
 sky130_fd_sc_hd__or3b_4 _4103_ (.A(_1616_),
    .B(_1693_),
    .C_N(_1539_),
    .X(_1704_));
 sky130_fd_sc_hd__a21oi_4 _4104_ (.A1(_1286_),
    .A2(_1704_),
    .B1(_1440_),
    .Y(_1715_));
 sky130_fd_sc_hd__a21o_4 _4105_ (.A1(_1286_),
    .A2(_1704_),
    .B1(_1440_),
    .X(_1726_));
 sky130_fd_sc_hd__o211a_1 _4106_ (.A1(net235),
    .A2(_1088_),
    .B1(_1495_),
    .C1(_1528_),
    .X(_1737_));
 sky130_fd_sc_hd__nor2_1 _4107_ (.A(_1693_),
    .B(_1737_),
    .Y(_1748_));
 sky130_fd_sc_hd__o21ai_2 _4108_ (.A1(_1616_),
    .A2(_1748_),
    .B1(_1187_),
    .Y(_1759_));
 sky130_fd_sc_hd__a21oi_4 _4109_ (.A1(_1264_),
    .A2(_1759_),
    .B1(_1429_),
    .Y(_1770_));
 sky130_fd_sc_hd__nor2_2 _4110_ (.A(_1341_),
    .B(_1770_),
    .Y(_1781_));
 sky130_fd_sc_hd__or2_1 _4111_ (.A(_1341_),
    .B(_1770_),
    .X(_1792_));
 sky130_fd_sc_hd__nand2b_1 _4112_ (.A_N(net235),
    .B(\posit_add.in1[1] ),
    .Y(_1803_));
 sky130_fd_sc_hd__mux2_1 _4113_ (.A0(_1803_),
    .A1(_1517_),
    .S(net204),
    .X(_1814_));
 sky130_fd_sc_hd__a21oi_1 _4114_ (.A1(_1495_),
    .A2(_1814_),
    .B1(_1682_),
    .Y(_1825_));
 sky130_fd_sc_hd__o21ai_2 _4115_ (.A1(_1649_),
    .A2(_1825_),
    .B1(_1605_),
    .Y(_1836_));
 sky130_fd_sc_hd__a21oi_4 _4116_ (.A1(_1572_),
    .A2(_1836_),
    .B1(_1275_),
    .Y(_1847_));
 sky130_fd_sc_hd__nor3_4 _4117_ (.A(_1132_),
    .B(_1176_),
    .C(_1253_),
    .Y(_1858_));
 sky130_fd_sc_hd__o31a_4 _4118_ (.A1(_1220_),
    .A2(_1847_),
    .A3(_1858_),
    .B1(_1418_),
    .X(_1869_));
 sky130_fd_sc_hd__o31ai_4 _4119_ (.A1(_1220_),
    .A2(_1847_),
    .A3(_1858_),
    .B1(_1418_),
    .Y(_1880_));
 sky130_fd_sc_hd__a21oi_4 _4120_ (.A1(_1374_),
    .A2(_1880_),
    .B1(_1341_),
    .Y(_1891_));
 sky130_fd_sc_hd__a21o_1 _4121_ (.A1(_1374_),
    .A2(_1880_),
    .B1(_1341_),
    .X(_1902_));
 sky130_fd_sc_hd__o211a_1 _4122_ (.A1(_1385_),
    .A2(_1869_),
    .B1(_1671_),
    .C1(_1352_),
    .X(_1913_));
 sky130_fd_sc_hd__o211a_1 _4123_ (.A1(_1385_),
    .A2(_1869_),
    .B1(_1594_),
    .C1(_1352_),
    .X(_1924_));
 sky130_fd_sc_hd__a211o_2 _4124_ (.A1(_1638_),
    .A2(net130),
    .B1(_1924_),
    .C1(_1781_),
    .X(_1935_));
 sky130_fd_sc_hd__a211o_2 _4125_ (.A1(_1484_),
    .A2(net130),
    .B1(_1913_),
    .C1(net131),
    .X(_1946_));
 sky130_fd_sc_hd__a211o_1 _4126_ (.A1(_1374_),
    .A2(_1880_),
    .B1(_1517_),
    .C1(_1341_),
    .X(_1957_));
 sky130_fd_sc_hd__o211a_1 _4127_ (.A1(_1385_),
    .A2(_1869_),
    .B1(_1517_),
    .C1(_1352_),
    .X(_1968_));
 sky130_fd_sc_hd__o2111a_1 _4128_ (.A1(net235),
    .A2(_1891_),
    .B1(_1957_),
    .C1(_1715_),
    .D1(net131),
    .X(_1979_));
 sky130_fd_sc_hd__a31o_4 _4129_ (.A1(net169),
    .A2(_1935_),
    .A3(_1946_),
    .B1(_1979_),
    .X(_1990_));
 sky130_fd_sc_hd__a211o_1 _4130_ (.A1(_1374_),
    .A2(_1880_),
    .B1(_1242_),
    .C1(_1341_),
    .X(_2001_));
 sky130_fd_sc_hd__o211a_1 _4131_ (.A1(_1121_),
    .A2(_1891_),
    .B1(_2001_),
    .C1(net132),
    .X(_2012_));
 sky130_fd_sc_hd__o211a_1 _4132_ (.A1(_1385_),
    .A2(_1869_),
    .B1(_1165_),
    .C1(_1352_),
    .X(_2023_));
 sky130_fd_sc_hd__a21o_1 _4133_ (.A1(_1561_),
    .A2(net129),
    .B1(_2023_),
    .X(_2034_));
 sky130_fd_sc_hd__a21o_1 _4134_ (.A1(net133),
    .A2(_2034_),
    .B1(_2012_),
    .X(_2045_));
 sky130_fd_sc_hd__a211o_1 _4135_ (.A1(_1374_),
    .A2(_1880_),
    .B1(_1407_),
    .C1(_1341_),
    .X(_2056_));
 sky130_fd_sc_hd__o21a_1 _4136_ (.A1(_1209_),
    .A2(_1891_),
    .B1(_2056_),
    .X(_2067_));
 sky130_fd_sc_hd__mux2_1 _4137_ (.A0(_1363_),
    .A1(_2067_),
    .S(net133),
    .X(_2078_));
 sky130_fd_sc_hd__mux2_1 _4138_ (.A0(_2045_),
    .A1(_2078_),
    .S(_1726_),
    .X(_2089_));
 sky130_fd_sc_hd__mux2_8 _4139_ (.A0(_1990_),
    .A1(_2089_),
    .S(net171),
    .X(_2100_));
 sky130_fd_sc_hd__or2_4 _4140_ (.A(\posit_add.in2[0] ),
    .B(\posit_add.in2[1] ),
    .X(_2111_));
 sky130_fd_sc_hd__or4_4 _4141_ (.A(\posit_add.in2[0] ),
    .B(\posit_add.in2[1] ),
    .C(\posit_add.in2[3] ),
    .D(\posit_add.in2[2] ),
    .X(_2122_));
 sky130_fd_sc_hd__or4_4 _4142_ (.A(\posit_add.in2[7] ),
    .B(\posit_add.in2[5] ),
    .C(\posit_add.in2[4] ),
    .D(\posit_add.in2[6] ),
    .X(_2133_));
 sky130_fd_sc_hd__nor2_1 _4143_ (.A(net227),
    .B(_2133_),
    .Y(_2144_));
 sky130_fd_sc_hd__or3_1 _4144_ (.A(\posit_add.in2[9] ),
    .B(\posit_add.in2[8] ),
    .C(\posit_add.in2[10] ),
    .X(_2155_));
 sky130_fd_sc_hd__or4_4 _4145_ (.A(\posit_add.in2[11] ),
    .B(\posit_add.in2[9] ),
    .C(\posit_add.in2[8] ),
    .D(\posit_add.in2[10] ),
    .X(_2166_));
 sky130_fd_sc_hd__or2_1 _4146_ (.A(\posit_add.in2[13] ),
    .B(\posit_add.in2[12] ),
    .X(_2177_));
 sky130_fd_sc_hd__or4_4 _4147_ (.A(net227),
    .B(_2133_),
    .C(_2166_),
    .D(_2177_),
    .X(_2188_));
 sky130_fd_sc_hd__o41a_2 _4148_ (.A1(_2122_),
    .A2(_2133_),
    .A3(_2166_),
    .A4(_2177_),
    .B1(net229),
    .X(_2199_));
 sky130_fd_sc_hd__xnor2_2 _4149_ (.A(\posit_add.in2[14] ),
    .B(_2199_),
    .Y(_2210_));
 sky130_fd_sc_hd__inv_6 _4150_ (.A(net216),
    .Y(_2221_));
 sky130_fd_sc_hd__o31a_2 _4151_ (.A1(net227),
    .A2(_2133_),
    .A3(_2166_),
    .B1(net229),
    .X(_2232_));
 sky130_fd_sc_hd__xnor2_4 _4152_ (.A(\posit_add.in2[12] ),
    .B(_2232_),
    .Y(_2243_));
 sky130_fd_sc_hd__nor2_1 _4153_ (.A(net214),
    .B(_2243_),
    .Y(_2254_));
 sky130_fd_sc_hd__o21a_2 _4154_ (.A1(net227),
    .A2(_2133_),
    .B1(net230),
    .X(_2265_));
 sky130_fd_sc_hd__o31a_2 _4155_ (.A1(net227),
    .A2(_2133_),
    .A3(_2155_),
    .B1(net230),
    .X(_2276_));
 sky130_fd_sc_hd__xnor2_4 _4156_ (.A(\posit_add.in2[11] ),
    .B(_2276_),
    .Y(_2287_));
 sky130_fd_sc_hd__and2_1 _4157_ (.A(net214),
    .B(_2243_),
    .X(_2298_));
 sky130_fd_sc_hd__or3_4 _4158_ (.A(net214),
    .B(_2243_),
    .C(_2287_),
    .X(_2309_));
 sky130_fd_sc_hd__nand3_4 _4159_ (.A(net215),
    .B(_2243_),
    .C(_2287_),
    .Y(_2320_));
 sky130_fd_sc_hd__o41a_4 _4160_ (.A1(\posit_add.in2[12] ),
    .A2(_2122_),
    .A3(_2133_),
    .A4(_2166_),
    .B1(net229),
    .X(_2331_));
 sky130_fd_sc_hd__xnor2_4 _4161_ (.A(\posit_add.in2[13] ),
    .B(_2331_),
    .Y(_2342_));
 sky130_fd_sc_hd__xor2_4 _4162_ (.A(net214),
    .B(_2342_),
    .X(_2353_));
 sky130_fd_sc_hd__a21oi_4 _4163_ (.A1(_2309_),
    .A2(_2320_),
    .B1(_2353_),
    .Y(_2364_));
 sky130_fd_sc_hd__a21o_1 _4164_ (.A1(_2309_),
    .A2(_2320_),
    .B1(_2353_),
    .X(_2375_));
 sky130_fd_sc_hd__o41a_4 _4165_ (.A1(\posit_add.in2[9] ),
    .A2(\posit_add.in2[8] ),
    .A3(net227),
    .A4(_2133_),
    .B1(net230),
    .X(_2386_));
 sky130_fd_sc_hd__xnor2_4 _4166_ (.A(\posit_add.in2[10] ),
    .B(_2386_),
    .Y(_2397_));
 sky130_fd_sc_hd__nor2_1 _4167_ (.A(net214),
    .B(_2397_),
    .Y(_2408_));
 sky130_fd_sc_hd__o31a_4 _4168_ (.A1(\posit_add.in2[8] ),
    .A2(_2122_),
    .A3(_2133_),
    .B1(net230),
    .X(_2419_));
 sky130_fd_sc_hd__xnor2_2 _4169_ (.A(\posit_add.in2[9] ),
    .B(_2419_),
    .Y(_2430_));
 sky130_fd_sc_hd__xor2_4 _4170_ (.A(\posit_add.in2[9] ),
    .B(_2419_),
    .X(_2441_));
 sky130_fd_sc_hd__o21a_2 _4171_ (.A1(net214),
    .A2(_2397_),
    .B1(_2441_),
    .X(_2452_));
 sky130_fd_sc_hd__and2_1 _4172_ (.A(net216),
    .B(_2397_),
    .X(_2463_));
 sky130_fd_sc_hd__a21oi_4 _4173_ (.A1(net214),
    .A2(_2397_),
    .B1(_2441_),
    .Y(_2474_));
 sky130_fd_sc_hd__nor2_4 _4174_ (.A(_2452_),
    .B(_2474_),
    .Y(_2485_));
 sky130_fd_sc_hd__nand2_2 _4175_ (.A(net229),
    .B(net227),
    .Y(_2496_));
 sky130_fd_sc_hd__o31a_2 _4176_ (.A1(\posit_add.in2[5] ),
    .A2(\posit_add.in2[4] ),
    .A3(net227),
    .B1(net229),
    .X(_2507_));
 sky130_fd_sc_hd__o41a_4 _4177_ (.A1(\posit_add.in2[5] ),
    .A2(\posit_add.in2[4] ),
    .A3(\posit_add.in2[6] ),
    .A4(net227),
    .B1(net229),
    .X(_2518_));
 sky130_fd_sc_hd__xor2_4 _4178_ (.A(\posit_add.in2[7] ),
    .B(_2518_),
    .X(_2529_));
 sky130_fd_sc_hd__xnor2_4 _4179_ (.A(\posit_add.in2[8] ),
    .B(_2265_),
    .Y(_2540_));
 sky130_fd_sc_hd__clkinv_2 _4180_ (.A(_2540_),
    .Y(_2551_));
 sky130_fd_sc_hd__a21oi_1 _4181_ (.A1(net214),
    .A2(_2540_),
    .B1(_2529_),
    .Y(_2562_));
 sky130_fd_sc_hd__o21a_1 _4182_ (.A1(net214),
    .A2(_2540_),
    .B1(_2529_),
    .X(_2573_));
 sky130_fd_sc_hd__nor2_2 _4183_ (.A(_2562_),
    .B(_2573_),
    .Y(_2584_));
 sky130_fd_sc_hd__nand2_2 _4184_ (.A(_2485_),
    .B(_2584_),
    .Y(_2595_));
 sky130_fd_sc_hd__xor2_4 _4185_ (.A(\posit_add.in2[6] ),
    .B(_2507_),
    .X(_2606_));
 sky130_fd_sc_hd__inv_2 _4186_ (.A(_2606_),
    .Y(_2617_));
 sky130_fd_sc_hd__xnor2_4 _4187_ (.A(net215),
    .B(_2606_),
    .Y(_2628_));
 sky130_fd_sc_hd__o21ai_4 _4188_ (.A1(\posit_add.in2[4] ),
    .A2(net227),
    .B1(net229),
    .Y(_2639_));
 sky130_fd_sc_hd__xnor2_4 _4189_ (.A(\posit_add.in2[5] ),
    .B(_2639_),
    .Y(_2650_));
 sky130_fd_sc_hd__inv_2 _4190_ (.A(_2650_),
    .Y(_2661_));
 sky130_fd_sc_hd__xnor2_2 _4191_ (.A(net215),
    .B(_2650_),
    .Y(_2672_));
 sky130_fd_sc_hd__xor2_4 _4192_ (.A(net215),
    .B(_2650_),
    .X(_2683_));
 sky130_fd_sc_hd__nor2_2 _4193_ (.A(_2628_),
    .B(_2672_),
    .Y(_2694_));
 sky130_fd_sc_hd__xor2_4 _4194_ (.A(\posit_add.in2[4] ),
    .B(_2496_),
    .X(_2705_));
 sky130_fd_sc_hd__or2_2 _4195_ (.A(net215),
    .B(_2705_),
    .X(_2716_));
 sky130_fd_sc_hd__nand2_4 _4196_ (.A(net229),
    .B(_2111_),
    .Y(_2727_));
 sky130_fd_sc_hd__o21a_4 _4197_ (.A1(\posit_add.in2[2] ),
    .A2(_2111_),
    .B1(net229),
    .X(_2738_));
 sky130_fd_sc_hd__xnor2_4 _4198_ (.A(\posit_add.in2[3] ),
    .B(_2738_),
    .Y(_2749_));
 sky130_fd_sc_hd__xor2_4 _4199_ (.A(\posit_add.in2[3] ),
    .B(_2738_),
    .X(_2760_));
 sky130_fd_sc_hd__nand2_2 _4200_ (.A(net215),
    .B(_2705_),
    .Y(_2771_));
 sky130_fd_sc_hd__o21a_1 _4201_ (.A1(net215),
    .A2(_2705_),
    .B1(_2760_),
    .X(_2782_));
 sky130_fd_sc_hd__a2111o_4 _4202_ (.A1(_2749_),
    .A2(_2771_),
    .B1(_2782_),
    .C1(_2672_),
    .D1(_2628_),
    .X(_2793_));
 sky130_fd_sc_hd__xor2_4 _4203_ (.A(\posit_add.in2[2] ),
    .B(_2727_),
    .X(_2804_));
 sky130_fd_sc_hd__xnor2_2 _4204_ (.A(\posit_add.in2[2] ),
    .B(_2727_),
    .Y(_2815_));
 sky130_fd_sc_hd__nand2_2 _4205_ (.A(net215),
    .B(_2804_),
    .Y(_2826_));
 sky130_fd_sc_hd__o21ba_2 _4206_ (.A1(_2111_),
    .A2(_2826_),
    .B1_N(_2793_),
    .X(_2837_));
 sky130_fd_sc_hd__o21a_1 _4207_ (.A1(_2595_),
    .A2(_2837_),
    .B1(_2364_),
    .X(_2848_));
 sky130_fd_sc_hd__o21ai_4 _4208_ (.A1(_2595_),
    .A2(_2837_),
    .B1(_2364_),
    .Y(_2859_));
 sky130_fd_sc_hd__and3_4 _4209_ (.A(_2364_),
    .B(_2485_),
    .C(_2584_),
    .X(_2870_));
 sky130_fd_sc_hd__nand3_4 _4210_ (.A(_2364_),
    .B(_2485_),
    .C(_2584_),
    .Y(_2881_));
 sky130_fd_sc_hd__nand2_4 _4211_ (.A(\posit_add.in2[0] ),
    .B(net229),
    .Y(_2892_));
 sky130_fd_sc_hd__xnor2_2 _4212_ (.A(\posit_add.in2[1] ),
    .B(_2892_),
    .Y(_2903_));
 sky130_fd_sc_hd__xor2_4 _4213_ (.A(\posit_add.in2[1] ),
    .B(_2892_),
    .X(_2914_));
 sky130_fd_sc_hd__or2_2 _4214_ (.A(net215),
    .B(_2804_),
    .X(_2925_));
 sky130_fd_sc_hd__nor2_1 _4215_ (.A(_2914_),
    .B(_2925_),
    .Y(_2936_));
 sky130_fd_sc_hd__and4_1 _4216_ (.A(\posit_add.in2[0] ),
    .B(net214),
    .C(_2804_),
    .D(_2914_),
    .X(_2947_));
 sky130_fd_sc_hd__o31ai_4 _4217_ (.A1(_2793_),
    .A2(_2936_),
    .A3(_2947_),
    .B1(_2694_),
    .Y(_2958_));
 sky130_fd_sc_hd__a21oi_4 _4218_ (.A1(_2309_),
    .A2(_2320_),
    .B1(_2485_),
    .Y(_2969_));
 sky130_fd_sc_hd__a211oi_4 _4219_ (.A1(_2870_),
    .A2(_2958_),
    .B1(_2969_),
    .C1(_2353_),
    .Y(_2980_));
 sky130_fd_sc_hd__a211o_2 _4220_ (.A1(_2870_),
    .A2(_2958_),
    .B1(_2969_),
    .C1(_2353_),
    .X(_2990_));
 sky130_fd_sc_hd__nor2_2 _4221_ (.A(\posit_add.in2[0] ),
    .B(_2914_),
    .Y(_3001_));
 sky130_fd_sc_hd__o22a_1 _4222_ (.A1(_2826_),
    .A2(_2914_),
    .B1(_2925_),
    .B2(_3001_),
    .X(_3012_));
 sky130_fd_sc_hd__o22ai_4 _4223_ (.A1(_2826_),
    .A2(_2914_),
    .B1(_2925_),
    .B2(_3001_),
    .Y(_3023_));
 sky130_fd_sc_hd__a31oi_4 _4224_ (.A1(_2683_),
    .A2(_2716_),
    .A3(_2771_),
    .B1(_2628_),
    .Y(_3033_));
 sky130_fd_sc_hd__a31o_1 _4225_ (.A1(_2683_),
    .A2(_2716_),
    .A3(_2771_),
    .B1(_2628_),
    .X(_3044_));
 sky130_fd_sc_hd__mux2_8 _4226_ (.A0(_3012_),
    .A1(_3044_),
    .S(_2793_),
    .X(_3055_));
 sky130_fd_sc_hd__mux2_8 _4227_ (.A0(_3023_),
    .A1(_3033_),
    .S(_2793_),
    .X(_3065_));
 sky130_fd_sc_hd__xnor2_1 _4228_ (.A(net216),
    .B(_2540_),
    .Y(_3076_));
 sky130_fd_sc_hd__o32a_2 _4229_ (.A1(_2452_),
    .A2(_2474_),
    .A3(_3076_),
    .B1(_2463_),
    .B2(_2408_),
    .X(_3087_));
 sky130_fd_sc_hd__or3_4 _4230_ (.A(_2254_),
    .B(_2298_),
    .C(_2353_),
    .X(_3097_));
 sky130_fd_sc_hd__o21a_2 _4231_ (.A1(_2375_),
    .A2(_3087_),
    .B1(_3097_),
    .X(_3108_));
 sky130_fd_sc_hd__o21ai_4 _4232_ (.A1(_2375_),
    .A2(_3087_),
    .B1(_3097_),
    .Y(_3119_));
 sky130_fd_sc_hd__a21oi_4 _4233_ (.A1(_2870_),
    .A2(_3055_),
    .B1(_3119_),
    .Y(_3129_));
 sky130_fd_sc_hd__a21o_1 _4234_ (.A1(_2870_),
    .A2(_3055_),
    .B1(_3119_),
    .X(_3140_));
 sky130_fd_sc_hd__o211a_1 _4235_ (.A1(_2881_),
    .A2(_3065_),
    .B1(_3108_),
    .C1(_2606_),
    .X(_3151_));
 sky130_fd_sc_hd__o211a_1 _4236_ (.A1(_2881_),
    .A2(_3065_),
    .B1(_3108_),
    .C1(_2551_),
    .X(_3161_));
 sky130_fd_sc_hd__a211o_1 _4237_ (.A1(_2441_),
    .A2(net189),
    .B1(_3161_),
    .C1(net193),
    .X(_3172_));
 sky130_fd_sc_hd__a211o_1 _4238_ (.A1(_2529_),
    .A2(net189),
    .B1(_3151_),
    .C1(net191),
    .X(_3183_));
 sky130_fd_sc_hd__nand3_1 _4239_ (.A(net198),
    .B(_3172_),
    .C(_3183_),
    .Y(_3193_));
 sky130_fd_sc_hd__nor2_1 _4240_ (.A(_2144_),
    .B(_2881_),
    .Y(_3204_));
 sky130_fd_sc_hd__or2_1 _4241_ (.A(_2144_),
    .B(_2881_),
    .X(_3215_));
 sky130_fd_sc_hd__or2_1 _4242_ (.A(_2287_),
    .B(_3129_),
    .X(_3225_));
 sky130_fd_sc_hd__o21ai_1 _4243_ (.A1(_2397_),
    .A2(net188),
    .B1(_3225_),
    .Y(_3236_));
 sky130_fd_sc_hd__nor2_1 _4244_ (.A(net192),
    .B(_3236_),
    .Y(_3246_));
 sky130_fd_sc_hd__a211o_1 _4245_ (.A1(_2243_),
    .A2(net192),
    .B1(_3246_),
    .C1(net197),
    .X(_3257_));
 sky130_fd_sc_hd__a211o_1 _4246_ (.A1(_2870_),
    .A2(_3055_),
    .B1(_3119_),
    .C1(\posit_add.in2[0] ),
    .X(_3268_));
 sky130_fd_sc_hd__o21a_1 _4247_ (.A1(_2903_),
    .A2(net190),
    .B1(_3268_),
    .X(_3278_));
 sky130_fd_sc_hd__o2111a_2 _4248_ (.A1(_2903_),
    .A2(net190),
    .B1(_3268_),
    .C1(net191),
    .D1(net198),
    .X(_3289_));
 sky130_fd_sc_hd__o211a_1 _4249_ (.A1(_2881_),
    .A2(_3065_),
    .B1(_3108_),
    .C1(_2815_),
    .X(_3299_));
 sky130_fd_sc_hd__a211o_1 _4250_ (.A1(_2870_),
    .A2(_3055_),
    .B1(_3119_),
    .C1(_2815_),
    .X(_3310_));
 sky130_fd_sc_hd__a211oi_2 _4251_ (.A1(_2870_),
    .A2(_3055_),
    .B1(_3119_),
    .C1(_2705_),
    .Y(_3321_));
 sky130_fd_sc_hd__a211o_2 _4252_ (.A1(_2650_),
    .A2(net189),
    .B1(_3321_),
    .C1(net193),
    .X(_3331_));
 sky130_fd_sc_hd__a211o_4 _4253_ (.A1(_2760_),
    .A2(net189),
    .B1(_3299_),
    .C1(net191),
    .X(_3342_));
 sky130_fd_sc_hd__a31oi_4 _4254_ (.A1(net194),
    .A2(_3331_),
    .A3(_3342_),
    .B1(_3289_),
    .Y(_3352_));
 sky130_fd_sc_hd__a31o_4 _4255_ (.A1(net194),
    .A2(_3331_),
    .A3(_3342_),
    .B1(_3289_),
    .X(_3363_));
 sky130_fd_sc_hd__nor2_1 _4256_ (.A(net185),
    .B(_3363_),
    .Y(_3373_));
 sky130_fd_sc_hd__a31o_4 _4257_ (.A1(_3193_),
    .A2(net185),
    .A3(_3257_),
    .B1(_3373_),
    .X(_3384_));
 sky130_fd_sc_hd__or2_2 _4258_ (.A(_2100_),
    .B(_3384_),
    .X(_3394_));
 sky130_fd_sc_hd__nand2_1 _4259_ (.A(net192),
    .B(net188),
    .Y(_3403_));
 sky130_fd_sc_hd__and3_1 _4260_ (.A(\posit_add.in2[0] ),
    .B(net192),
    .C(net188),
    .X(_3410_));
 sky130_fd_sc_hd__o211a_1 _4261_ (.A1(_2881_),
    .A2(_3065_),
    .B1(_3108_),
    .C1(_2914_),
    .X(_3415_));
 sky130_fd_sc_hd__a211o_4 _4262_ (.A1(_2804_),
    .A2(net189),
    .B1(_3415_),
    .C1(net191),
    .X(_3416_));
 sky130_fd_sc_hd__a211o_1 _4263_ (.A1(_2870_),
    .A2(_3055_),
    .B1(_3119_),
    .C1(_2749_),
    .X(_3418_));
 sky130_fd_sc_hd__o211a_1 _4264_ (.A1(_2881_),
    .A2(_3065_),
    .B1(_3108_),
    .C1(_2749_),
    .X(_3419_));
 sky130_fd_sc_hd__a211o_4 _4265_ (.A1(_2705_),
    .A2(net189),
    .B1(_3419_),
    .C1(net193),
    .X(_3420_));
 sky130_fd_sc_hd__and2_2 _4266_ (.A(_3416_),
    .B(_3420_),
    .X(_3421_));
 sky130_fd_sc_hd__o31a_4 _4267_ (.A1(_0657_),
    .A2(net193),
    .A3(net190),
    .B1(net196),
    .X(_3422_));
 sky130_fd_sc_hd__a31o_1 _4268_ (.A1(net194),
    .A2(_3416_),
    .A3(_3420_),
    .B1(_3422_),
    .X(_3423_));
 sky130_fd_sc_hd__a21oi_4 _4269_ (.A1(net194),
    .A2(_3421_),
    .B1(_3422_),
    .Y(_3424_));
 sky130_fd_sc_hd__o211a_1 _4270_ (.A1(_2881_),
    .A2(_3065_),
    .B1(_3108_),
    .C1(_2650_),
    .X(_3425_));
 sky130_fd_sc_hd__o211a_1 _4271_ (.A1(_2881_),
    .A2(_3065_),
    .B1(_3108_),
    .C1(_2529_),
    .X(_3426_));
 sky130_fd_sc_hd__a21oi_1 _4272_ (.A1(_2551_),
    .A2(net188),
    .B1(_3426_),
    .Y(_3427_));
 sky130_fd_sc_hd__a211o_1 _4273_ (.A1(_2551_),
    .A2(net188),
    .B1(_3426_),
    .C1(_2980_),
    .X(_3428_));
 sky130_fd_sc_hd__a211o_1 _4274_ (.A1(_2606_),
    .A2(net188),
    .B1(_3425_),
    .C1(net191),
    .X(_3429_));
 sky130_fd_sc_hd__and3_1 _4275_ (.A(net184),
    .B(_3428_),
    .C(_3429_),
    .X(_3430_));
 sky130_fd_sc_hd__mux2_2 _4276_ (.A0(_2397_),
    .A1(_2430_),
    .S(net190),
    .X(_3431_));
 sky130_fd_sc_hd__a211o_1 _4277_ (.A1(_2287_),
    .A2(net192),
    .B1(net187),
    .C1(net197),
    .X(_3432_));
 sky130_fd_sc_hd__a21oi_2 _4278_ (.A1(_2980_),
    .A2(_3431_),
    .B1(_3432_),
    .Y(_3433_));
 sky130_fd_sc_hd__a221oi_4 _4279_ (.A1(net186),
    .A2(_3424_),
    .B1(_3430_),
    .B2(net197),
    .C1(_3433_),
    .Y(_3434_));
 sky130_fd_sc_hd__clkinv_4 _4280_ (.A(_3434_),
    .Y(_3435_));
 sky130_fd_sc_hd__a211o_1 _4281_ (.A1(_2529_),
    .A2(net189),
    .B1(_3151_),
    .C1(net193),
    .X(_3436_));
 sky130_fd_sc_hd__a211o_1 _4282_ (.A1(_2650_),
    .A2(net189),
    .B1(_3321_),
    .C1(net191),
    .X(_3437_));
 sky130_fd_sc_hd__a21o_1 _4283_ (.A1(_3436_),
    .A2(_3437_),
    .B1(net194),
    .X(_3438_));
 sky130_fd_sc_hd__a211o_1 _4284_ (.A1(_2441_),
    .A2(net188),
    .B1(_3161_),
    .C1(net191),
    .X(_3439_));
 sky130_fd_sc_hd__o21a_1 _4285_ (.A1(_2980_),
    .A2(_3236_),
    .B1(_3439_),
    .X(_3440_));
 sky130_fd_sc_hd__o21ai_1 _4286_ (.A1(net196),
    .A2(_3440_),
    .B1(_3438_),
    .Y(_3441_));
 sky130_fd_sc_hd__o211a_2 _4287_ (.A1(_2903_),
    .A2(net190),
    .B1(_3268_),
    .C1(net193),
    .X(_3442_));
 sky130_fd_sc_hd__o211a_2 _4288_ (.A1(_2760_),
    .A2(net190),
    .B1(_3310_),
    .C1(net191),
    .X(_3443_));
 sky130_fd_sc_hd__o21ai_4 _4289_ (.A1(_3442_),
    .A2(_3443_),
    .B1(net194),
    .Y(_3444_));
 sky130_fd_sc_hd__mux2_8 _4290_ (.A0(_3441_),
    .A1(_3444_),
    .S(net186),
    .X(_3445_));
 sky130_fd_sc_hd__inv_2 _4291_ (.A(_3445_),
    .Y(_3446_));
 sky130_fd_sc_hd__o211a_1 _4292_ (.A1(_1385_),
    .A2(_1869_),
    .B1(_1638_),
    .C1(_1352_),
    .X(_3447_));
 sky130_fd_sc_hd__o211a_1 _4293_ (.A1(_1385_),
    .A2(_1869_),
    .B1(_1561_),
    .C1(_1352_),
    .X(_3448_));
 sky130_fd_sc_hd__a211o_1 _4294_ (.A1(_1594_),
    .A2(net129),
    .B1(_3448_),
    .C1(net133),
    .X(_3449_));
 sky130_fd_sc_hd__a211o_1 _4295_ (.A1(_1671_),
    .A2(net129),
    .B1(_3447_),
    .C1(net131),
    .X(_3450_));
 sky130_fd_sc_hd__nand2_4 _4296_ (.A(_3449_),
    .B(_3450_),
    .Y(_3451_));
 sky130_fd_sc_hd__o211a_1 _4297_ (.A1(_1385_),
    .A2(_1869_),
    .B1(_1209_),
    .C1(_1352_),
    .X(_3452_));
 sky130_fd_sc_hd__o211a_1 _4298_ (.A1(_1385_),
    .A2(_1869_),
    .B1(_1121_),
    .C1(_1352_),
    .X(_3453_));
 sky130_fd_sc_hd__a211o_1 _4299_ (.A1(_1165_),
    .A2(net129),
    .B1(_3453_),
    .C1(net131),
    .X(_3454_));
 sky130_fd_sc_hd__a211o_1 _4300_ (.A1(_1242_),
    .A2(net129),
    .B1(_3452_),
    .C1(net133),
    .X(_3455_));
 sky130_fd_sc_hd__nand2_1 _4301_ (.A(_3454_),
    .B(_3455_),
    .Y(_3456_));
 sky130_fd_sc_hd__mux2_1 _4302_ (.A0(_3451_),
    .A1(_3456_),
    .S(net167),
    .X(_3457_));
 sky130_fd_sc_hd__nand3_2 _4303_ (.A(\posit_add.in1[0] ),
    .B(net133),
    .C(_1891_),
    .Y(_3458_));
 sky130_fd_sc_hd__a211o_1 _4304_ (.A1(_1374_),
    .A2(_1880_),
    .B1(_1484_),
    .C1(_1341_),
    .X(_3459_));
 sky130_fd_sc_hd__o211a_1 _4305_ (.A1(_1385_),
    .A2(_1869_),
    .B1(_1484_),
    .C1(_1352_),
    .X(_3460_));
 sky130_fd_sc_hd__o211ai_4 _4306_ (.A1(_1517_),
    .A2(_1891_),
    .B1(_3459_),
    .C1(net132),
    .Y(_3461_));
 sky130_fd_sc_hd__a21o_2 _4307_ (.A1(_3458_),
    .A2(_3461_),
    .B1(_1715_),
    .X(_3462_));
 sky130_fd_sc_hd__mux2_2 _4308_ (.A0(_3457_),
    .A1(_3462_),
    .S(net172),
    .X(_3463_));
 sky130_fd_sc_hd__inv_8 _4309_ (.A(net70),
    .Y(_3464_));
 sky130_fd_sc_hd__a211o_2 _4310_ (.A1(_2606_),
    .A2(net188),
    .B1(_3425_),
    .C1(net193),
    .X(_3465_));
 sky130_fd_sc_hd__o211ai_4 _4311_ (.A1(_2705_),
    .A2(net190),
    .B1(_3418_),
    .C1(net193),
    .Y(_3466_));
 sky130_fd_sc_hd__and3_2 _4312_ (.A(net196),
    .B(_3465_),
    .C(_3466_),
    .X(_3467_));
 sky130_fd_sc_hd__mux2_1 _4313_ (.A0(_3427_),
    .A1(_3431_),
    .S(_2990_),
    .X(_3468_));
 sky130_fd_sc_hd__o21ai_2 _4314_ (.A1(net196),
    .A2(_3468_),
    .B1(net185),
    .Y(_3469_));
 sky130_fd_sc_hd__or3_4 _4315_ (.A(_0657_),
    .B(net191),
    .C(net190),
    .X(_3470_));
 sky130_fd_sc_hd__a211o_2 _4316_ (.A1(_2804_),
    .A2(net188),
    .B1(_3415_),
    .C1(net193),
    .X(_3471_));
 sky130_fd_sc_hd__and2_1 _4317_ (.A(_3470_),
    .B(_3471_),
    .X(_3472_));
 sky130_fd_sc_hd__nor2_2 _4318_ (.A(net197),
    .B(_3472_),
    .Y(_3473_));
 sky130_fd_sc_hd__or2_2 _4319_ (.A(net197),
    .B(_3472_),
    .X(_3474_));
 sky130_fd_sc_hd__o22a_4 _4320_ (.A1(_3467_),
    .A2(_3469_),
    .B1(_3473_),
    .B2(net184),
    .X(_3475_));
 sky130_fd_sc_hd__a2bb2o_4 _4321_ (.A1_N(_3467_),
    .A2_N(_3469_),
    .B1(_3474_),
    .B2(net186),
    .X(_3476_));
 sky130_fd_sc_hd__and3_2 _4322_ (.A(net198),
    .B(_3331_),
    .C(_3342_),
    .X(_3477_));
 sky130_fd_sc_hd__a31o_2 _4323_ (.A1(net195),
    .A2(_3172_),
    .A3(_3183_),
    .B1(net187),
    .X(_3478_));
 sky130_fd_sc_hd__a31o_2 _4324_ (.A1(net194),
    .A2(net191),
    .A3(_3278_),
    .B1(net184),
    .X(_3479_));
 sky130_fd_sc_hd__o21ai_4 _4325_ (.A1(_3477_),
    .A2(_3478_),
    .B1(_3479_),
    .Y(_3480_));
 sky130_fd_sc_hd__o21a_4 _4326_ (.A1(_3477_),
    .A2(_3478_),
    .B1(_3479_),
    .X(_3481_));
 sky130_fd_sc_hd__a31o_1 _4327_ (.A1(net184),
    .A2(_3428_),
    .A3(_3429_),
    .B1(_3410_),
    .X(_3482_));
 sky130_fd_sc_hd__nand2_1 _4328_ (.A(net196),
    .B(net185),
    .Y(_3483_));
 sky130_fd_sc_hd__o2bb2a_1 _4329_ (.A1_N(net195),
    .A2_N(_3482_),
    .B1(_3483_),
    .B2(_3421_),
    .X(_3484_));
 sky130_fd_sc_hd__a2bb2o_1 _4330_ (.A1_N(_3421_),
    .A2_N(_3483_),
    .B1(_3482_),
    .B2(net195),
    .X(_3485_));
 sky130_fd_sc_hd__a21o_1 _4331_ (.A1(_3436_),
    .A2(_3437_),
    .B1(net198),
    .X(_3486_));
 sky130_fd_sc_hd__o31a_1 _4332_ (.A1(net194),
    .A2(_3442_),
    .A3(_3443_),
    .B1(net184),
    .X(_3487_));
 sky130_fd_sc_hd__and2_1 _4333_ (.A(_3486_),
    .B(_3487_),
    .X(_3488_));
 sky130_fd_sc_hd__nand2_1 _4334_ (.A(_3486_),
    .B(_3487_),
    .Y(_3489_));
 sky130_fd_sc_hd__a21oi_4 _4335_ (.A1(_3465_),
    .A2(_3466_),
    .B1(net196),
    .Y(_3490_));
 sky130_fd_sc_hd__a21o_1 _4336_ (.A1(_3465_),
    .A2(_3466_),
    .B1(net196),
    .X(_3491_));
 sky130_fd_sc_hd__a31oi_4 _4337_ (.A1(net196),
    .A2(_3470_),
    .A3(_3471_),
    .B1(net187),
    .Y(_3492_));
 sky130_fd_sc_hd__a31o_2 _4338_ (.A1(net196),
    .A2(_3470_),
    .A3(_3471_),
    .B1(net187),
    .X(_3493_));
 sky130_fd_sc_hd__nor2_1 _4339_ (.A(_3490_),
    .B(_3493_),
    .Y(_3494_));
 sky130_fd_sc_hd__nand2_1 _4340_ (.A(_3491_),
    .B(_3492_),
    .Y(_3495_));
 sky130_fd_sc_hd__a311oi_4 _4341_ (.A1(net194),
    .A2(_3416_),
    .A3(_3420_),
    .B1(_3422_),
    .C1(net186),
    .Y(_3496_));
 sky130_fd_sc_hd__a311o_4 _4342_ (.A1(net194),
    .A2(_3416_),
    .A3(_3420_),
    .B1(_3422_),
    .C1(net186),
    .X(_3497_));
 sky130_fd_sc_hd__nor2_8 _4343_ (.A(net186),
    .B(_3352_),
    .Y(_3498_));
 sky130_fd_sc_hd__nand2_4 _4344_ (.A(net184),
    .B(_3363_),
    .Y(_3499_));
 sky130_fd_sc_hd__nor2_1 _4345_ (.A(_3352_),
    .B(net178),
    .Y(_3500_));
 sky130_fd_sc_hd__nand2_4 _4346_ (.A(_3363_),
    .B(net180),
    .Y(_3501_));
 sky130_fd_sc_hd__a22o_4 _4347_ (.A1(_3491_),
    .A2(_3492_),
    .B1(net180),
    .B2(_3363_),
    .X(_3502_));
 sky130_fd_sc_hd__and2_1 _4348_ (.A(net151),
    .B(_3502_),
    .X(_3503_));
 sky130_fd_sc_hd__a21oi_4 _4349_ (.A1(net150),
    .A2(_3502_),
    .B1(net155),
    .Y(_3504_));
 sky130_fd_sc_hd__o21a_1 _4350_ (.A1(net164),
    .A2(_3504_),
    .B1(net125),
    .X(_3505_));
 sky130_fd_sc_hd__o21ai_4 _4351_ (.A1(net164),
    .A2(_3504_),
    .B1(net126),
    .Y(_3506_));
 sky130_fd_sc_hd__nor2_8 _4352_ (.A(\posit_add.in2[14] ),
    .B(_2188_),
    .Y(_3507_));
 sky130_fd_sc_hd__nor2_2 _4353_ (.A(net186),
    .B(_3444_),
    .Y(_3508_));
 sky130_fd_sc_hd__or2_4 _4354_ (.A(net186),
    .B(_3444_),
    .X(_3509_));
 sky130_fd_sc_hd__nor2_4 _4355_ (.A(net187),
    .B(_3474_),
    .Y(_3510_));
 sky130_fd_sc_hd__nand2_2 _4356_ (.A(net184),
    .B(_3473_),
    .Y(_3511_));
 sky130_fd_sc_hd__a21oi_4 _4357_ (.A1(net184),
    .A2(_3363_),
    .B1(net181),
    .Y(_3512_));
 sky130_fd_sc_hd__a21o_4 _4358_ (.A1(net184),
    .A2(_3363_),
    .B1(net180),
    .X(_3513_));
 sky130_fd_sc_hd__nand2_1 _4359_ (.A(net145),
    .B(_3513_),
    .Y(_3514_));
 sky130_fd_sc_hd__nand2_1 _4360_ (.A(net165),
    .B(net160),
    .Y(_3515_));
 sky130_fd_sc_hd__a31o_1 _4361_ (.A1(net151),
    .A2(net145),
    .A3(_3513_),
    .B1(net162),
    .X(_3516_));
 sky130_fd_sc_hd__o311a_1 _4362_ (.A1(net148),
    .A2(net141),
    .A3(_3512_),
    .B1(net158),
    .C1(net165),
    .X(_3517_));
 sky130_fd_sc_hd__a211o_1 _4363_ (.A1(net150),
    .A2(_3502_),
    .B1(net164),
    .C1(net155),
    .X(_3518_));
 sky130_fd_sc_hd__o2bb2a_4 _4364_ (.A1_N(_3486_),
    .A2_N(_3487_),
    .B1(_3490_),
    .B2(_3493_),
    .X(_3519_));
 sky130_fd_sc_hd__nor2_1 _4365_ (.A(net151),
    .B(_3502_),
    .Y(_3520_));
 sky130_fd_sc_hd__a211o_1 _4366_ (.A1(_3501_),
    .A2(_3519_),
    .B1(net162),
    .C1(net158),
    .X(_3521_));
 sky130_fd_sc_hd__a31o_1 _4367_ (.A1(net126),
    .A2(_3518_),
    .A3(_3521_),
    .B1(_3517_),
    .X(_3522_));
 sky130_fd_sc_hd__or4b_4 _4368_ (.A(_3506_),
    .B(net135),
    .C(net122),
    .D_N(net118),
    .X(_3523_));
 sky130_fd_sc_hd__nand2_1 _4369_ (.A(net141),
    .B(net177),
    .Y(_3524_));
 sky130_fd_sc_hd__nor2_1 _4370_ (.A(net145),
    .B(_3513_),
    .Y(_3525_));
 sky130_fd_sc_hd__a21o_1 _4371_ (.A1(net142),
    .A2(_3512_),
    .B1(net165),
    .X(_3526_));
 sky130_fd_sc_hd__a21o_1 _4372_ (.A1(net165),
    .A2(net142),
    .B1(net155),
    .X(_3527_));
 sky130_fd_sc_hd__nor2_1 _4373_ (.A(net155),
    .B(_3519_),
    .Y(_3528_));
 sky130_fd_sc_hd__a32o_1 _4374_ (.A1(net147),
    .A2(_3526_),
    .A3(_3527_),
    .B1(_3528_),
    .B2(_3516_),
    .X(_3529_));
 sky130_fd_sc_hd__nor2_4 _4375_ (.A(net156),
    .B(net150),
    .Y(_3530_));
 sky130_fd_sc_hd__or3_4 _4376_ (.A(_3352_),
    .B(_3490_),
    .C(_3493_),
    .X(_3531_));
 sky130_fd_sc_hd__and3_1 _4377_ (.A(net158),
    .B(net150),
    .C(_3531_),
    .X(_3532_));
 sky130_fd_sc_hd__o2111a_1 _4378_ (.A1(net145),
    .A2(_3513_),
    .B1(_3531_),
    .C1(net150),
    .D1(net158),
    .X(_3533_));
 sky130_fd_sc_hd__a221oi_4 _4379_ (.A1(_3501_),
    .A2(_3519_),
    .B1(_3531_),
    .B2(net151),
    .C1(net159),
    .Y(_3534_));
 sky130_fd_sc_hd__a2111o_1 _4380_ (.A1(_3514_),
    .A2(_3530_),
    .B1(_3533_),
    .C1(_3534_),
    .D1(net162),
    .X(_3535_));
 sky130_fd_sc_hd__a21o_1 _4381_ (.A1(net159),
    .A2(_3519_),
    .B1(net164),
    .X(_3536_));
 sky130_fd_sc_hd__o31a_1 _4382_ (.A1(_3503_),
    .A2(_3520_),
    .A3(_3536_),
    .B1(net125),
    .X(_3537_));
 sky130_fd_sc_hd__a22o_2 _4383_ (.A1(net128),
    .A2(_3529_),
    .B1(_3535_),
    .B2(_3537_),
    .X(_3538_));
 sky130_fd_sc_hd__inv_4 _4384_ (.A(net115),
    .Y(_3539_));
 sky130_fd_sc_hd__a22o_2 _4385_ (.A1(net120),
    .A2(net124),
    .B1(net118),
    .B2(net136),
    .X(_3540_));
 sky130_fd_sc_hd__nand4_4 _4386_ (.A(net140),
    .B(_3523_),
    .C(net116),
    .D(_3540_),
    .Y(_3541_));
 sky130_fd_sc_hd__nand2_4 _4387_ (.A(_3523_),
    .B(_3541_),
    .Y(_3542_));
 sky130_fd_sc_hd__nand2_4 _4388_ (.A(net145),
    .B(net115),
    .Y(_3543_));
 sky130_fd_sc_hd__nand2_2 _4389_ (.A(net180),
    .B(net118),
    .Y(_3544_));
 sky130_fd_sc_hd__or4b_4 _4390_ (.A(net177),
    .B(_3506_),
    .C(net135),
    .D_N(net118),
    .X(_3545_));
 sky130_fd_sc_hd__a22o_1 _4391_ (.A1(net121),
    .A2(net137),
    .B1(net118),
    .B2(net180),
    .X(_3546_));
 sky130_fd_sc_hd__nand2_4 _4392_ (.A(_3545_),
    .B(_3546_),
    .Y(_3547_));
 sky130_fd_sc_hd__xnor2_4 _4393_ (.A(_3543_),
    .B(_3547_),
    .Y(_3548_));
 sky130_fd_sc_hd__nand2b_2 _4394_ (.A_N(_3548_),
    .B(_3542_),
    .Y(_3549_));
 sky130_fd_sc_hd__xnor2_4 _4395_ (.A(_3542_),
    .B(_3548_),
    .Y(_3550_));
 sky130_fd_sc_hd__nor2_1 _4396_ (.A(net147),
    .B(_3531_),
    .Y(_3551_));
 sky130_fd_sc_hd__a21oi_4 _4397_ (.A1(_3502_),
    .A2(_3531_),
    .B1(net147),
    .Y(_3552_));
 sky130_fd_sc_hd__a221o_2 _4398_ (.A1(_3352_),
    .A2(_3423_),
    .B1(_3491_),
    .B2(_3492_),
    .C1(net186),
    .X(_3553_));
 sky130_fd_sc_hd__a21oi_1 _4399_ (.A1(_3501_),
    .A2(_3553_),
    .B1(net152),
    .Y(_3554_));
 sky130_fd_sc_hd__a21o_1 _4400_ (.A1(net146),
    .A2(_3513_),
    .B1(net159),
    .X(_3555_));
 sky130_fd_sc_hd__o32a_1 _4401_ (.A1(net156),
    .A2(_3552_),
    .A3(_3554_),
    .B1(_3555_),
    .B2(_3525_),
    .X(_3556_));
 sky130_fd_sc_hd__o21a_1 _4402_ (.A1(net142),
    .A2(_3512_),
    .B1(_3502_),
    .X(_3557_));
 sky130_fd_sc_hd__o211a_1 _4403_ (.A1(net142),
    .A2(_3512_),
    .B1(_3502_),
    .C1(net148),
    .X(_3558_));
 sky130_fd_sc_hd__o31ai_4 _4404_ (.A1(net160),
    .A2(_3552_),
    .A3(_3558_),
    .B1(net165),
    .Y(_3559_));
 sky130_fd_sc_hd__nand2_1 _4405_ (.A(net147),
    .B(net145),
    .Y(_3560_));
 sky130_fd_sc_hd__or3_1 _4406_ (.A(_3363_),
    .B(net152),
    .C(net142),
    .X(_3561_));
 sky130_fd_sc_hd__and2_4 _4407_ (.A(_3512_),
    .B(_3519_),
    .X(_3562_));
 sky130_fd_sc_hd__a21oi_1 _4408_ (.A1(_3512_),
    .A2(_3519_),
    .B1(net155),
    .Y(_3563_));
 sky130_fd_sc_hd__o211a_1 _4409_ (.A1(net148),
    .A2(_3557_),
    .B1(_3561_),
    .C1(_3563_),
    .X(_3564_));
 sky130_fd_sc_hd__o22a_1 _4410_ (.A1(net165),
    .A2(_3556_),
    .B1(_3559_),
    .B2(_3564_),
    .X(_3565_));
 sky130_fd_sc_hd__or2_4 _4411_ (.A(net125),
    .B(_3565_),
    .X(_3566_));
 sky130_fd_sc_hd__nand2_1 _4412_ (.A(_3501_),
    .B(_3513_),
    .Y(_3567_));
 sky130_fd_sc_hd__or2_2 _4413_ (.A(_3500_),
    .B(_3553_),
    .X(_3568_));
 sky130_fd_sc_hd__a21o_1 _4414_ (.A1(_3501_),
    .A2(_3513_),
    .B1(net141),
    .X(_3569_));
 sky130_fd_sc_hd__a21o_1 _4415_ (.A1(_3568_),
    .A2(_3569_),
    .B1(net153),
    .X(_3570_));
 sky130_fd_sc_hd__a211oi_1 _4416_ (.A1(_3568_),
    .A2(_3569_),
    .B1(net158),
    .C1(net153),
    .Y(_3571_));
 sky130_fd_sc_hd__mux2_2 _4417_ (.A0(_3424_),
    .A1(net178),
    .S(net141),
    .X(_3572_));
 sky130_fd_sc_hd__a21o_1 _4418_ (.A1(_3501_),
    .A2(_3513_),
    .B1(net158),
    .X(_3573_));
 sky130_fd_sc_hd__a21o_1 _4419_ (.A1(net141),
    .A2(net139),
    .B1(_3424_),
    .X(_3574_));
 sky130_fd_sc_hd__o2111a_1 _4420_ (.A1(net146),
    .A2(net140),
    .B1(_3423_),
    .C1(net158),
    .D1(net147),
    .X(_3575_));
 sky130_fd_sc_hd__a311o_1 _4421_ (.A1(net152),
    .A2(_3572_),
    .A3(_3573_),
    .B1(_3575_),
    .C1(net162),
    .X(_3576_));
 sky130_fd_sc_hd__a21oi_1 _4422_ (.A1(net141),
    .A2(net177),
    .B1(net139),
    .Y(_3577_));
 sky130_fd_sc_hd__o21a_1 _4423_ (.A1(_3525_),
    .A2(_3577_),
    .B1(_3530_),
    .X(_3578_));
 sky130_fd_sc_hd__nor2_1 _4424_ (.A(_3530_),
    .B(_3567_),
    .Y(_3579_));
 sky130_fd_sc_hd__o32a_1 _4425_ (.A1(net165),
    .A2(_3578_),
    .A3(_3579_),
    .B1(_3571_),
    .B2(_3576_),
    .X(_3580_));
 sky130_fd_sc_hd__mux2_2 _4426_ (.A0(_3565_),
    .A1(_3580_),
    .S(net125),
    .X(_3581_));
 sky130_fd_sc_hd__inv_2 _4427_ (.A(net95),
    .Y(_3582_));
 sky130_fd_sc_hd__nor2_2 _4428_ (.A(net159),
    .B(net96),
    .Y(_3583_));
 sky130_fd_sc_hd__and2b_1 _4429_ (.A_N(_3517_),
    .B(_3536_),
    .X(_3584_));
 sky130_fd_sc_hd__and3_1 _4430_ (.A(net155),
    .B(net151),
    .C(_3502_),
    .X(_3585_));
 sky130_fd_sc_hd__o31a_1 _4431_ (.A1(net164),
    .A2(_3504_),
    .A3(_3585_),
    .B1(net126),
    .X(_3586_));
 sky130_fd_sc_hd__a21oi_1 _4432_ (.A1(net142),
    .A2(_3512_),
    .B1(net148),
    .Y(_3587_));
 sky130_fd_sc_hd__o22a_1 _4433_ (.A1(_3521_),
    .A2(_3551_),
    .B1(_3587_),
    .B2(_3515_),
    .X(_3588_));
 sky130_fd_sc_hd__a2bb2o_4 _4434_ (.A1_N(net125),
    .A2_N(_3584_),
    .B1(_3586_),
    .B2(_3588_),
    .X(_3589_));
 sky130_fd_sc_hd__inv_6 _4435_ (.A(net114),
    .Y(_3590_));
 sky130_fd_sc_hd__nor2_8 _4436_ (.A(net148),
    .B(net114),
    .Y(_3591_));
 sky130_fd_sc_hd__a211o_1 _4437_ (.A1(net150),
    .A2(_3502_),
    .B1(_3519_),
    .C1(net155),
    .X(_3592_));
 sky130_fd_sc_hd__o311a_1 _4438_ (.A1(net158),
    .A2(_3562_),
    .A3(_3587_),
    .B1(_3592_),
    .C1(net162),
    .X(_3593_));
 sky130_fd_sc_hd__a31o_1 _4439_ (.A1(net159),
    .A2(_3514_),
    .A3(_3560_),
    .B1(_3534_),
    .X(_3594_));
 sky130_fd_sc_hd__a211o_2 _4440_ (.A1(net164),
    .A2(_3594_),
    .B1(_3593_),
    .C1(net125),
    .X(_3595_));
 sky130_fd_sc_hd__nand2_1 _4441_ (.A(net141),
    .B(_3500_),
    .Y(_3596_));
 sky130_fd_sc_hd__o221a_1 _4442_ (.A1(net155),
    .A2(net151),
    .B1(net177),
    .B2(_3531_),
    .C1(_3502_),
    .X(_3597_));
 sky130_fd_sc_hd__a21oi_1 _4443_ (.A1(_3530_),
    .A2(_3553_),
    .B1(_3597_),
    .Y(_3598_));
 sky130_fd_sc_hd__a32o_1 _4444_ (.A1(_3524_),
    .A2(_3530_),
    .A3(_3567_),
    .B1(_3568_),
    .B2(_3532_),
    .X(_3599_));
 sky130_fd_sc_hd__o22a_1 _4445_ (.A1(net165),
    .A2(_3598_),
    .B1(_3599_),
    .B2(_3559_),
    .X(_3600_));
 sky130_fd_sc_hd__o21a_2 _4446_ (.A1(net128),
    .A2(_3600_),
    .B1(_3595_),
    .X(_3601_));
 sky130_fd_sc_hd__o21ai_2 _4447_ (.A1(net128),
    .A2(_3600_),
    .B1(_3595_),
    .Y(_3602_));
 sky130_fd_sc_hd__nor2_1 _4448_ (.A(net139),
    .B(net114),
    .Y(_3603_));
 sky130_fd_sc_hd__or3b_2 _4449_ (.A(net148),
    .B(net94),
    .C_N(_3603_),
    .X(_3604_));
 sky130_fd_sc_hd__a21o_2 _4450_ (.A1(net150),
    .A2(net92),
    .B1(_3603_),
    .X(_3605_));
 sky130_fd_sc_hd__nand3_2 _4451_ (.A(_3583_),
    .B(_3604_),
    .C(_3605_),
    .Y(_3606_));
 sky130_fd_sc_hd__a21o_1 _4452_ (.A1(_3604_),
    .A2(_3605_),
    .B1(_3583_),
    .X(_3607_));
 sky130_fd_sc_hd__nand3_4 _4453_ (.A(_3550_),
    .B(_3606_),
    .C(_3607_),
    .Y(_3608_));
 sky130_fd_sc_hd__o21ai_4 _4454_ (.A1(_3543_),
    .A2(_3547_),
    .B1(_3545_),
    .Y(_3609_));
 sky130_fd_sc_hd__nand2_2 _4455_ (.A(net150),
    .B(net115),
    .Y(_3610_));
 sky130_fd_sc_hd__nand2_8 _4456_ (.A(net140),
    .B(net121),
    .Y(_3611_));
 sky130_fd_sc_hd__nor2_1 _4457_ (.A(_3544_),
    .B(_3611_),
    .Y(_3612_));
 sky130_fd_sc_hd__a22o_2 _4458_ (.A1(net180),
    .A2(net121),
    .B1(net118),
    .B2(net140),
    .X(_3613_));
 sky130_fd_sc_hd__o21ai_4 _4459_ (.A1(_3544_),
    .A2(_3611_),
    .B1(_3613_),
    .Y(_3614_));
 sky130_fd_sc_hd__xor2_4 _4460_ (.A(_3610_),
    .B(_3614_),
    .X(_3615_));
 sky130_fd_sc_hd__xor2_4 _4461_ (.A(_3609_),
    .B(_3615_),
    .X(_3616_));
 sky130_fd_sc_hd__nor2_2 _4462_ (.A(net164),
    .B(net96),
    .Y(_3617_));
 sky130_fd_sc_hd__or4_4 _4463_ (.A(net159),
    .B(net143),
    .C(net114),
    .D(net94),
    .X(_3618_));
 sky130_fd_sc_hd__a22o_2 _4464_ (.A1(net145),
    .A2(_3590_),
    .B1(net92),
    .B2(net155),
    .X(_3619_));
 sky130_fd_sc_hd__nand3_4 _4465_ (.A(_3617_),
    .B(_3618_),
    .C(_3619_),
    .Y(_3620_));
 sky130_fd_sc_hd__a21o_1 _4466_ (.A1(_3618_),
    .A2(_3619_),
    .B1(_3617_),
    .X(_3621_));
 sky130_fd_sc_hd__and3_2 _4467_ (.A(_3616_),
    .B(_3620_),
    .C(_3621_),
    .X(_3622_));
 sky130_fd_sc_hd__a21oi_4 _4468_ (.A1(_3620_),
    .A2(_3621_),
    .B1(_3616_),
    .Y(_3623_));
 sky130_fd_sc_hd__a211oi_4 _4469_ (.A1(_3549_),
    .A2(_3608_),
    .B1(_3622_),
    .C1(_3623_),
    .Y(_3624_));
 sky130_fd_sc_hd__o211a_2 _4470_ (.A1(_3622_),
    .A2(_3623_),
    .B1(_3549_),
    .C1(_3608_),
    .X(_3625_));
 sky130_fd_sc_hd__a21boi_4 _4471_ (.A1(_3583_),
    .A2(_3605_),
    .B1_N(_3604_),
    .Y(_3626_));
 sky130_fd_sc_hd__nor2_1 _4472_ (.A(net152),
    .B(_3572_),
    .Y(_3627_));
 sky130_fd_sc_hd__a21o_1 _4473_ (.A1(net152),
    .A2(_3574_),
    .B1(net157),
    .X(_3628_));
 sky130_fd_sc_hd__o221a_1 _4474_ (.A1(net158),
    .A2(net180),
    .B1(_3627_),
    .B2(_3628_),
    .C1(net126),
    .X(_3629_));
 sky130_fd_sc_hd__a21o_1 _4475_ (.A1(_3423_),
    .A2(net140),
    .B1(net141),
    .X(_3630_));
 sky130_fd_sc_hd__a22o_1 _4476_ (.A1(_3363_),
    .A2(net141),
    .B1(net178),
    .B2(_3630_),
    .X(_3631_));
 sky130_fd_sc_hd__a221o_1 _4477_ (.A1(net156),
    .A2(_3567_),
    .B1(_3596_),
    .B2(_3533_),
    .C1(net125),
    .X(_3632_));
 sky130_fd_sc_hd__a21oi_1 _4478_ (.A1(_3530_),
    .A2(_3631_),
    .B1(_3632_),
    .Y(_3633_));
 sky130_fd_sc_hd__o21a_4 _4479_ (.A1(_3629_),
    .A2(_3633_),
    .B1(net162),
    .X(_3634_));
 sky130_fd_sc_hd__a21o_1 _4480_ (.A1(_3568_),
    .A2(_3630_),
    .B1(net147),
    .X(_3635_));
 sky130_fd_sc_hd__a211o_1 _4481_ (.A1(_3424_),
    .A2(net146),
    .B1(net139),
    .C1(net152),
    .X(_3636_));
 sky130_fd_sc_hd__a21oi_1 _4482_ (.A1(_3501_),
    .A2(_3553_),
    .B1(net147),
    .Y(_3637_));
 sky130_fd_sc_hd__or3_1 _4483_ (.A(_3424_),
    .B(net146),
    .C(net139),
    .X(_3638_));
 sky130_fd_sc_hd__a21o_1 _4484_ (.A1(_3630_),
    .A2(_3638_),
    .B1(net147),
    .X(_3639_));
 sky130_fd_sc_hd__a211oi_1 _4485_ (.A1(_3363_),
    .A2(net141),
    .B1(_3572_),
    .C1(net152),
    .Y(_3640_));
 sky130_fd_sc_hd__o21a_1 _4486_ (.A1(_3562_),
    .A2(_3637_),
    .B1(net159),
    .X(_3641_));
 sky130_fd_sc_hd__a311o_4 _4487_ (.A1(net156),
    .A2(_3635_),
    .A3(_3636_),
    .B1(_3641_),
    .C1(net128),
    .X(_3642_));
 sky130_fd_sc_hd__and3_1 _4488_ (.A(net156),
    .B(_3570_),
    .C(_3639_),
    .X(_3643_));
 sky130_fd_sc_hd__a31o_1 _4489_ (.A1(net152),
    .A2(_3569_),
    .A3(_3638_),
    .B1(_3640_),
    .X(_3644_));
 sky130_fd_sc_hd__a211o_2 _4490_ (.A1(net158),
    .A2(_3644_),
    .B1(_3643_),
    .C1(net125),
    .X(_3645_));
 sky130_fd_sc_hd__a31oi_4 _4491_ (.A1(net165),
    .A2(_3642_),
    .A3(_3645_),
    .B1(_3634_),
    .Y(_3646_));
 sky130_fd_sc_hd__a31o_4 _4492_ (.A1(net165),
    .A2(_3642_),
    .A3(_3645_),
    .B1(_3634_),
    .X(_3647_));
 sky130_fd_sc_hd__nor2_2 _4493_ (.A(net125),
    .B(net68),
    .Y(_3648_));
 sky130_fd_sc_hd__or3_1 _4494_ (.A(net125),
    .B(_3626_),
    .C(_3646_),
    .X(_3649_));
 sky130_fd_sc_hd__xor2_4 _4495_ (.A(_3626_),
    .B(_3648_),
    .X(_3650_));
 sky130_fd_sc_hd__xnor2_4 _4496_ (.A(net135),
    .B(_3650_),
    .Y(_3651_));
 sky130_fd_sc_hd__or3_4 _4497_ (.A(_3624_),
    .B(_3625_),
    .C(_3651_),
    .X(_3652_));
 sky130_fd_sc_hd__and2b_2 _4498_ (.A_N(_3624_),
    .B(_3652_),
    .X(_3653_));
 sky130_fd_sc_hd__a21o_2 _4499_ (.A1(_3609_),
    .A2(_3615_),
    .B1(_3622_),
    .X(_3654_));
 sky130_fd_sc_hd__a31o_4 _4500_ (.A1(net150),
    .A2(net116),
    .A3(_3613_),
    .B1(_3612_),
    .X(_3655_));
 sky130_fd_sc_hd__nand2_4 _4501_ (.A(net156),
    .B(net116),
    .Y(_3656_));
 sky130_fd_sc_hd__nand2_4 _4502_ (.A(net145),
    .B(net118),
    .Y(_3657_));
 sky130_fd_sc_hd__xor2_4 _4503_ (.A(_3611_),
    .B(_3657_),
    .X(_3658_));
 sky130_fd_sc_hd__nand2b_1 _4504_ (.A_N(_3656_),
    .B(_3658_),
    .Y(_3659_));
 sky130_fd_sc_hd__xnor2_4 _4505_ (.A(_3656_),
    .B(_3658_),
    .Y(_3660_));
 sky130_fd_sc_hd__xnor2_4 _4506_ (.A(_3655_),
    .B(_3660_),
    .Y(_3661_));
 sky130_fd_sc_hd__nor2_4 _4507_ (.A(net164),
    .B(net94),
    .Y(_3662_));
 sky130_fd_sc_hd__xnor2_4 _4508_ (.A(_3591_),
    .B(_3662_),
    .Y(_3663_));
 sky130_fd_sc_hd__xnor2_4 _4509_ (.A(_3566_),
    .B(_3663_),
    .Y(_3664_));
 sky130_fd_sc_hd__nor2_1 _4510_ (.A(_3661_),
    .B(_3664_),
    .Y(_3665_));
 sky130_fd_sc_hd__xor2_4 _4511_ (.A(_3661_),
    .B(_3664_),
    .X(_3666_));
 sky130_fd_sc_hd__nand2_1 _4512_ (.A(_3654_),
    .B(_3666_),
    .Y(_3667_));
 sky130_fd_sc_hd__xnor2_4 _4513_ (.A(_3654_),
    .B(_3666_),
    .Y(_3668_));
 sky130_fd_sc_hd__or2_4 _4514_ (.A(net211),
    .B(_3646_),
    .X(_3669_));
 sky130_fd_sc_hd__a21o_2 _4515_ (.A1(_3618_),
    .A2(_3620_),
    .B1(_3669_),
    .X(_3670_));
 sky130_fd_sc_hd__nand3_2 _4516_ (.A(_3618_),
    .B(_3620_),
    .C(_3669_),
    .Y(_3671_));
 sky130_fd_sc_hd__nand2_4 _4517_ (.A(_3670_),
    .B(_3671_),
    .Y(_3672_));
 sky130_fd_sc_hd__xnor2_4 _4518_ (.A(net177),
    .B(_3672_),
    .Y(_3673_));
 sky130_fd_sc_hd__xnor2_4 _4519_ (.A(_3668_),
    .B(_3673_),
    .Y(_3674_));
 sky130_fd_sc_hd__o21ai_2 _4520_ (.A1(net135),
    .A2(_3650_),
    .B1(_3649_),
    .Y(_3675_));
 sky130_fd_sc_hd__xnor2_2 _4521_ (.A(_3653_),
    .B(_3674_),
    .Y(_3676_));
 sky130_fd_sc_hd__nand2b_1 _4522_ (.A_N(_3676_),
    .B(_3675_),
    .Y(_3677_));
 sky130_fd_sc_hd__o21a_2 _4523_ (.A1(_3653_),
    .A2(_3674_),
    .B1(_3677_),
    .X(_3678_));
 sky130_fd_sc_hd__o21a_2 _4524_ (.A1(_3611_),
    .A2(_3657_),
    .B1(_3659_),
    .X(_3679_));
 sky130_fd_sc_hd__nand2_2 _4525_ (.A(net162),
    .B(net116),
    .Y(_3680_));
 sky130_fd_sc_hd__a22o_1 _4526_ (.A1(net145),
    .A2(net121),
    .B1(net119),
    .B2(net150),
    .X(_3681_));
 sky130_fd_sc_hd__or4b_1 _4527_ (.A(net148),
    .B(net143),
    .C(_3506_),
    .D_N(net119),
    .X(_3682_));
 sky130_fd_sc_hd__nand2_2 _4528_ (.A(_3681_),
    .B(_3682_),
    .Y(_3683_));
 sky130_fd_sc_hd__xnor2_4 _4529_ (.A(_3680_),
    .B(_3683_),
    .Y(_3684_));
 sky130_fd_sc_hd__xnor2_4 _4530_ (.A(_3679_),
    .B(_3684_),
    .Y(_3685_));
 sky130_fd_sc_hd__or2_4 _4531_ (.A(net210),
    .B(net96),
    .X(_3686_));
 sky130_fd_sc_hd__o21a_1 _4532_ (.A1(net159),
    .A2(net114),
    .B1(_3595_),
    .X(_3687_));
 sky130_fd_sc_hd__a41o_2 _4533_ (.A1(net128),
    .A2(net164),
    .A3(net155),
    .A4(net92),
    .B1(_3687_),
    .X(_3688_));
 sky130_fd_sc_hd__xnor2_4 _4534_ (.A(_3686_),
    .B(_3688_),
    .Y(_3689_));
 sky130_fd_sc_hd__o2bb2ai_4 _4535_ (.A1_N(_3591_),
    .A2_N(_3662_),
    .B1(_3663_),
    .B2(_3566_),
    .Y(_3690_));
 sky130_fd_sc_hd__xnor2_4 _4536_ (.A(_3689_),
    .B(_3690_),
    .Y(_3691_));
 sky130_fd_sc_hd__xnor2_4 _4537_ (.A(_3685_),
    .B(_3691_),
    .Y(_3692_));
 sky130_fd_sc_hd__a21oi_4 _4538_ (.A1(_3655_),
    .A2(_3660_),
    .B1(_3665_),
    .Y(_3693_));
 sky130_fd_sc_hd__xnor2_4 _4539_ (.A(net139),
    .B(_3693_),
    .Y(_3694_));
 sky130_fd_sc_hd__xnor2_4 _4540_ (.A(_3692_),
    .B(_3694_),
    .Y(_3695_));
 sky130_fd_sc_hd__o21ai_4 _4541_ (.A1(net178),
    .A2(_3672_),
    .B1(_3670_),
    .Y(_3696_));
 sky130_fd_sc_hd__o21a_2 _4542_ (.A1(_3668_),
    .A2(_3673_),
    .B1(_3667_),
    .X(_3697_));
 sky130_fd_sc_hd__xnor2_4 _4543_ (.A(_3696_),
    .B(_3697_),
    .Y(_3698_));
 sky130_fd_sc_hd__xnor2_4 _4544_ (.A(_3695_),
    .B(_3698_),
    .Y(_3699_));
 sky130_fd_sc_hd__xnor2_4 _4545_ (.A(_3678_),
    .B(_3699_),
    .Y(_3700_));
 sky130_fd_sc_hd__xnor2_1 _4546_ (.A(_3675_),
    .B(_3676_),
    .Y(_3701_));
 sky130_fd_sc_hd__and4_4 _4547_ (.A(net195),
    .B(net192),
    .C(net184),
    .D(_3278_),
    .X(_3702_));
 sky130_fd_sc_hd__or4b_2 _4548_ (.A(net196),
    .B(net193),
    .C(net186),
    .D_N(_3278_),
    .X(_3703_));
 sky130_fd_sc_hd__or4b_4 _4549_ (.A(_3506_),
    .B(net123),
    .C(net174),
    .D_N(net118),
    .X(_3704_));
 sky130_fd_sc_hd__a22o_2 _4550_ (.A1(net124),
    .A2(net118),
    .B1(_3702_),
    .B2(net121),
    .X(_3705_));
 sky130_fd_sc_hd__nand4_4 _4551_ (.A(net180),
    .B(net116),
    .C(_3704_),
    .D(_3705_),
    .Y(_3706_));
 sky130_fd_sc_hd__nand2_4 _4552_ (.A(_3704_),
    .B(_3706_),
    .Y(_3707_));
 sky130_fd_sc_hd__a22o_1 _4553_ (.A1(net140),
    .A2(net116),
    .B1(_3540_),
    .B2(_3523_),
    .X(_3708_));
 sky130_fd_sc_hd__nand2_2 _4554_ (.A(_3541_),
    .B(_3708_),
    .Y(_3709_));
 sky130_fd_sc_hd__and3_1 _4555_ (.A(_3541_),
    .B(_3707_),
    .C(_3708_),
    .X(_3710_));
 sky130_fd_sc_hd__xnor2_4 _4556_ (.A(_3707_),
    .B(_3709_),
    .Y(_3711_));
 sky130_fd_sc_hd__nor2_2 _4557_ (.A(net148),
    .B(net96),
    .Y(_3712_));
 sky130_fd_sc_hd__or2_2 _4558_ (.A(net177),
    .B(net114),
    .X(_3713_));
 sky130_fd_sc_hd__or3_2 _4559_ (.A(net143),
    .B(net94),
    .C(_3713_),
    .X(_3714_));
 sky130_fd_sc_hd__o21ai_4 _4560_ (.A1(net143),
    .A2(net94),
    .B1(_3713_),
    .Y(_3715_));
 sky130_fd_sc_hd__nand3_2 _4561_ (.A(_3712_),
    .B(_3714_),
    .C(_3715_),
    .Y(_3716_));
 sky130_fd_sc_hd__a21o_1 _4562_ (.A1(_3714_),
    .A2(_3715_),
    .B1(_3712_),
    .X(_3717_));
 sky130_fd_sc_hd__nand3_2 _4563_ (.A(_3711_),
    .B(_3716_),
    .C(_3717_),
    .Y(_3718_));
 sky130_fd_sc_hd__a31o_2 _4564_ (.A1(_3711_),
    .A2(_3716_),
    .A3(_3717_),
    .B1(_3710_),
    .X(_3719_));
 sky130_fd_sc_hd__a21o_2 _4565_ (.A1(_3606_),
    .A2(_3607_),
    .B1(_3550_),
    .X(_3720_));
 sky130_fd_sc_hd__and3_4 _4566_ (.A(_3608_),
    .B(_3719_),
    .C(_3720_),
    .X(_3721_));
 sky130_fd_sc_hd__a21oi_4 _4567_ (.A1(_3608_),
    .A2(_3720_),
    .B1(_3719_),
    .Y(_3722_));
 sky130_fd_sc_hd__a21boi_4 _4568_ (.A1(_3712_),
    .A2(_3715_),
    .B1_N(_3714_),
    .Y(_3723_));
 sky130_fd_sc_hd__and2b_2 _4569_ (.A_N(_3723_),
    .B(_3634_),
    .X(_3724_));
 sky130_fd_sc_hd__xor2_4 _4570_ (.A(_3634_),
    .B(_3723_),
    .X(_3725_));
 sky130_fd_sc_hd__nor2_2 _4571_ (.A(net122),
    .B(_3725_),
    .Y(_3726_));
 sky130_fd_sc_hd__xnor2_4 _4572_ (.A(net122),
    .B(_3725_),
    .Y(_3727_));
 sky130_fd_sc_hd__nor3_2 _4573_ (.A(_3721_),
    .B(_3722_),
    .C(_3727_),
    .Y(_3728_));
 sky130_fd_sc_hd__or3_4 _4574_ (.A(_3721_),
    .B(_3722_),
    .C(_3727_),
    .X(_3729_));
 sky130_fd_sc_hd__o21ai_4 _4575_ (.A1(_3624_),
    .A2(_3625_),
    .B1(_3651_),
    .Y(_3730_));
 sky130_fd_sc_hd__o211ai_4 _4576_ (.A1(_3721_),
    .A2(_3728_),
    .B1(_3730_),
    .C1(_3652_),
    .Y(_3731_));
 sky130_fd_sc_hd__inv_2 _4577_ (.A(_3731_),
    .Y(_3732_));
 sky130_fd_sc_hd__a211o_2 _4578_ (.A1(_3652_),
    .A2(_3730_),
    .B1(_3728_),
    .C1(_3721_),
    .X(_3733_));
 sky130_fd_sc_hd__o211a_2 _4579_ (.A1(_3724_),
    .A2(_3726_),
    .B1(_3731_),
    .C1(_3733_),
    .X(_3734_));
 sky130_fd_sc_hd__o21a_1 _4580_ (.A1(_3732_),
    .A2(_3734_),
    .B1(_3701_),
    .X(_3735_));
 sky130_fd_sc_hd__or3_1 _4581_ (.A(_3701_),
    .B(_3732_),
    .C(_3734_),
    .X(_3736_));
 sky130_fd_sc_hd__a211oi_4 _4582_ (.A1(_3731_),
    .A2(_3733_),
    .B1(_3724_),
    .C1(_3726_),
    .Y(_3737_));
 sky130_fd_sc_hd__nor2_4 _4583_ (.A(_3734_),
    .B(_3737_),
    .Y(_3738_));
 sky130_fd_sc_hd__nand2_1 _4584_ (.A(net115),
    .B(_3702_),
    .Y(_3739_));
 sky130_fd_sc_hd__and4_4 _4585_ (.A(net136),
    .B(net118),
    .C(net115),
    .D(_3702_),
    .X(_3740_));
 sky130_fd_sc_hd__a22o_1 _4586_ (.A1(net180),
    .A2(net116),
    .B1(_3704_),
    .B2(_3705_),
    .X(_3741_));
 sky130_fd_sc_hd__and2_2 _4587_ (.A(_3706_),
    .B(_3741_),
    .X(_3742_));
 sky130_fd_sc_hd__and2_1 _4588_ (.A(_3740_),
    .B(_3742_),
    .X(_3743_));
 sky130_fd_sc_hd__xor2_4 _4589_ (.A(_3740_),
    .B(_3742_),
    .X(_3744_));
 sky130_fd_sc_hd__nor2_2 _4590_ (.A(net143),
    .B(net96),
    .Y(_3745_));
 sky130_fd_sc_hd__or2_2 _4591_ (.A(net135),
    .B(net114),
    .X(_3746_));
 sky130_fd_sc_hd__o21ai_4 _4592_ (.A1(net139),
    .A2(net93),
    .B1(_3746_),
    .Y(_3747_));
 sky130_fd_sc_hd__or3_2 _4593_ (.A(net139),
    .B(net93),
    .C(_3746_),
    .X(_3748_));
 sky130_fd_sc_hd__nand3_2 _4594_ (.A(_3745_),
    .B(_3747_),
    .C(_3748_),
    .Y(_3749_));
 sky130_fd_sc_hd__a21o_1 _4595_ (.A1(_3747_),
    .A2(_3748_),
    .B1(_3745_),
    .X(_3750_));
 sky130_fd_sc_hd__nand3_2 _4596_ (.A(_3744_),
    .B(_3749_),
    .C(_3750_),
    .Y(_3751_));
 sky130_fd_sc_hd__a31o_2 _4597_ (.A1(_3744_),
    .A2(_3749_),
    .A3(_3750_),
    .B1(_3743_),
    .X(_3752_));
 sky130_fd_sc_hd__a21o_2 _4598_ (.A1(_3716_),
    .A2(_3717_),
    .B1(_3711_),
    .X(_3753_));
 sky130_fd_sc_hd__and3_4 _4599_ (.A(_3718_),
    .B(_3752_),
    .C(_3753_),
    .X(_3754_));
 sky130_fd_sc_hd__a21oi_4 _4600_ (.A1(_3718_),
    .A2(_3753_),
    .B1(_3752_),
    .Y(_3755_));
 sky130_fd_sc_hd__a21bo_4 _4601_ (.A1(_3745_),
    .A2(_3747_),
    .B1_N(_3748_),
    .X(_3756_));
 sky130_fd_sc_hd__nor2_4 _4602_ (.A(net159),
    .B(net68),
    .Y(_3757_));
 sky130_fd_sc_hd__nand2_1 _4603_ (.A(_3756_),
    .B(_3757_),
    .Y(_3758_));
 sky130_fd_sc_hd__xnor2_4 _4604_ (.A(_3756_),
    .B(_3757_),
    .Y(_3759_));
 sky130_fd_sc_hd__xnor2_4 _4605_ (.A(net174),
    .B(_3759_),
    .Y(_3760_));
 sky130_fd_sc_hd__nor3_4 _4606_ (.A(_3754_),
    .B(_3755_),
    .C(_3760_),
    .Y(_3761_));
 sky130_fd_sc_hd__o21ai_4 _4607_ (.A1(_3721_),
    .A2(_3722_),
    .B1(_3727_),
    .Y(_3762_));
 sky130_fd_sc_hd__o211ai_4 _4608_ (.A1(_3754_),
    .A2(_3761_),
    .B1(_3762_),
    .C1(_3729_),
    .Y(_3763_));
 sky130_fd_sc_hd__o21ai_4 _4609_ (.A1(net174),
    .A2(_3759_),
    .B1(_3758_),
    .Y(_3764_));
 sky130_fd_sc_hd__a211o_4 _4610_ (.A1(_3729_),
    .A2(_3762_),
    .B1(_3761_),
    .C1(_3754_),
    .X(_3765_));
 sky130_fd_sc_hd__and3_2 _4611_ (.A(_3763_),
    .B(_3764_),
    .C(_3765_),
    .X(_3766_));
 sky130_fd_sc_hd__a21boi_4 _4612_ (.A1(_3764_),
    .A2(_3765_),
    .B1_N(_3763_),
    .Y(_3767_));
 sky130_fd_sc_hd__and2b_2 _4613_ (.A_N(_3767_),
    .B(_3738_),
    .X(_3768_));
 sky130_fd_sc_hd__xnor2_4 _4614_ (.A(_3738_),
    .B(_3767_),
    .Y(_3769_));
 sky130_fd_sc_hd__nor2_1 _4615_ (.A(net93),
    .B(net174),
    .Y(_3770_));
 sky130_fd_sc_hd__or3_4 _4616_ (.A(net93),
    .B(net174),
    .C(_3746_),
    .X(_3771_));
 sky130_fd_sc_hd__nor2_2 _4617_ (.A(net177),
    .B(net95),
    .Y(_3772_));
 sky130_fd_sc_hd__a22o_2 _4618_ (.A1(net136),
    .A2(net92),
    .B1(_3702_),
    .B2(_3590_),
    .X(_3773_));
 sky130_fd_sc_hd__nand3_4 _4619_ (.A(_3771_),
    .B(_3772_),
    .C(_3773_),
    .Y(_3774_));
 sky130_fd_sc_hd__nand2_4 _4620_ (.A(_3771_),
    .B(_3774_),
    .Y(_3775_));
 sky130_fd_sc_hd__nor2_4 _4621_ (.A(net143),
    .B(_3646_),
    .Y(_3776_));
 sky130_fd_sc_hd__and2_1 _4622_ (.A(_3775_),
    .B(_3776_),
    .X(_3777_));
 sky130_fd_sc_hd__nor2_1 _4623_ (.A(net122),
    .B(_3539_),
    .Y(_3778_));
 sky130_fd_sc_hd__a21o_1 _4624_ (.A1(_3771_),
    .A2(_3773_),
    .B1(_3772_),
    .X(_3779_));
 sky130_fd_sc_hd__and3_2 _4625_ (.A(_3774_),
    .B(_3778_),
    .C(_3779_),
    .X(_3780_));
 sky130_fd_sc_hd__o2bb2a_1 _4626_ (.A1_N(net119),
    .A2_N(_3702_),
    .B1(_3539_),
    .B2(net135),
    .X(_3781_));
 sky130_fd_sc_hd__nor2_2 _4627_ (.A(_3740_),
    .B(_3781_),
    .Y(_3782_));
 sky130_fd_sc_hd__nor2_2 _4628_ (.A(net139),
    .B(net96),
    .Y(_3783_));
 sky130_fd_sc_hd__nor2_1 _4629_ (.A(net122),
    .B(net93),
    .Y(_3784_));
 sky130_fd_sc_hd__or3_4 _4630_ (.A(net122),
    .B(net94),
    .C(_3713_),
    .X(_3785_));
 sky130_fd_sc_hd__a22o_2 _4631_ (.A1(net124),
    .A2(_3590_),
    .B1(_3602_),
    .B2(net180),
    .X(_3786_));
 sky130_fd_sc_hd__nand3_4 _4632_ (.A(_3783_),
    .B(_3785_),
    .C(_3786_),
    .Y(_3787_));
 sky130_fd_sc_hd__a21o_1 _4633_ (.A1(_3785_),
    .A2(_3786_),
    .B1(_3783_),
    .X(_3788_));
 sky130_fd_sc_hd__nand3_4 _4634_ (.A(_3782_),
    .B(_3787_),
    .C(_3788_),
    .Y(_3789_));
 sky130_fd_sc_hd__a21o_1 _4635_ (.A1(_3787_),
    .A2(_3788_),
    .B1(_3782_),
    .X(_3790_));
 sky130_fd_sc_hd__nand3_2 _4636_ (.A(_3780_),
    .B(_3789_),
    .C(_3790_),
    .Y(_3791_));
 sky130_fd_sc_hd__a21o_1 _4637_ (.A1(_3789_),
    .A2(_3790_),
    .B1(_3780_),
    .X(_3792_));
 sky130_fd_sc_hd__xor2_4 _4638_ (.A(_3775_),
    .B(_3776_),
    .X(_3793_));
 sky130_fd_sc_hd__nand3_2 _4639_ (.A(_3791_),
    .B(_3792_),
    .C(_3793_),
    .Y(_3794_));
 sky130_fd_sc_hd__a21bo_1 _4640_ (.A1(_3792_),
    .A2(_3793_),
    .B1_N(_3791_),
    .X(_3795_));
 sky130_fd_sc_hd__nand2_4 _4641_ (.A(_3785_),
    .B(_3787_),
    .Y(_3796_));
 sky130_fd_sc_hd__nor2_4 _4642_ (.A(net148),
    .B(net68),
    .Y(_3797_));
 sky130_fd_sc_hd__nand2_1 _4643_ (.A(_3796_),
    .B(_3797_),
    .Y(_3798_));
 sky130_fd_sc_hd__xor2_4 _4644_ (.A(_3796_),
    .B(_3797_),
    .X(_3799_));
 sky130_fd_sc_hd__a21o_1 _4645_ (.A1(_3749_),
    .A2(_3750_),
    .B1(_3744_),
    .X(_3800_));
 sky130_fd_sc_hd__nand3b_4 _4646_ (.A_N(_3789_),
    .B(_3800_),
    .C(_3751_),
    .Y(_3801_));
 sky130_fd_sc_hd__a21bo_2 _4647_ (.A1(_3751_),
    .A2(_3800_),
    .B1_N(_3789_),
    .X(_3802_));
 sky130_fd_sc_hd__nand3_4 _4648_ (.A(_3799_),
    .B(_3801_),
    .C(_3802_),
    .Y(_3803_));
 sky130_fd_sc_hd__a21o_1 _4649_ (.A1(_3801_),
    .A2(_3802_),
    .B1(_3799_),
    .X(_3804_));
 sky130_fd_sc_hd__nand3_2 _4650_ (.A(_3795_),
    .B(_3803_),
    .C(_3804_),
    .Y(_3805_));
 sky130_fd_sc_hd__a21o_1 _4651_ (.A1(_3803_),
    .A2(_3804_),
    .B1(_3795_),
    .X(_3806_));
 sky130_fd_sc_hd__nand3_1 _4652_ (.A(_3777_),
    .B(_3805_),
    .C(_3806_),
    .Y(_3807_));
 sky130_fd_sc_hd__a21o_1 _4653_ (.A1(_3805_),
    .A2(_3806_),
    .B1(_3777_),
    .X(_3808_));
 sky130_fd_sc_hd__nor2_1 _4654_ (.A(net122),
    .B(net95),
    .Y(_3809_));
 sky130_fd_sc_hd__nor2_1 _4655_ (.A(net135),
    .B(net95),
    .Y(_3810_));
 sky130_fd_sc_hd__nand2_1 _4656_ (.A(_3784_),
    .B(_3810_),
    .Y(_3811_));
 sky130_fd_sc_hd__xnor2_1 _4657_ (.A(_3784_),
    .B(_3810_),
    .Y(_3812_));
 sky130_fd_sc_hd__nor2_1 _4658_ (.A(_3739_),
    .B(_3812_),
    .Y(_3813_));
 sky130_fd_sc_hd__a21oi_2 _4659_ (.A1(_3774_),
    .A2(_3779_),
    .B1(_3778_),
    .Y(_3814_));
 sky130_fd_sc_hd__or3b_2 _4660_ (.A(_3780_),
    .B(_3814_),
    .C_N(_3813_),
    .X(_3815_));
 sky130_fd_sc_hd__o21bai_2 _4661_ (.A1(_3780_),
    .A2(_3814_),
    .B1_N(_3813_),
    .Y(_3816_));
 sky130_fd_sc_hd__nor2_2 _4662_ (.A(net139),
    .B(net68),
    .Y(_3817_));
 sky130_fd_sc_hd__and3_1 _4663_ (.A(_3784_),
    .B(_3810_),
    .C(_3817_),
    .X(_3818_));
 sky130_fd_sc_hd__xnor2_2 _4664_ (.A(_3811_),
    .B(_3817_),
    .Y(_3819_));
 sky130_fd_sc_hd__nand3_1 _4665_ (.A(_3815_),
    .B(_3816_),
    .C(_3819_),
    .Y(_3820_));
 sky130_fd_sc_hd__a21bo_1 _4666_ (.A1(_3816_),
    .A2(_3819_),
    .B1_N(_3815_),
    .X(_3821_));
 sky130_fd_sc_hd__a21o_1 _4667_ (.A1(_3791_),
    .A2(_3792_),
    .B1(_3793_),
    .X(_3822_));
 sky130_fd_sc_hd__nand3_2 _4668_ (.A(_3794_),
    .B(_3821_),
    .C(_3822_),
    .Y(_3823_));
 sky130_fd_sc_hd__a21o_1 _4669_ (.A1(_3794_),
    .A2(_3822_),
    .B1(_3821_),
    .X(_3824_));
 sky130_fd_sc_hd__nand3_1 _4670_ (.A(_3818_),
    .B(_3823_),
    .C(_3824_),
    .Y(_3825_));
 sky130_fd_sc_hd__a21bo_1 _4671_ (.A1(_3818_),
    .A2(_3824_),
    .B1_N(_3823_),
    .X(_3826_));
 sky130_fd_sc_hd__a21o_2 _4672_ (.A1(_3807_),
    .A2(_3808_),
    .B1(_3826_),
    .X(_3827_));
 sky130_fd_sc_hd__and3_2 _4673_ (.A(_3807_),
    .B(_3808_),
    .C(_3826_),
    .X(_3828_));
 sky130_fd_sc_hd__a21o_1 _4674_ (.A1(_3823_),
    .A2(_3824_),
    .B1(_3818_),
    .X(_3829_));
 sky130_fd_sc_hd__and2_1 _4675_ (.A(_3739_),
    .B(_3812_),
    .X(_3830_));
 sky130_fd_sc_hd__nor2_1 _4676_ (.A(_3813_),
    .B(_3830_),
    .Y(_3831_));
 sky130_fd_sc_hd__nor2_1 _4677_ (.A(net177),
    .B(net68),
    .Y(_3832_));
 sky130_fd_sc_hd__nand2_1 _4678_ (.A(_3770_),
    .B(_3809_),
    .Y(_3833_));
 sky130_fd_sc_hd__and3_1 _4679_ (.A(_3770_),
    .B(_3809_),
    .C(_3832_),
    .X(_3834_));
 sky130_fd_sc_hd__and2b_1 _4680_ (.A_N(_3832_),
    .B(_3833_),
    .X(_3835_));
 sky130_fd_sc_hd__nor2_1 _4681_ (.A(_3834_),
    .B(_3835_),
    .Y(_3836_));
 sky130_fd_sc_hd__and2_2 _4682_ (.A(_3831_),
    .B(_3836_),
    .X(_3837_));
 sky130_fd_sc_hd__a21o_1 _4683_ (.A1(_3815_),
    .A2(_3816_),
    .B1(_3819_),
    .X(_3838_));
 sky130_fd_sc_hd__and2_1 _4684_ (.A(_3820_),
    .B(_3838_),
    .X(_3839_));
 sky130_fd_sc_hd__and3_1 _4685_ (.A(_3820_),
    .B(_3837_),
    .C(_3838_),
    .X(_3840_));
 sky130_fd_sc_hd__a21oi_1 _4686_ (.A1(_3820_),
    .A2(_3838_),
    .B1(_3837_),
    .Y(_3841_));
 sky130_fd_sc_hd__nand2_1 _4687_ (.A(_3834_),
    .B(_3839_),
    .Y(_3842_));
 sky130_fd_sc_hd__o21a_1 _4688_ (.A1(_3834_),
    .A2(_3837_),
    .B1(_3839_),
    .X(_3843_));
 sky130_fd_sc_hd__and3_4 _4689_ (.A(_3825_),
    .B(_3829_),
    .C(_3843_),
    .X(_3844_));
 sky130_fd_sc_hd__nor2_1 _4690_ (.A(_3828_),
    .B(_3844_),
    .Y(_3845_));
 sky130_fd_sc_hd__and2_1 _4691_ (.A(_3827_),
    .B(_3844_),
    .X(_3846_));
 sky130_fd_sc_hd__a21oi_4 _4692_ (.A1(_3827_),
    .A2(_3844_),
    .B1(_3828_),
    .Y(_3847_));
 sky130_fd_sc_hd__o21a_1 _4693_ (.A1(_3754_),
    .A2(_3755_),
    .B1(_3760_),
    .X(_3848_));
 sky130_fd_sc_hd__a211oi_2 _4694_ (.A1(_3801_),
    .A2(_3803_),
    .B1(_3848_),
    .C1(_3761_),
    .Y(_3849_));
 sky130_fd_sc_hd__a211o_2 _4695_ (.A1(_3801_),
    .A2(_3803_),
    .B1(_3848_),
    .C1(_3761_),
    .X(_3850_));
 sky130_fd_sc_hd__o211a_1 _4696_ (.A1(_3761_),
    .A2(_3848_),
    .B1(_3803_),
    .C1(_3801_),
    .X(_3851_));
 sky130_fd_sc_hd__or3_4 _4697_ (.A(_3798_),
    .B(_3849_),
    .C(_3851_),
    .X(_3852_));
 sky130_fd_sc_hd__o21ai_1 _4698_ (.A1(_3849_),
    .A2(_3851_),
    .B1(_3798_),
    .Y(_3853_));
 sky130_fd_sc_hd__a21bo_1 _4699_ (.A1(_3777_),
    .A2(_3806_),
    .B1_N(_3805_),
    .X(_3854_));
 sky130_fd_sc_hd__and3_2 _4700_ (.A(_3852_),
    .B(_3853_),
    .C(_3854_),
    .X(_3855_));
 sky130_fd_sc_hd__a21oi_1 _4701_ (.A1(_3852_),
    .A2(_3853_),
    .B1(_3854_),
    .Y(_3856_));
 sky130_fd_sc_hd__nor2_1 _4702_ (.A(_3855_),
    .B(_3856_),
    .Y(_3857_));
 sky130_fd_sc_hd__or2_4 _4703_ (.A(_3855_),
    .B(_3856_),
    .X(_3858_));
 sky130_fd_sc_hd__a21oi_4 _4704_ (.A1(_3763_),
    .A2(_3765_),
    .B1(_3764_),
    .Y(_3859_));
 sky130_fd_sc_hd__a211oi_4 _4705_ (.A1(_3850_),
    .A2(_3852_),
    .B1(_3859_),
    .C1(_3766_),
    .Y(_3860_));
 sky130_fd_sc_hd__o211a_1 _4706_ (.A1(_3766_),
    .A2(_3859_),
    .B1(_3852_),
    .C1(_3850_),
    .X(_3861_));
 sky130_fd_sc_hd__nor2_1 _4707_ (.A(_3860_),
    .B(_3861_),
    .Y(_3862_));
 sky130_fd_sc_hd__or2_2 _4708_ (.A(_3860_),
    .B(_3861_),
    .X(_3863_));
 sky130_fd_sc_hd__nand2b_1 _4709_ (.A_N(_3861_),
    .B(_3855_),
    .Y(_3864_));
 sky130_fd_sc_hd__o21bai_2 _4710_ (.A1(_3855_),
    .A2(_3860_),
    .B1_N(_3861_),
    .Y(_3865_));
 sky130_fd_sc_hd__a21oi_1 _4711_ (.A1(_3825_),
    .A2(_3829_),
    .B1(_3843_),
    .Y(_3866_));
 sky130_fd_sc_hd__nor2_2 _4712_ (.A(_3844_),
    .B(_3866_),
    .Y(_3867_));
 sky130_fd_sc_hd__o21bai_2 _4713_ (.A1(_3840_),
    .A2(_3841_),
    .B1_N(_3834_),
    .Y(_3868_));
 sky130_fd_sc_hd__nor2_1 _4714_ (.A(_3831_),
    .B(_3836_),
    .Y(_3869_));
 sky130_fd_sc_hd__nor2_1 _4715_ (.A(_3837_),
    .B(_3869_),
    .Y(_3870_));
 sky130_fd_sc_hd__or2_1 _4716_ (.A(_3770_),
    .B(_3809_),
    .X(_3871_));
 sky130_fd_sc_hd__and2_1 _4717_ (.A(_3833_),
    .B(_3871_),
    .X(_3872_));
 sky130_fd_sc_hd__and3_1 _4718_ (.A(net136),
    .B(_3647_),
    .C(_3872_),
    .X(_3873_));
 sky130_fd_sc_hd__and2_1 _4719_ (.A(_3870_),
    .B(_3873_),
    .X(_3874_));
 sky130_fd_sc_hd__and3_1 _4720_ (.A(_3842_),
    .B(_3868_),
    .C(_3874_),
    .X(_3875_));
 sky130_fd_sc_hd__a21oi_1 _4721_ (.A1(_3842_),
    .A2(_3868_),
    .B1(_3874_),
    .Y(_3876_));
 sky130_fd_sc_hd__a21o_1 _4722_ (.A1(_3842_),
    .A2(_3868_),
    .B1(_3874_),
    .X(_3877_));
 sky130_fd_sc_hd__or3b_2 _4723_ (.A(net68),
    .B(net174),
    .C_N(_3809_),
    .X(_3878_));
 sky130_fd_sc_hd__a21oi_1 _4724_ (.A1(net136),
    .A2(_3647_),
    .B1(_3872_),
    .Y(_3879_));
 sky130_fd_sc_hd__or2_1 _4725_ (.A(_3873_),
    .B(_3879_),
    .X(_3880_));
 sky130_fd_sc_hd__nor2_1 _4726_ (.A(_3870_),
    .B(_3873_),
    .Y(_3881_));
 sky130_fd_sc_hd__nor4_2 _4727_ (.A(_3837_),
    .B(_3869_),
    .C(_3878_),
    .D(_3880_),
    .Y(_3882_));
 sky130_fd_sc_hd__and3b_1 _4728_ (.A_N(_3875_),
    .B(_3877_),
    .C(_3882_),
    .X(_3883_));
 sky130_fd_sc_hd__a21o_1 _4729_ (.A1(_3877_),
    .A2(_3882_),
    .B1(_3875_),
    .X(_3884_));
 sky130_fd_sc_hd__nand2_1 _4730_ (.A(_3867_),
    .B(_3884_),
    .Y(_3885_));
 sky130_fd_sc_hd__a311o_4 _4731_ (.A1(_3827_),
    .A2(_3867_),
    .A3(_3884_),
    .B1(_3828_),
    .C1(_3846_),
    .X(_3886_));
 sky130_fd_sc_hd__o31a_2 _4732_ (.A1(_3847_),
    .A2(_3858_),
    .A3(_3863_),
    .B1(_3864_),
    .X(_3887_));
 sky130_fd_sc_hd__o31ai_4 _4733_ (.A1(_3847_),
    .A2(_3858_),
    .A3(_3863_),
    .B1(_3865_),
    .Y(_3888_));
 sky130_fd_sc_hd__a21oi_4 _4734_ (.A1(_3769_),
    .A2(_3888_),
    .B1(_3768_),
    .Y(_3889_));
 sky130_fd_sc_hd__and2b_2 _4735_ (.A_N(_3735_),
    .B(_3736_),
    .X(_3890_));
 sky130_fd_sc_hd__o21a_1 _4736_ (.A1(_3735_),
    .A2(_3768_),
    .B1(_3736_),
    .X(_3891_));
 sky130_fd_sc_hd__a31o_2 _4737_ (.A1(_3769_),
    .A2(_3888_),
    .A3(_3890_),
    .B1(_3891_),
    .X(_3892_));
 sky130_fd_sc_hd__xnor2_4 _4738_ (.A(_3700_),
    .B(_3892_),
    .Y(_3893_));
 sky130_fd_sc_hd__nor2_8 _4739_ (.A(net211),
    .B(net59),
    .Y(_3894_));
 sky130_fd_sc_hd__nand2_2 _4740_ (.A(net120),
    .B(_3894_),
    .Y(_3895_));
 sky130_fd_sc_hd__or3_4 _4741_ (.A(net210),
    .B(_3539_),
    .C(net58),
    .X(_3896_));
 sky130_fd_sc_hd__and3_2 _4742_ (.A(net115),
    .B(_3590_),
    .C(_3894_),
    .X(_3897_));
 sky130_fd_sc_hd__or4_4 _4743_ (.A(net210),
    .B(_3539_),
    .C(net114),
    .D(net59),
    .X(_3898_));
 sky130_fd_sc_hd__a211oi_4 _4744_ (.A1(_3539_),
    .A2(_3589_),
    .B1(net59),
    .C1(net210),
    .Y(_3899_));
 sky130_fd_sc_hd__nand4_4 _4745_ (.A(net117),
    .B(_3894_),
    .C(_3898_),
    .D(_3899_),
    .Y(_3900_));
 sky130_fd_sc_hd__and3_4 _4746_ (.A(_3895_),
    .B(_3898_),
    .C(_3900_),
    .X(_3901_));
 sky130_fd_sc_hd__a21oi_2 _4747_ (.A1(_3898_),
    .A2(_3900_),
    .B1(_3895_),
    .Y(_3902_));
 sky130_fd_sc_hd__nor2_2 _4748_ (.A(_3901_),
    .B(_3902_),
    .Y(_3903_));
 sky130_fd_sc_hd__or3_4 _4749_ (.A(net211),
    .B(net59),
    .C(_3903_),
    .X(_3904_));
 sky130_fd_sc_hd__a22o_1 _4750_ (.A1(net115),
    .A2(net59),
    .B1(_3894_),
    .B2(_3590_),
    .X(_3905_));
 sky130_fd_sc_hd__or4b_4 _4751_ (.A(net210),
    .B(_3589_),
    .C(net59),
    .D_N(net117),
    .X(_3906_));
 sky130_fd_sc_hd__inv_2 _4752_ (.A(_3906_),
    .Y(_3907_));
 sky130_fd_sc_hd__a21o_1 _4753_ (.A1(net119),
    .A2(_3894_),
    .B1(_3905_),
    .X(_3908_));
 sky130_fd_sc_hd__nand2_2 _4754_ (.A(_3906_),
    .B(_3908_),
    .Y(_3909_));
 sky130_fd_sc_hd__or2_1 _4755_ (.A(_3904_),
    .B(_3909_),
    .X(_3910_));
 sky130_fd_sc_hd__a22o_1 _4756_ (.A1(_3590_),
    .A2(net59),
    .B1(_3894_),
    .B2(net117),
    .X(_3911_));
 sky130_fd_sc_hd__nand2_1 _4757_ (.A(_3506_),
    .B(_3906_),
    .Y(_3912_));
 sky130_fd_sc_hd__o21ai_1 _4758_ (.A1(_3895_),
    .A2(_3906_),
    .B1(_3912_),
    .Y(_3913_));
 sky130_fd_sc_hd__nand2_1 _4759_ (.A(_3894_),
    .B(_3913_),
    .Y(_3914_));
 sky130_fd_sc_hd__nand2b_1 _4760_ (.A_N(_3914_),
    .B(_3911_),
    .Y(_3915_));
 sky130_fd_sc_hd__xor2_1 _4761_ (.A(_3911_),
    .B(_3914_),
    .X(_3916_));
 sky130_fd_sc_hd__or2_2 _4762_ (.A(_3910_),
    .B(_3916_),
    .X(_3917_));
 sky130_fd_sc_hd__nand2_1 _4763_ (.A(_3910_),
    .B(_3916_),
    .Y(_3918_));
 sky130_fd_sc_hd__nand2_1 _4764_ (.A(_3917_),
    .B(_3918_),
    .Y(_3919_));
 sky130_fd_sc_hd__or2_2 _4765_ (.A(_3901_),
    .B(_3919_),
    .X(_3920_));
 sky130_fd_sc_hd__nand2_1 _4766_ (.A(_3901_),
    .B(_3919_),
    .Y(_3921_));
 sky130_fd_sc_hd__and2_1 _4767_ (.A(_3920_),
    .B(_3921_),
    .X(_3922_));
 sky130_fd_sc_hd__xor2_2 _4768_ (.A(_3904_),
    .B(_3909_),
    .X(_3923_));
 sky130_fd_sc_hd__a22o_2 _4769_ (.A1(net117),
    .A2(_3894_),
    .B1(_3898_),
    .B2(_3899_),
    .X(_3924_));
 sky130_fd_sc_hd__and2_4 _4770_ (.A(_3900_),
    .B(_3924_),
    .X(_3925_));
 sky130_fd_sc_hd__or3_4 _4771_ (.A(net210),
    .B(net93),
    .C(net58),
    .X(_3926_));
 sky130_fd_sc_hd__nand2_1 _4772_ (.A(_3647_),
    .B(net58),
    .Y(_3927_));
 sky130_fd_sc_hd__or4_4 _4773_ (.A(net210),
    .B(net95),
    .C(net93),
    .D(net58),
    .X(_3928_));
 sky130_fd_sc_hd__a21bo_1 _4774_ (.A1(_3582_),
    .A2(net58),
    .B1_N(_3926_),
    .X(_3929_));
 sky130_fd_sc_hd__nand4_2 _4775_ (.A(_3900_),
    .B(_3924_),
    .C(_3928_),
    .D(_3929_),
    .Y(_3930_));
 sky130_fd_sc_hd__a22oi_2 _4776_ (.A1(net92),
    .A2(net59),
    .B1(_3900_),
    .B2(_3924_),
    .Y(_3931_));
 sky130_fd_sc_hd__a21oi_1 _4777_ (.A1(_3928_),
    .A2(_3930_),
    .B1(_3931_),
    .Y(_3932_));
 sky130_fd_sc_hd__and2_1 _4778_ (.A(_3928_),
    .B(_3931_),
    .X(_3933_));
 sky130_fd_sc_hd__nor2_2 _4779_ (.A(_3932_),
    .B(_3933_),
    .Y(_3934_));
 sky130_fd_sc_hd__o21ba_1 _4780_ (.A1(_3904_),
    .A2(_3933_),
    .B1_N(_3932_),
    .X(_3935_));
 sky130_fd_sc_hd__and2b_1 _4781_ (.A_N(_3935_),
    .B(_3923_),
    .X(_3936_));
 sky130_fd_sc_hd__xnor2_1 _4782_ (.A(_3923_),
    .B(_3935_),
    .Y(_3937_));
 sky130_fd_sc_hd__and2b_1 _4783_ (.A_N(_3901_),
    .B(_3937_),
    .X(_3938_));
 sky130_fd_sc_hd__o21ai_2 _4784_ (.A1(_3936_),
    .A2(_3938_),
    .B1(_3922_),
    .Y(_3939_));
 sky130_fd_sc_hd__or3_1 _4785_ (.A(_3922_),
    .B(_3936_),
    .C(_3938_),
    .X(_3940_));
 sky130_fd_sc_hd__nand2_1 _4786_ (.A(_3939_),
    .B(_3940_),
    .Y(_3941_));
 sky130_fd_sc_hd__inv_2 _4787_ (.A(_3941_),
    .Y(_3942_));
 sky130_fd_sc_hd__and2b_1 _4788_ (.A_N(_3937_),
    .B(_3901_),
    .X(_3943_));
 sky130_fd_sc_hd__nor2_1 _4789_ (.A(_3938_),
    .B(_3943_),
    .Y(_3944_));
 sky130_fd_sc_hd__xnor2_4 _4790_ (.A(_3904_),
    .B(_3934_),
    .Y(_3945_));
 sky130_fd_sc_hd__a22o_1 _4791_ (.A1(_3900_),
    .A2(_3924_),
    .B1(_3928_),
    .B2(_3929_),
    .X(_3946_));
 sky130_fd_sc_hd__nand2_1 _4792_ (.A(_3930_),
    .B(_3946_),
    .Y(_3947_));
 sky130_fd_sc_hd__o211a_1 _4793_ (.A1(_3686_),
    .A2(net58),
    .B1(_3926_),
    .C1(_3927_),
    .X(_3948_));
 sky130_fd_sc_hd__nor2_4 _4794_ (.A(_3669_),
    .B(net58),
    .Y(_3949_));
 sky130_fd_sc_hd__or3_4 _4795_ (.A(_3669_),
    .B(_3686_),
    .C(net58),
    .X(_3950_));
 sky130_fd_sc_hd__a21o_2 _4796_ (.A1(_3669_),
    .A2(_3686_),
    .B1(net58),
    .X(_3951_));
 sky130_fd_sc_hd__a21oi_2 _4797_ (.A1(_3669_),
    .A2(_3686_),
    .B1(net58),
    .Y(_3952_));
 sky130_fd_sc_hd__or3b_1 _4798_ (.A(_3951_),
    .B(_3926_),
    .C_N(_3950_),
    .X(_3953_));
 sky130_fd_sc_hd__o21ai_4 _4799_ (.A1(_3926_),
    .A2(_3951_),
    .B1(_3950_),
    .Y(_3954_));
 sky130_fd_sc_hd__nand2_1 _4800_ (.A(_3928_),
    .B(_3954_),
    .Y(_3955_));
 sky130_fd_sc_hd__a21oi_4 _4801_ (.A1(_3928_),
    .A2(_3954_),
    .B1(_3948_),
    .Y(_3956_));
 sky130_fd_sc_hd__nand2_1 _4802_ (.A(_3925_),
    .B(_3956_),
    .Y(_3957_));
 sky130_fd_sc_hd__a21bo_1 _4803_ (.A1(_3925_),
    .A2(_3956_),
    .B1_N(_3955_),
    .X(_3958_));
 sky130_fd_sc_hd__nand2b_1 _4804_ (.A_N(_3947_),
    .B(_3958_),
    .Y(_3959_));
 sky130_fd_sc_hd__and3_1 _4805_ (.A(_3947_),
    .B(_3955_),
    .C(_3957_),
    .X(_3960_));
 sky130_fd_sc_hd__xnor2_1 _4806_ (.A(_3947_),
    .B(_3958_),
    .Y(_3961_));
 sky130_fd_sc_hd__o21a_1 _4807_ (.A1(_3904_),
    .A2(_3960_),
    .B1(_3959_),
    .X(_3962_));
 sky130_fd_sc_hd__and2b_1 _4808_ (.A_N(_3962_),
    .B(_3945_),
    .X(_3963_));
 sky130_fd_sc_hd__xor2_2 _4809_ (.A(_3945_),
    .B(_3962_),
    .X(_3964_));
 sky130_fd_sc_hd__nor2_2 _4810_ (.A(_3901_),
    .B(_3964_),
    .Y(_3965_));
 sky130_fd_sc_hd__o21a_1 _4811_ (.A1(_3963_),
    .A2(_3965_),
    .B1(_3944_),
    .X(_3966_));
 sky130_fd_sc_hd__inv_2 _4812_ (.A(_3966_),
    .Y(_3967_));
 sky130_fd_sc_hd__nor3_1 _4813_ (.A(_3944_),
    .B(_3963_),
    .C(_3965_),
    .Y(_3968_));
 sky130_fd_sc_hd__or2_4 _4814_ (.A(_3966_),
    .B(_3968_),
    .X(_3969_));
 sky130_fd_sc_hd__and2_1 _4815_ (.A(_3901_),
    .B(_3964_),
    .X(_3970_));
 sky130_fd_sc_hd__nor2_2 _4816_ (.A(_3965_),
    .B(_3970_),
    .Y(_3971_));
 sky130_fd_sc_hd__xnor2_1 _4817_ (.A(_3904_),
    .B(_3961_),
    .Y(_3972_));
 sky130_fd_sc_hd__nor2_1 _4818_ (.A(_3925_),
    .B(_3956_),
    .Y(_3973_));
 sky130_fd_sc_hd__nor2_8 _4819_ (.A(net93),
    .B(_3950_),
    .Y(_3974_));
 sky130_fd_sc_hd__mux2_8 _4820_ (.A0(_3950_),
    .A1(_3952_),
    .S(_3926_),
    .X(_3975_));
 sky130_fd_sc_hd__a21o_2 _4821_ (.A1(_3926_),
    .A2(_3951_),
    .B1(_3974_),
    .X(_3976_));
 sky130_fd_sc_hd__a21o_1 _4822_ (.A1(_3925_),
    .A2(_3975_),
    .B1(_3974_),
    .X(_3977_));
 sky130_fd_sc_hd__a21o_1 _4823_ (.A1(_3957_),
    .A2(_3977_),
    .B1(_3973_),
    .X(_3978_));
 sky130_fd_sc_hd__a2bb2o_1 _4824_ (.A1_N(_3904_),
    .A2_N(_3973_),
    .B1(_3977_),
    .B2(_3957_),
    .X(_3979_));
 sky130_fd_sc_hd__and2_2 _4825_ (.A(_3972_),
    .B(_3979_),
    .X(_3980_));
 sky130_fd_sc_hd__xnor2_1 _4826_ (.A(_3972_),
    .B(_3979_),
    .Y(_3981_));
 sky130_fd_sc_hd__nor2_2 _4827_ (.A(_3901_),
    .B(_3981_),
    .Y(_3982_));
 sky130_fd_sc_hd__o21ai_4 _4828_ (.A1(_3980_),
    .A2(_3982_),
    .B1(_3971_),
    .Y(_3983_));
 sky130_fd_sc_hd__or3_2 _4829_ (.A(_3971_),
    .B(_3980_),
    .C(_3982_),
    .X(_3984_));
 sky130_fd_sc_hd__nand2_4 _4830_ (.A(_3983_),
    .B(_3984_),
    .Y(_3985_));
 sky130_fd_sc_hd__or2_1 _4831_ (.A(_3969_),
    .B(_3985_),
    .X(_3986_));
 sky130_fd_sc_hd__and2_1 _4832_ (.A(_3901_),
    .B(_3981_),
    .X(_3987_));
 sky130_fd_sc_hd__nor2_1 _4833_ (.A(_3982_),
    .B(_3987_),
    .Y(_3988_));
 sky130_fd_sc_hd__xnor2_1 _4834_ (.A(_3925_),
    .B(_3975_),
    .Y(_3989_));
 sky130_fd_sc_hd__nand2_2 _4835_ (.A(_3925_),
    .B(_3974_),
    .Y(_3990_));
 sky130_fd_sc_hd__xnor2_4 _4836_ (.A(_3858_),
    .B(_3886_),
    .Y(_3991_));
 sky130_fd_sc_hd__and2_1 _4837_ (.A(_3878_),
    .B(_3880_),
    .X(_3992_));
 sky130_fd_sc_hd__o221a_1 _4838_ (.A1(_3875_),
    .A2(_3876_),
    .B1(_3881_),
    .B2(_3874_),
    .C1(_3992_),
    .X(_3993_));
 sky130_fd_sc_hd__a21o_1 _4839_ (.A1(net122),
    .A2(net174),
    .B1(net68),
    .X(_3994_));
 sky130_fd_sc_hd__o221a_1 _4840_ (.A1(net95),
    .A2(net174),
    .B1(_3883_),
    .B2(_3993_),
    .C1(_3994_),
    .X(_3995_));
 sky130_fd_sc_hd__a211o_1 _4841_ (.A1(_3827_),
    .A2(_3845_),
    .B1(_3867_),
    .C1(_3884_),
    .X(_3996_));
 sky130_fd_sc_hd__a21bo_4 _4842_ (.A1(_3885_),
    .A2(_3996_),
    .B1_N(_3995_),
    .X(_3997_));
 sky130_fd_sc_hd__nor2_1 _4843_ (.A(_3991_),
    .B(net60),
    .Y(_3998_));
 sky130_fd_sc_hd__a211o_2 _4844_ (.A1(_3857_),
    .A2(_3886_),
    .B1(_3862_),
    .C1(_3855_),
    .X(_3999_));
 sky130_fd_sc_hd__a211o_4 _4845_ (.A1(_3887_),
    .A2(_3999_),
    .B1(net60),
    .C1(_3991_),
    .X(_4000_));
 sky130_fd_sc_hd__xor2_4 _4846_ (.A(_3769_),
    .B(_3888_),
    .X(_4001_));
 sky130_fd_sc_hd__a2111o_4 _4847_ (.A1(_3887_),
    .A2(_3999_),
    .B1(_4001_),
    .C1(_3991_),
    .D1(net60),
    .X(_4002_));
 sky130_fd_sc_hd__xnor2_4 _4848_ (.A(_3889_),
    .B(_3890_),
    .Y(_4003_));
 sky130_fd_sc_hd__a21oi_4 _4849_ (.A1(_4002_),
    .A2(_4003_),
    .B1(net210),
    .Y(_0075_));
 sky130_fd_sc_hd__xor2_2 _4850_ (.A(_3903_),
    .B(_0075_),
    .X(_0076_));
 sky130_fd_sc_hd__or3_1 _4851_ (.A(_3925_),
    .B(_3974_),
    .C(_3975_),
    .X(_0077_));
 sky130_fd_sc_hd__and2_1 _4852_ (.A(_3990_),
    .B(_0077_),
    .X(_0078_));
 sky130_fd_sc_hd__nand2_2 _4853_ (.A(_0076_),
    .B(_0078_),
    .Y(_0079_));
 sky130_fd_sc_hd__xnor2_2 _4854_ (.A(_3904_),
    .B(_3978_),
    .Y(_0080_));
 sky130_fd_sc_hd__a21oi_4 _4855_ (.A1(_3990_),
    .A2(_0079_),
    .B1(_0080_),
    .Y(_0081_));
 sky130_fd_sc_hd__a21o_2 _4856_ (.A1(_3903_),
    .A2(net57),
    .B1(_3902_),
    .X(_0082_));
 sky130_fd_sc_hd__and3_1 _4857_ (.A(_3990_),
    .B(_0079_),
    .C(_0080_),
    .X(_0083_));
 sky130_fd_sc_hd__nor2_2 _4858_ (.A(_0081_),
    .B(_0083_),
    .Y(_0084_));
 sky130_fd_sc_hd__and2_1 _4859_ (.A(_0082_),
    .B(_0084_),
    .X(_0085_));
 sky130_fd_sc_hd__nor3_1 _4860_ (.A(_3988_),
    .B(_0081_),
    .C(_0085_),
    .Y(_0086_));
 sky130_fd_sc_hd__o21ai_2 _4861_ (.A1(_0081_),
    .A2(_0085_),
    .B1(_3988_),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _4862_ (.A(_0087_),
    .Y(_0088_));
 sky130_fd_sc_hd__nand2b_2 _4863_ (.A_N(_0086_),
    .B(_0087_),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _4864_ (.A(_0089_),
    .Y(_0090_));
 sky130_fd_sc_hd__xnor2_2 _4865_ (.A(_0082_),
    .B(_0084_),
    .Y(_0091_));
 sky130_fd_sc_hd__or2_1 _4866_ (.A(_0076_),
    .B(_0078_),
    .X(_0092_));
 sky130_fd_sc_hd__and2_2 _4867_ (.A(_0079_),
    .B(_0092_),
    .X(_0093_));
 sky130_fd_sc_hd__and4_1 _4868_ (.A(net117),
    .B(_3898_),
    .C(_3899_),
    .D(_0075_),
    .X(_0094_));
 sky130_fd_sc_hd__a22o_1 _4869_ (.A1(_3898_),
    .A2(_3899_),
    .B1(_0075_),
    .B2(net117),
    .X(_0095_));
 sky130_fd_sc_hd__and2b_2 _4870_ (.A_N(_0094_),
    .B(_0095_),
    .X(_0096_));
 sky130_fd_sc_hd__a21oi_1 _4871_ (.A1(_3975_),
    .A2(_0096_),
    .B1(_3974_),
    .Y(_0097_));
 sky130_fd_sc_hd__nor2_1 _4872_ (.A(_3989_),
    .B(_0097_),
    .Y(_0098_));
 sky130_fd_sc_hd__xnor2_4 _4873_ (.A(_4000_),
    .B(_4001_),
    .Y(_0099_));
 sky130_fd_sc_hd__or2_4 _4874_ (.A(_3897_),
    .B(_0094_),
    .X(_0100_));
 sky130_fd_sc_hd__nand2_2 _4875_ (.A(net120),
    .B(net57),
    .Y(_0101_));
 sky130_fd_sc_hd__xnor2_4 _4876_ (.A(_0100_),
    .B(_0101_),
    .Y(_0102_));
 sky130_fd_sc_hd__and2b_1 _4877_ (.A_N(_0099_),
    .B(_0102_),
    .X(_0103_));
 sky130_fd_sc_hd__xnor2_4 _4878_ (.A(_0099_),
    .B(_0102_),
    .Y(_0104_));
 sky130_fd_sc_hd__nand2_1 _4879_ (.A(_3989_),
    .B(_0097_),
    .Y(_0105_));
 sky130_fd_sc_hd__nand2b_2 _4880_ (.A_N(_0098_),
    .B(_0105_),
    .Y(_0106_));
 sky130_fd_sc_hd__a21o_2 _4881_ (.A1(_0104_),
    .A2(_0105_),
    .B1(_0098_),
    .X(_0107_));
 sky130_fd_sc_hd__nand2_1 _4882_ (.A(_0093_),
    .B(_0107_),
    .Y(_0108_));
 sky130_fd_sc_hd__a31o_4 _4883_ (.A1(net120),
    .A2(net57),
    .A3(_0100_),
    .B1(_0103_),
    .X(_0109_));
 sky130_fd_sc_hd__xor2_4 _4884_ (.A(_0093_),
    .B(_0107_),
    .X(_0110_));
 sky130_fd_sc_hd__a21boi_4 _4885_ (.A1(_0109_),
    .A2(_0110_),
    .B1_N(_0108_),
    .Y(_0111_));
 sky130_fd_sc_hd__nor2_4 _4886_ (.A(_0091_),
    .B(_0111_),
    .Y(_0112_));
 sky130_fd_sc_hd__and2_1 _4887_ (.A(_0091_),
    .B(_0111_),
    .X(_0113_));
 sky130_fd_sc_hd__or2_4 _4888_ (.A(_0112_),
    .B(_0113_),
    .X(_0114_));
 sky130_fd_sc_hd__a211o_4 _4889_ (.A1(_4002_),
    .A2(_4003_),
    .B1(net210),
    .C1(net114),
    .X(_0115_));
 sky130_fd_sc_hd__xnor2_4 _4890_ (.A(_3896_),
    .B(_0115_),
    .Y(_0116_));
 sky130_fd_sc_hd__nand2b_4 _4891_ (.A_N(net56),
    .B(net117),
    .Y(_0117_));
 sky130_fd_sc_hd__xnor2_4 _4892_ (.A(_0116_),
    .B(_0117_),
    .Y(_0118_));
 sky130_fd_sc_hd__o21ba_1 _4893_ (.A1(_3976_),
    .A2(_0118_),
    .B1_N(_3974_),
    .X(_0119_));
 sky130_fd_sc_hd__xnor2_2 _4894_ (.A(_3976_),
    .B(_0096_),
    .Y(_0120_));
 sky130_fd_sc_hd__nand2b_1 _4895_ (.A_N(_0119_),
    .B(_0120_),
    .Y(_0121_));
 sky130_fd_sc_hd__o211ai_1 _4896_ (.A1(_3991_),
    .A2(net60),
    .B1(_3999_),
    .C1(_3887_),
    .Y(_0122_));
 sky130_fd_sc_hd__and2_2 _4897_ (.A(_4000_),
    .B(_0122_),
    .X(_0123_));
 sky130_fd_sc_hd__o2bb2a_4 _4898_ (.A1_N(_3897_),
    .A2_N(net57),
    .B1(_0116_),
    .B2(_0117_),
    .X(_0124_));
 sky130_fd_sc_hd__nor2_1 _4899_ (.A(_3506_),
    .B(net56),
    .Y(_0125_));
 sky130_fd_sc_hd__xnor2_2 _4900_ (.A(_0124_),
    .B(_0125_),
    .Y(_0126_));
 sky130_fd_sc_hd__nand2_1 _4901_ (.A(net55),
    .B(_0126_),
    .Y(_0127_));
 sky130_fd_sc_hd__xor2_2 _4902_ (.A(net55),
    .B(_0126_),
    .X(_0128_));
 sky130_fd_sc_hd__xnor2_1 _4903_ (.A(_0119_),
    .B(_0120_),
    .Y(_0129_));
 sky130_fd_sc_hd__nand2_2 _4904_ (.A(_0128_),
    .B(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__nand2_4 _4905_ (.A(_0121_),
    .B(_0130_),
    .Y(_0131_));
 sky130_fd_sc_hd__xor2_4 _4906_ (.A(_0104_),
    .B(_0106_),
    .X(_0132_));
 sky130_fd_sc_hd__nand2b_1 _4907_ (.A_N(_0132_),
    .B(_0131_),
    .Y(_0133_));
 sky130_fd_sc_hd__o31ai_4 _4908_ (.A1(_3506_),
    .A2(net56),
    .A3(_0124_),
    .B1(_0127_),
    .Y(_0134_));
 sky130_fd_sc_hd__xor2_4 _4909_ (.A(_0131_),
    .B(_0132_),
    .X(_0135_));
 sky130_fd_sc_hd__nand2b_1 _4910_ (.A_N(_0135_),
    .B(_0134_),
    .Y(_0136_));
 sky130_fd_sc_hd__xnor2_2 _4911_ (.A(_0109_),
    .B(_0110_),
    .Y(_0137_));
 sky130_fd_sc_hd__a21oi_2 _4912_ (.A1(_0133_),
    .A2(_0136_),
    .B1(_0137_),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _4913_ (.A(_0138_),
    .Y(_0139_));
 sky130_fd_sc_hd__and3_1 _4914_ (.A(_0133_),
    .B(_0136_),
    .C(_0137_),
    .X(_0140_));
 sky130_fd_sc_hd__or2_4 _4915_ (.A(_0138_),
    .B(_0140_),
    .X(_0141_));
 sky130_fd_sc_hd__xor2_4 _4916_ (.A(_0134_),
    .B(_0135_),
    .X(_0142_));
 sky130_fd_sc_hd__a2bb2o_2 _4917_ (.A1_N(net114),
    .A2_N(net56),
    .B1(net57),
    .B2(net115),
    .X(_0143_));
 sky130_fd_sc_hd__or2_4 _4918_ (.A(_3539_),
    .B(_0099_),
    .X(_0144_));
 sky130_fd_sc_hd__or3_4 _4919_ (.A(_3539_),
    .B(net56),
    .C(_0115_),
    .X(_0145_));
 sky130_fd_sc_hd__and2_2 _4920_ (.A(net119),
    .B(net55),
    .X(_0146_));
 sky130_fd_sc_hd__nand3_4 _4921_ (.A(_0143_),
    .B(_0145_),
    .C(_0146_),
    .Y(_0147_));
 sky130_fd_sc_hd__a21o_1 _4922_ (.A1(_0143_),
    .A2(_0145_),
    .B1(_0146_),
    .X(_0148_));
 sky130_fd_sc_hd__and4_1 _4923_ (.A(net92),
    .B(_3950_),
    .C(_3952_),
    .D(net57),
    .X(_0149_));
 sky130_fd_sc_hd__a21o_1 _4924_ (.A1(_3953_),
    .A2(_3975_),
    .B1(_0149_),
    .X(_0150_));
 sky130_fd_sc_hd__and3_2 _4925_ (.A(_0147_),
    .B(_0148_),
    .C(_0150_),
    .X(_0151_));
 sky130_fd_sc_hd__nor2_4 _4926_ (.A(_3974_),
    .B(_0151_),
    .Y(_0152_));
 sky130_fd_sc_hd__xnor2_4 _4927_ (.A(_3975_),
    .B(_0118_),
    .Y(_0153_));
 sky130_fd_sc_hd__and2b_1 _4928_ (.A_N(_0152_),
    .B(_0153_),
    .X(_0154_));
 sky130_fd_sc_hd__and2_1 _4929_ (.A(_3991_),
    .B(net60),
    .X(_0155_));
 sky130_fd_sc_hd__or2_4 _4930_ (.A(_3998_),
    .B(_0155_),
    .X(_0156_));
 sky130_fd_sc_hd__nand2_4 _4931_ (.A(_0145_),
    .B(_0147_),
    .Y(_0157_));
 sky130_fd_sc_hd__nand2_2 _4932_ (.A(net120),
    .B(net55),
    .Y(_0158_));
 sky130_fd_sc_hd__xnor2_4 _4933_ (.A(_0157_),
    .B(_0158_),
    .Y(_0159_));
 sky130_fd_sc_hd__and2b_1 _4934_ (.A_N(_0156_),
    .B(_0159_),
    .X(_0160_));
 sky130_fd_sc_hd__xnor2_4 _4935_ (.A(_0156_),
    .B(_0159_),
    .Y(_0161_));
 sky130_fd_sc_hd__xnor2_4 _4936_ (.A(_0152_),
    .B(_0153_),
    .Y(_0162_));
 sky130_fd_sc_hd__a21oi_4 _4937_ (.A1(_0161_),
    .A2(_0162_),
    .B1(_0154_),
    .Y(_0163_));
 sky130_fd_sc_hd__or2_1 _4938_ (.A(_0128_),
    .B(_0129_),
    .X(_0164_));
 sky130_fd_sc_hd__nand2_2 _4939_ (.A(_0130_),
    .B(_0164_),
    .Y(_0165_));
 sky130_fd_sc_hd__nor2_1 _4940_ (.A(_0163_),
    .B(_0165_),
    .Y(_0166_));
 sky130_fd_sc_hd__a31o_4 _4941_ (.A1(net120),
    .A2(net55),
    .A3(_0157_),
    .B1(_0160_),
    .X(_0167_));
 sky130_fd_sc_hd__xor2_4 _4942_ (.A(_0163_),
    .B(_0165_),
    .X(_0168_));
 sky130_fd_sc_hd__a21oi_4 _4943_ (.A1(_0167_),
    .A2(_0168_),
    .B1(_0166_),
    .Y(_0169_));
 sky130_fd_sc_hd__or2_1 _4944_ (.A(_0142_),
    .B(_0169_),
    .X(_0170_));
 sky130_fd_sc_hd__xnor2_2 _4945_ (.A(_0142_),
    .B(_0169_),
    .Y(_0171_));
 sky130_fd_sc_hd__a211o_4 _4946_ (.A1(_4002_),
    .A2(_4003_),
    .B1(net210),
    .C1(net95),
    .X(_0172_));
 sky130_fd_sc_hd__and3_1 _4947_ (.A(_3582_),
    .B(_3949_),
    .C(net57),
    .X(_0173_));
 sky130_fd_sc_hd__nor2_4 _4948_ (.A(net93),
    .B(net56),
    .Y(_0174_));
 sky130_fd_sc_hd__xnor2_4 _4949_ (.A(_3949_),
    .B(_0172_),
    .Y(_0175_));
 sky130_fd_sc_hd__a21o_2 _4950_ (.A1(_0174_),
    .A2(_0175_),
    .B1(_0173_),
    .X(_0176_));
 sky130_fd_sc_hd__a22o_1 _4951_ (.A1(_3950_),
    .A2(_3952_),
    .B1(net57),
    .B2(net92),
    .X(_0177_));
 sky130_fd_sc_hd__and2b_2 _4952_ (.A_N(_0149_),
    .B(_0177_),
    .X(_0178_));
 sky130_fd_sc_hd__and2_1 _4953_ (.A(_0176_),
    .B(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__nand2_4 _4954_ (.A(_3590_),
    .B(net55),
    .Y(_0180_));
 sky130_fd_sc_hd__nand2_2 _4955_ (.A(net115),
    .B(net55),
    .Y(_0181_));
 sky130_fd_sc_hd__or2_1 _4956_ (.A(_0144_),
    .B(_0180_),
    .X(_0182_));
 sky130_fd_sc_hd__xnor2_4 _4957_ (.A(_0144_),
    .B(_0180_),
    .Y(_0183_));
 sky130_fd_sc_hd__nand2b_4 _4958_ (.A_N(_0156_),
    .B(net117),
    .Y(_0184_));
 sky130_fd_sc_hd__xor2_4 _4959_ (.A(_0183_),
    .B(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__xor2_4 _4960_ (.A(_0176_),
    .B(_0178_),
    .X(_0186_));
 sky130_fd_sc_hd__a21oi_4 _4961_ (.A1(_0185_),
    .A2(_0186_),
    .B1(_0179_),
    .Y(_0187_));
 sky130_fd_sc_hd__a21oi_2 _4962_ (.A1(_0147_),
    .A2(_0148_),
    .B1(_0150_),
    .Y(_0188_));
 sky130_fd_sc_hd__nor2_4 _4963_ (.A(_0151_),
    .B(_0188_),
    .Y(_0189_));
 sky130_fd_sc_hd__and2b_1 _4964_ (.A_N(_0187_),
    .B(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__xnor2_4 _4965_ (.A(_0187_),
    .B(_0189_),
    .Y(_0191_));
 sky130_fd_sc_hd__o21a_4 _4966_ (.A1(_0183_),
    .A2(_0184_),
    .B1(_0182_),
    .X(_0192_));
 sky130_fd_sc_hd__or2_4 _4967_ (.A(_3506_),
    .B(_0156_),
    .X(_0193_));
 sky130_fd_sc_hd__xor2_4 _4968_ (.A(_0192_),
    .B(_0193_),
    .X(_0194_));
 sky130_fd_sc_hd__xor2_4 _4969_ (.A(_3997_),
    .B(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__a21o_2 _4970_ (.A1(_0191_),
    .A2(_0195_),
    .B1(_0190_),
    .X(_0196_));
 sky130_fd_sc_hd__xor2_4 _4971_ (.A(_0161_),
    .B(_0162_),
    .X(_0197_));
 sky130_fd_sc_hd__nand2_1 _4972_ (.A(_0196_),
    .B(_0197_),
    .Y(_0198_));
 sky130_fd_sc_hd__a2bb2o_4 _4973_ (.A1_N(_0192_),
    .A2_N(_0193_),
    .B1(_0194_),
    .B2(_3997_),
    .X(_0199_));
 sky130_fd_sc_hd__xnor2_4 _4974_ (.A(_0196_),
    .B(_0197_),
    .Y(_0200_));
 sky130_fd_sc_hd__nand2b_1 _4975_ (.A_N(_0200_),
    .B(_0199_),
    .Y(_0201_));
 sky130_fd_sc_hd__xnor2_2 _4976_ (.A(_0167_),
    .B(_0168_),
    .Y(_0202_));
 sky130_fd_sc_hd__a21oi_1 _4977_ (.A1(_0198_),
    .A2(_0201_),
    .B1(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__a21o_1 _4978_ (.A1(_0198_),
    .A2(_0201_),
    .B1(_0202_),
    .X(_0204_));
 sky130_fd_sc_hd__and3_2 _4979_ (.A(_0198_),
    .B(_0201_),
    .C(_0202_),
    .X(_0205_));
 sky130_fd_sc_hd__xor2_4 _4980_ (.A(_0199_),
    .B(_0200_),
    .X(_0206_));
 sky130_fd_sc_hd__or4b_2 _4981_ (.A(net95),
    .B(net56),
    .C(net68),
    .D_N(net57),
    .X(_0207_));
 sky130_fd_sc_hd__and2_2 _4982_ (.A(net92),
    .B(net55),
    .X(_0208_));
 sky130_fd_sc_hd__a2bb2o_2 _4983_ (.A1_N(net95),
    .A2_N(net56),
    .B1(_3647_),
    .B2(net57),
    .X(_0209_));
 sky130_fd_sc_hd__nand3_1 _4984_ (.A(_0207_),
    .B(_0208_),
    .C(_0209_),
    .Y(_0210_));
 sky130_fd_sc_hd__a21bo_4 _4985_ (.A1(_0208_),
    .A2(_0209_),
    .B1_N(_0207_),
    .X(_0211_));
 sky130_fd_sc_hd__xnor2_4 _4986_ (.A(_0174_),
    .B(_0175_),
    .Y(_0212_));
 sky130_fd_sc_hd__nand2b_2 _4987_ (.A_N(_0212_),
    .B(_0211_),
    .Y(_0213_));
 sky130_fd_sc_hd__nor2_2 _4988_ (.A(_3589_),
    .B(_0156_),
    .Y(_0214_));
 sky130_fd_sc_hd__or2_4 _4989_ (.A(_3539_),
    .B(_0156_),
    .X(_0215_));
 sky130_fd_sc_hd__xor2_4 _4990_ (.A(_0181_),
    .B(_0214_),
    .X(_0216_));
 sky130_fd_sc_hd__nand2_4 _4991_ (.A(net117),
    .B(net60),
    .Y(_0217_));
 sky130_fd_sc_hd__xnor2_4 _4992_ (.A(_0216_),
    .B(_0217_),
    .Y(_0218_));
 sky130_fd_sc_hd__xor2_4 _4993_ (.A(_0211_),
    .B(_0212_),
    .X(_0219_));
 sky130_fd_sc_hd__o21ai_4 _4994_ (.A1(_0218_),
    .A2(_0219_),
    .B1(_0213_),
    .Y(_0220_));
 sky130_fd_sc_hd__xor2_4 _4995_ (.A(_0185_),
    .B(_0186_),
    .X(_0221_));
 sky130_fd_sc_hd__nand2_1 _4996_ (.A(_0220_),
    .B(_0221_),
    .Y(_0222_));
 sky130_fd_sc_hd__o22ai_4 _4997_ (.A1(_0180_),
    .A2(_0215_),
    .B1(_0216_),
    .B2(_0217_),
    .Y(_0223_));
 sky130_fd_sc_hd__and3_4 _4998_ (.A(net120),
    .B(net60),
    .C(_0223_),
    .X(_0224_));
 sky130_fd_sc_hd__a21oi_2 _4999_ (.A1(net120),
    .A2(net60),
    .B1(_0223_),
    .Y(_0225_));
 sky130_fd_sc_hd__nor2_4 _5000_ (.A(_0224_),
    .B(_0225_),
    .Y(_0226_));
 sky130_fd_sc_hd__xor2_4 _5001_ (.A(_0220_),
    .B(_0221_),
    .X(_0227_));
 sky130_fd_sc_hd__a21boi_4 _5002_ (.A1(_0226_),
    .A2(_0227_),
    .B1_N(_0222_),
    .Y(_0228_));
 sky130_fd_sc_hd__xnor2_4 _5003_ (.A(_0191_),
    .B(_0195_),
    .Y(_0229_));
 sky130_fd_sc_hd__nor2_1 _5004_ (.A(_0228_),
    .B(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__xor2_4 _5005_ (.A(_0228_),
    .B(_0229_),
    .X(_0231_));
 sky130_fd_sc_hd__a21oi_4 _5006_ (.A1(_0224_),
    .A2(_0231_),
    .B1(_0230_),
    .Y(_0232_));
 sky130_fd_sc_hd__or2_1 _5007_ (.A(_0206_),
    .B(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__xnor2_4 _5008_ (.A(_0206_),
    .B(_0232_),
    .Y(_0234_));
 sky130_fd_sc_hd__xnor2_1 _5009_ (.A(_0224_),
    .B(_0231_),
    .Y(_0235_));
 sky130_fd_sc_hd__xnor2_4 _5010_ (.A(_0226_),
    .B(_0227_),
    .Y(_0236_));
 sky130_fd_sc_hd__xor2_4 _5011_ (.A(_0218_),
    .B(_0219_),
    .X(_0237_));
 sky130_fd_sc_hd__a21o_1 _5012_ (.A1(_0207_),
    .A2(_0209_),
    .B1(_0208_),
    .X(_0238_));
 sky130_fd_sc_hd__or4b_2 _5013_ (.A(net95),
    .B(net68),
    .C(net56),
    .D_N(net55),
    .X(_0239_));
 sky130_fd_sc_hd__nor2_1 _5014_ (.A(net93),
    .B(_0156_),
    .Y(_0240_));
 sky130_fd_sc_hd__a2bb2o_1 _5015_ (.A1_N(net68),
    .A2_N(net56),
    .B1(net55),
    .B2(_3582_),
    .X(_0241_));
 sky130_fd_sc_hd__and3_1 _5016_ (.A(_0239_),
    .B(_0240_),
    .C(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__a21bo_1 _5017_ (.A1(_0240_),
    .A2(_0241_),
    .B1_N(_0239_),
    .X(_0243_));
 sky130_fd_sc_hd__and3_2 _5018_ (.A(_0210_),
    .B(_0238_),
    .C(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__and2_1 _5019_ (.A(net115),
    .B(net60),
    .X(_0245_));
 sky130_fd_sc_hd__nand2_4 _5020_ (.A(_3590_),
    .B(net60),
    .Y(_0246_));
 sky130_fd_sc_hd__nor2_4 _5021_ (.A(_0215_),
    .B(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__xor2_4 _5022_ (.A(_0215_),
    .B(_0246_),
    .X(_0248_));
 sky130_fd_sc_hd__a21o_1 _5023_ (.A1(_0210_),
    .A2(_0238_),
    .B1(_0243_),
    .X(_0249_));
 sky130_fd_sc_hd__and2b_1 _5024_ (.A_N(_0244_),
    .B(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__a21oi_4 _5025_ (.A1(_0248_),
    .A2(_0249_),
    .B1(_0244_),
    .Y(_0251_));
 sky130_fd_sc_hd__and2b_1 _5026_ (.A_N(_0251_),
    .B(_0237_),
    .X(_0252_));
 sky130_fd_sc_hd__xnor2_4 _5027_ (.A(_0237_),
    .B(_0251_),
    .Y(_0253_));
 sky130_fd_sc_hd__a21oi_4 _5028_ (.A1(_0247_),
    .A2(_0253_),
    .B1(_0252_),
    .Y(_0254_));
 sky130_fd_sc_hd__or2_1 _5029_ (.A(_0236_),
    .B(_0254_),
    .X(_0255_));
 sky130_fd_sc_hd__xnor2_4 _5030_ (.A(_0236_),
    .B(_0254_),
    .Y(_0256_));
 sky130_fd_sc_hd__a21oi_1 _5031_ (.A1(_0239_),
    .A2(_0241_),
    .B1(_0240_),
    .Y(_0257_));
 sky130_fd_sc_hd__nor2_1 _5032_ (.A(_0242_),
    .B(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hd__nor2_1 _5033_ (.A(net96),
    .B(_0156_),
    .Y(_0259_));
 sky130_fd_sc_hd__and3_1 _5034_ (.A(_3647_),
    .B(_0123_),
    .C(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__a21o_1 _5035_ (.A1(_3647_),
    .A2(_0123_),
    .B1(_0259_),
    .X(_0261_));
 sky130_fd_sc_hd__a31o_1 _5036_ (.A1(net92),
    .A2(_3997_),
    .A3(_0261_),
    .B1(_0260_),
    .X(_0262_));
 sky130_fd_sc_hd__nand2_1 _5037_ (.A(_0258_),
    .B(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__xor2_1 _5038_ (.A(_0258_),
    .B(_0262_),
    .X(_0264_));
 sky130_fd_sc_hd__nand2_1 _5039_ (.A(_0245_),
    .B(_0264_),
    .Y(_0265_));
 sky130_fd_sc_hd__nor2_1 _5040_ (.A(net92),
    .B(_0123_),
    .Y(_0266_));
 sky130_fd_sc_hd__o2111a_1 _5041_ (.A1(_0208_),
    .A2(_0266_),
    .B1(_0259_),
    .C1(_3647_),
    .D1(_3997_),
    .X(_0267_));
 sky130_fd_sc_hd__o21ai_1 _5042_ (.A1(_0245_),
    .A2(_0264_),
    .B1(_0267_),
    .Y(_0268_));
 sky130_fd_sc_hd__xnor2_1 _5043_ (.A(_0248_),
    .B(_0250_),
    .Y(_0269_));
 sky130_fd_sc_hd__o21a_1 _5044_ (.A1(_0263_),
    .A2(_0268_),
    .B1(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__a31o_2 _5045_ (.A1(_0263_),
    .A2(_0265_),
    .A3(_0268_),
    .B1(_0270_),
    .X(_0271_));
 sky130_fd_sc_hd__xnor2_4 _5046_ (.A(_0247_),
    .B(_0253_),
    .Y(_0272_));
 sky130_fd_sc_hd__or3_4 _5047_ (.A(_0256_),
    .B(_0271_),
    .C(_0272_),
    .X(_0273_));
 sky130_fd_sc_hd__a21o_2 _5048_ (.A1(_0255_),
    .A2(_0273_),
    .B1(_0235_),
    .X(_0274_));
 sky130_fd_sc_hd__or2_4 _5049_ (.A(_0234_),
    .B(_0274_),
    .X(_0275_));
 sky130_fd_sc_hd__or2_1 _5050_ (.A(_0203_),
    .B(_0205_),
    .X(_0276_));
 sky130_fd_sc_hd__a21oi_1 _5051_ (.A1(_0233_),
    .A2(_0275_),
    .B1(_0276_),
    .Y(_0277_));
 sky130_fd_sc_hd__o211a_2 _5052_ (.A1(_0234_),
    .A2(_0274_),
    .B1(_0204_),
    .C1(_0233_),
    .X(_0278_));
 sky130_fd_sc_hd__or3_1 _5053_ (.A(_0171_),
    .B(_0205_),
    .C(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__or4_4 _5054_ (.A(_0141_),
    .B(_0171_),
    .C(_0205_),
    .D(_0278_),
    .X(_0280_));
 sky130_fd_sc_hd__a21o_2 _5055_ (.A1(_0139_),
    .A2(_0170_),
    .B1(_0140_),
    .X(_0281_));
 sky130_fd_sc_hd__a21oi_4 _5056_ (.A1(_0280_),
    .A2(_0281_),
    .B1(_0114_),
    .Y(_0282_));
 sky130_fd_sc_hd__a211o_1 _5057_ (.A1(_0280_),
    .A2(_0281_),
    .B1(_0089_),
    .C1(_0114_),
    .X(_0283_));
 sky130_fd_sc_hd__or2_1 _5058_ (.A(_0089_),
    .B(_0114_),
    .X(_0284_));
 sky130_fd_sc_hd__a211o_2 _5059_ (.A1(_0280_),
    .A2(_0281_),
    .B1(_0284_),
    .C1(_3986_),
    .X(_0285_));
 sky130_fd_sc_hd__o21bai_4 _5060_ (.A1(_0088_),
    .A2(_0112_),
    .B1_N(_0086_),
    .Y(_0286_));
 sky130_fd_sc_hd__o221a_2 _5061_ (.A1(_3968_),
    .A2(_3983_),
    .B1(_3986_),
    .B2(_0286_),
    .C1(_3967_),
    .X(_0287_));
 sky130_fd_sc_hd__nand2_4 _5062_ (.A(_0285_),
    .B(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__xnor2_4 _5063_ (.A(_3942_),
    .B(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hd__or2_4 _5064_ (.A(net69),
    .B(net47),
    .X(_0290_));
 sky130_fd_sc_hd__a21oi_4 _5065_ (.A1(_1935_),
    .A2(_1946_),
    .B1(net169),
    .Y(_0291_));
 sky130_fd_sc_hd__nor2_2 _5066_ (.A(_1715_),
    .B(_2045_),
    .Y(_0292_));
 sky130_fd_sc_hd__o2111a_2 _5067_ (.A1(\posit_add.in1[0] ),
    .A2(_1891_),
    .B1(_1957_),
    .C1(net167),
    .D1(net131),
    .X(_0293_));
 sky130_fd_sc_hd__nand2_2 _5068_ (.A(net173),
    .B(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hd__o31a_4 _5069_ (.A1(net172),
    .A2(_0291_),
    .A3(_0292_),
    .B1(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__o31ai_4 _5070_ (.A1(net172),
    .A2(_0291_),
    .A3(_0292_),
    .B1(_0294_),
    .Y(_0296_));
 sky130_fd_sc_hd__nand2_2 _5071_ (.A(_0283_),
    .B(_0286_),
    .Y(_0297_));
 sky130_fd_sc_hd__a21o_2 _5072_ (.A1(_0283_),
    .A2(_0286_),
    .B1(_3985_),
    .X(_0298_));
 sky130_fd_sc_hd__a21o_4 _5073_ (.A1(_3983_),
    .A2(_0298_),
    .B1(_3969_),
    .X(_0299_));
 sky130_fd_sc_hd__nand3_4 _5074_ (.A(_3969_),
    .B(_3983_),
    .C(_0298_),
    .Y(_0300_));
 sky130_fd_sc_hd__nand2_2 _5075_ (.A(_0299_),
    .B(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__and3_4 _5076_ (.A(net65),
    .B(_0299_),
    .C(_0300_),
    .X(_0302_));
 sky130_fd_sc_hd__nand3_4 _5077_ (.A(_3464_),
    .B(_0299_),
    .C(_0300_),
    .Y(_0303_));
 sky130_fd_sc_hd__nor2_4 _5078_ (.A(net47),
    .B(net67),
    .Y(_0304_));
 sky130_fd_sc_hd__and2b_2 _5079_ (.A_N(_0290_),
    .B(_0302_),
    .X(_0305_));
 sky130_fd_sc_hd__a211o_2 _5080_ (.A1(_1165_),
    .A2(net129),
    .B1(_3453_),
    .C1(net133),
    .X(_0306_));
 sky130_fd_sc_hd__a211o_2 _5081_ (.A1(_1594_),
    .A2(net129),
    .B1(_3448_),
    .C1(net131),
    .X(_0307_));
 sky130_fd_sc_hd__a21o_2 _5082_ (.A1(_0306_),
    .A2(_0307_),
    .B1(_1715_),
    .X(_0308_));
 sky130_fd_sc_hd__a211o_4 _5083_ (.A1(_1671_),
    .A2(net130),
    .B1(_3447_),
    .C1(net133),
    .X(_0309_));
 sky130_fd_sc_hd__a211o_4 _5084_ (.A1(_1517_),
    .A2(net129),
    .B1(_3460_),
    .C1(net131),
    .X(_0310_));
 sky130_fd_sc_hd__a21o_1 _5085_ (.A1(_0309_),
    .A2(_0310_),
    .B1(net167),
    .X(_0311_));
 sky130_fd_sc_hd__o2111a_1 _5086_ (.A1(_1385_),
    .A2(_1869_),
    .B1(_1770_),
    .C1(\posit_add.in1[0] ),
    .D1(_1352_),
    .X(_0312_));
 sky130_fd_sc_hd__and3_2 _5087_ (.A(net172),
    .B(net167),
    .C(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__a31oi_4 _5088_ (.A1(net170),
    .A2(_0308_),
    .A3(_0311_),
    .B1(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__a31o_2 _5089_ (.A1(net170),
    .A2(_0308_),
    .A3(_0311_),
    .B1(_0313_),
    .X(_0315_));
 sky130_fd_sc_hd__and2_1 _5090_ (.A(_3506_),
    .B(_3894_),
    .X(_0316_));
 sky130_fd_sc_hd__a21o_1 _5091_ (.A1(net117),
    .A2(net59),
    .B1(_0316_),
    .X(_0317_));
 sky130_fd_sc_hd__inv_2 _5092_ (.A(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__xnor2_1 _5093_ (.A(_3915_),
    .B(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__a21o_1 _5094_ (.A1(_3895_),
    .A2(_0319_),
    .B1(_3907_),
    .X(_0320_));
 sky130_fd_sc_hd__and3_1 _5095_ (.A(_3917_),
    .B(_3920_),
    .C(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__a21oi_2 _5096_ (.A1(_3917_),
    .A2(_3920_),
    .B1(_0320_),
    .Y(_0322_));
 sky130_fd_sc_hd__inv_2 _5097_ (.A(_0322_),
    .Y(_0323_));
 sky130_fd_sc_hd__or2_4 _5098_ (.A(_0321_),
    .B(_0322_),
    .X(_0324_));
 sky130_fd_sc_hd__a21bo_2 _5099_ (.A1(_3942_),
    .A2(_0288_),
    .B1_N(_3939_),
    .X(_0325_));
 sky130_fd_sc_hd__xor2_4 _5100_ (.A(_0324_),
    .B(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__inv_2 _5101_ (.A(net43),
    .Y(_0327_));
 sky130_fd_sc_hd__or2_4 _5102_ (.A(net90),
    .B(net43),
    .X(_0328_));
 sky130_fd_sc_hd__xnor2_4 _5103_ (.A(_0303_),
    .B(_0304_),
    .Y(_0329_));
 sky130_fd_sc_hd__and3_2 _5104_ (.A(net87),
    .B(_0327_),
    .C(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__or2_4 _5105_ (.A(net67),
    .B(_0326_),
    .X(_0331_));
 sky130_fd_sc_hd__nor3_2 _5106_ (.A(\posit_add.in1[14] ),
    .B(_1044_),
    .C(_1055_),
    .Y(_0332_));
 sky130_fd_sc_hd__or3_4 _5107_ (.A(\posit_add.in1[14] ),
    .B(_1044_),
    .C(_1055_),
    .X(_0333_));
 sky130_fd_sc_hd__or2_1 _5108_ (.A(net47),
    .B(net200),
    .X(_0334_));
 sky130_fd_sc_hd__or2_4 _5109_ (.A(_0301_),
    .B(net200),
    .X(_0335_));
 sky130_fd_sc_hd__or2_1 _5110_ (.A(_0303_),
    .B(_0334_),
    .X(_0336_));
 sky130_fd_sc_hd__xnor2_4 _5111_ (.A(_0290_),
    .B(_0335_),
    .Y(_0337_));
 sky130_fd_sc_hd__or2_1 _5112_ (.A(_0331_),
    .B(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__xor2_4 _5113_ (.A(_0331_),
    .B(_0337_),
    .X(_0339_));
 sky130_fd_sc_hd__o21a_1 _5114_ (.A1(_0305_),
    .A2(_0330_),
    .B1(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__o21ai_4 _5115_ (.A1(_0305_),
    .A2(_0330_),
    .B1(_0339_),
    .Y(_0341_));
 sky130_fd_sc_hd__a21o_1 _5116_ (.A1(_3939_),
    .A2(_0323_),
    .B1(_0321_),
    .X(_0342_));
 sky130_fd_sc_hd__a211o_2 _5117_ (.A1(_0285_),
    .A2(_0287_),
    .B1(_0324_),
    .C1(_3941_),
    .X(_0343_));
 sky130_fd_sc_hd__a21o_1 _5118_ (.A1(net120),
    .A2(net59),
    .B1(_0316_),
    .X(_0344_));
 sky130_fd_sc_hd__o211a_1 _5119_ (.A1(_3915_),
    .A2(_0318_),
    .B1(_0344_),
    .C1(_3906_),
    .X(_0345_));
 sky130_fd_sc_hd__a21o_2 _5120_ (.A1(net120),
    .A2(_3907_),
    .B1(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__and3_2 _5121_ (.A(_0342_),
    .B(_0343_),
    .C(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__a21oi_4 _5122_ (.A1(_0342_),
    .A2(_0343_),
    .B1(_0346_),
    .Y(_0348_));
 sky130_fd_sc_hd__nor2_4 _5123_ (.A(_0347_),
    .B(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__nor2_1 _5124_ (.A(net89),
    .B(net42),
    .Y(_0350_));
 sky130_fd_sc_hd__or2_1 _5125_ (.A(net90),
    .B(net42),
    .X(_0351_));
 sky130_fd_sc_hd__nor2_2 _5126_ (.A(net212),
    .B(net67),
    .Y(_0352_));
 sky130_fd_sc_hd__or2_4 _5127_ (.A(net213),
    .B(net67),
    .X(_0353_));
 sky130_fd_sc_hd__nor2_1 _5128_ (.A(net212),
    .B(net90),
    .Y(_0354_));
 sky130_fd_sc_hd__or2_4 _5129_ (.A(net213),
    .B(net90),
    .X(_0355_));
 sky130_fd_sc_hd__nor2_2 _5130_ (.A(_0295_),
    .B(_0349_),
    .Y(_0356_));
 sky130_fd_sc_hd__a211o_2 _5131_ (.A1(_1561_),
    .A2(net130),
    .B1(_2023_),
    .C1(net133),
    .X(_0357_));
 sky130_fd_sc_hd__a211o_2 _5132_ (.A1(_1638_),
    .A2(net130),
    .B1(_1924_),
    .C1(net132),
    .X(_0358_));
 sky130_fd_sc_hd__nand2_2 _5133_ (.A(_0357_),
    .B(_0358_),
    .Y(_0359_));
 sky130_fd_sc_hd__a211o_4 _5134_ (.A1(_1484_),
    .A2(net130),
    .B1(_1913_),
    .C1(_1781_),
    .X(_0360_));
 sky130_fd_sc_hd__a211o_4 _5135_ (.A1(net235),
    .A2(net130),
    .B1(_1968_),
    .C1(net131),
    .X(_0361_));
 sky130_fd_sc_hd__a21oi_4 _5136_ (.A1(_0360_),
    .A2(_0361_),
    .B1(net168),
    .Y(_0362_));
 sky130_fd_sc_hd__a211o_4 _5137_ (.A1(net168),
    .A2(_0359_),
    .B1(_0362_),
    .C1(net173),
    .X(_0363_));
 sky130_fd_sc_hd__clkinv_4 _5138_ (.A(net86),
    .Y(_0364_));
 sky130_fd_sc_hd__or2_4 _5139_ (.A(net42),
    .B(net85),
    .X(_0365_));
 sky130_fd_sc_hd__nor2_2 _5140_ (.A(net212),
    .B(net85),
    .Y(_0366_));
 sky130_fd_sc_hd__or2_1 _5141_ (.A(net213),
    .B(net86),
    .X(_0367_));
 sky130_fd_sc_hd__and3_1 _5142_ (.A(_0350_),
    .B(_0353_),
    .C(_0366_),
    .X(_0368_));
 sky130_fd_sc_hd__a21o_1 _5143_ (.A1(_0354_),
    .A2(_0365_),
    .B1(_0356_),
    .X(_0369_));
 sky130_fd_sc_hd__o31a_2 _5144_ (.A1(_0351_),
    .A2(_0353_),
    .A3(_0366_),
    .B1(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__and3_4 _5145_ (.A(_1715_),
    .B(_3458_),
    .C(_3461_),
    .X(_0371_));
 sky130_fd_sc_hd__a211oi_4 _5146_ (.A1(net167),
    .A2(_3451_),
    .B1(_0371_),
    .C1(net172),
    .Y(_0372_));
 sky130_fd_sc_hd__a211o_4 _5147_ (.A1(net167),
    .A2(_3451_),
    .B1(_0371_),
    .C1(net172),
    .X(_0373_));
 sky130_fd_sc_hd__or2_2 _5148_ (.A(net42),
    .B(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__nor2_4 _5149_ (.A(net213),
    .B(net82),
    .Y(_0375_));
 sky130_fd_sc_hd__or2_2 _5150_ (.A(net212),
    .B(_0373_),
    .X(_0376_));
 sky130_fd_sc_hd__and3b_2 _5151_ (.A_N(_0365_),
    .B(_0375_),
    .C(_0355_),
    .X(_0377_));
 sky130_fd_sc_hd__xnor2_2 _5152_ (.A(_0341_),
    .B(_0370_),
    .Y(_0378_));
 sky130_fd_sc_hd__a22o_1 _5153_ (.A1(_0340_),
    .A2(_0370_),
    .B1(_0377_),
    .B2(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__xor2_2 _5154_ (.A(_0377_),
    .B(_0378_),
    .X(_0380_));
 sky130_fd_sc_hd__nand2_1 _5155_ (.A(_0336_),
    .B(_0338_),
    .Y(_0381_));
 sky130_fd_sc_hd__or3_4 _5156_ (.A(net69),
    .B(_0326_),
    .C(_0334_),
    .X(_0382_));
 sky130_fd_sc_hd__o21ai_1 _5157_ (.A1(net69),
    .A2(_0326_),
    .B1(_0334_),
    .Y(_0383_));
 sky130_fd_sc_hd__and2_1 _5158_ (.A(_0382_),
    .B(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__a21bo_1 _5159_ (.A1(_0336_),
    .A2(_0338_),
    .B1_N(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__or2_1 _5160_ (.A(_0381_),
    .B(_0384_),
    .X(_0386_));
 sky130_fd_sc_hd__and2_1 _5161_ (.A(_0385_),
    .B(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__nand2_2 _5162_ (.A(_0380_),
    .B(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__or2_4 _5163_ (.A(net70),
    .B(net42),
    .X(_0389_));
 sky130_fd_sc_hd__or2_1 _5164_ (.A(net69),
    .B(net213),
    .X(_0390_));
 sky130_fd_sc_hd__and3b_1 _5165_ (.A_N(_0389_),
    .B(_0351_),
    .C(_0352_),
    .X(_0391_));
 sky130_fd_sc_hd__and3_1 _5166_ (.A(net70),
    .B(_0350_),
    .C(_0352_),
    .X(_0392_));
 sky130_fd_sc_hd__a211o_1 _5167_ (.A1(_0353_),
    .A2(_0389_),
    .B1(_0391_),
    .C1(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__nor2_2 _5168_ (.A(_0385_),
    .B(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__and2_1 _5169_ (.A(_0385_),
    .B(_0393_),
    .X(_0395_));
 sky130_fd_sc_hd__nor2_1 _5170_ (.A(_0394_),
    .B(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__and2_1 _5171_ (.A(_0368_),
    .B(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__nor2_1 _5172_ (.A(_0368_),
    .B(_0396_),
    .Y(_0398_));
 sky130_fd_sc_hd__or2_2 _5173_ (.A(_0397_),
    .B(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__and3_2 _5174_ (.A(_0290_),
    .B(_0327_),
    .C(net199),
    .X(_0400_));
 sky130_fd_sc_hd__or3b_2 _5175_ (.A(_0397_),
    .B(_0398_),
    .C_N(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__xnor2_2 _5176_ (.A(_0399_),
    .B(_0400_),
    .Y(_0402_));
 sky130_fd_sc_hd__and3_1 _5177_ (.A(_0380_),
    .B(_0387_),
    .C(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__xnor2_2 _5178_ (.A(_0388_),
    .B(_0402_),
    .Y(_0404_));
 sky130_fd_sc_hd__xnor2_1 _5179_ (.A(_0379_),
    .B(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__or2_2 _5180_ (.A(_0380_),
    .B(_0387_),
    .X(_0406_));
 sky130_fd_sc_hd__nand2_4 _5181_ (.A(_0388_),
    .B(_0406_),
    .Y(_0407_));
 sky130_fd_sc_hd__or3_2 _5182_ (.A(_0305_),
    .B(_0330_),
    .C(_0339_),
    .X(_0408_));
 sky130_fd_sc_hd__nand2_4 _5183_ (.A(_0341_),
    .B(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__xor2_4 _5184_ (.A(_3985_),
    .B(_0297_),
    .X(_0410_));
 sky130_fd_sc_hd__inv_2 _5185_ (.A(net46),
    .Y(_0411_));
 sky130_fd_sc_hd__nor2_4 _5186_ (.A(net200),
    .B(_0410_),
    .Y(_0412_));
 sky130_fd_sc_hd__xnor2_4 _5187_ (.A(_0328_),
    .B(_0329_),
    .Y(_0413_));
 sky130_fd_sc_hd__o21ai_4 _5188_ (.A1(_0112_),
    .A2(_0282_),
    .B1(_0090_),
    .Y(_0414_));
 sky130_fd_sc_hd__or3_4 _5189_ (.A(_0090_),
    .B(_0112_),
    .C(_0282_),
    .X(_0415_));
 sky130_fd_sc_hd__nand2_4 _5190_ (.A(_0414_),
    .B(_0415_),
    .Y(_0416_));
 sky130_fd_sc_hd__or2_1 _5191_ (.A(net70),
    .B(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__or2_4 _5192_ (.A(net200),
    .B(_0416_),
    .X(_0418_));
 sky130_fd_sc_hd__nor2_4 _5193_ (.A(net69),
    .B(net46),
    .Y(_0419_));
 sky130_fd_sc_hd__and2b_4 _5194_ (.A_N(_0418_),
    .B(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__nand2_1 _5195_ (.A(_0413_),
    .B(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__xnor2_4 _5196_ (.A(_0413_),
    .B(_0420_),
    .Y(_0422_));
 sky130_fd_sc_hd__and3_4 _5197_ (.A(_0299_),
    .B(_0300_),
    .C(net87),
    .X(_0423_));
 sky130_fd_sc_hd__or2_4 _5198_ (.A(net47),
    .B(net90),
    .X(_0424_));
 sky130_fd_sc_hd__nor2_4 _5199_ (.A(net43),
    .B(net85),
    .Y(_0425_));
 sky130_fd_sc_hd__xnor2_4 _5200_ (.A(_0302_),
    .B(_0424_),
    .Y(_0426_));
 sky130_fd_sc_hd__a22oi_4 _5201_ (.A1(_0304_),
    .A2(_0423_),
    .B1(_0425_),
    .B2(_0426_),
    .Y(_0427_));
 sky130_fd_sc_hd__xor2_4 _5202_ (.A(_0422_),
    .B(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__nand2_4 _5203_ (.A(_0412_),
    .B(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__and2_4 _5204_ (.A(net170),
    .B(_1990_),
    .X(_0430_));
 sky130_fd_sc_hd__nand2_8 _5205_ (.A(net170),
    .B(_1990_),
    .Y(_0431_));
 sky130_fd_sc_hd__nor2_2 _5206_ (.A(net42),
    .B(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__or2_4 _5207_ (.A(net211),
    .B(_0431_),
    .X(_0433_));
 sky130_fd_sc_hd__or3_4 _5208_ (.A(_0366_),
    .B(_0374_),
    .C(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__o21ai_4 _5209_ (.A1(_0422_),
    .A2(_0427_),
    .B1(_0421_),
    .Y(_0435_));
 sky130_fd_sc_hd__a21o_1 _5210_ (.A1(_0366_),
    .A2(_0374_),
    .B1(_0350_),
    .X(_0436_));
 sky130_fd_sc_hd__o31a_4 _5211_ (.A1(_0355_),
    .A2(_0365_),
    .A3(_0375_),
    .B1(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__xor2_4 _5212_ (.A(_0435_),
    .B(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__and2b_1 _5213_ (.A_N(_0434_),
    .B(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__xnor2_4 _5214_ (.A(_0434_),
    .B(_0438_),
    .Y(_0440_));
 sky130_fd_sc_hd__xor2_4 _5215_ (.A(_0409_),
    .B(_0429_),
    .X(_0441_));
 sky130_fd_sc_hd__nand2_1 _5216_ (.A(_0440_),
    .B(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__o21a_2 _5217_ (.A1(_0409_),
    .A2(_0429_),
    .B1(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__nor2_1 _5218_ (.A(_0407_),
    .B(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__a21o_2 _5219_ (.A1(_0435_),
    .A2(_0437_),
    .B1(_0439_),
    .X(_0445_));
 sky130_fd_sc_hd__xor2_4 _5220_ (.A(_0407_),
    .B(_0443_),
    .X(_0446_));
 sky130_fd_sc_hd__a21oi_1 _5221_ (.A1(_0445_),
    .A2(_0446_),
    .B1(_0444_),
    .Y(_0447_));
 sky130_fd_sc_hd__or2_4 _5222_ (.A(_0405_),
    .B(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__o21ai_2 _5223_ (.A1(net201),
    .A2(net42),
    .B1(_0390_),
    .Y(_0449_));
 sky130_fd_sc_hd__o21ai_4 _5224_ (.A1(_0352_),
    .A2(_0389_),
    .B1(_0449_),
    .Y(_0450_));
 sky130_fd_sc_hd__o21bai_4 _5225_ (.A1(_0382_),
    .A2(_0450_),
    .B1_N(_0392_),
    .Y(_0451_));
 sky130_fd_sc_hd__inv_2 _5226_ (.A(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__and2_1 _5227_ (.A(_0382_),
    .B(_0450_),
    .X(_0453_));
 sky130_fd_sc_hd__nor2_1 _5228_ (.A(_0451_),
    .B(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__or3_1 _5229_ (.A(_0401_),
    .B(_0451_),
    .C(_0453_),
    .X(_0455_));
 sky130_fd_sc_hd__xnor2_1 _5230_ (.A(_0401_),
    .B(_0454_),
    .Y(_0456_));
 sky130_fd_sc_hd__o21ai_2 _5231_ (.A1(_0394_),
    .A2(_0397_),
    .B1(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__or3_1 _5232_ (.A(_0394_),
    .B(_0397_),
    .C(_0456_),
    .X(_0458_));
 sky130_fd_sc_hd__nand2_1 _5233_ (.A(_0457_),
    .B(_0458_),
    .Y(_0459_));
 sky130_fd_sc_hd__a21oi_1 _5234_ (.A1(_0379_),
    .A2(_0404_),
    .B1(_0403_),
    .Y(_0460_));
 sky130_fd_sc_hd__or2_2 _5235_ (.A(_0459_),
    .B(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__nand2_1 _5236_ (.A(_0459_),
    .B(_0460_),
    .Y(_0462_));
 sky130_fd_sc_hd__and2_2 _5237_ (.A(_0461_),
    .B(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__xor2_4 _5238_ (.A(_0448_),
    .B(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__xnor2_4 _5239_ (.A(_0445_),
    .B(_0446_),
    .Y(_0465_));
 sky130_fd_sc_hd__xnor2_2 _5240_ (.A(_0440_),
    .B(_0441_),
    .Y(_0466_));
 sky130_fd_sc_hd__xnor2_4 _5241_ (.A(_0412_),
    .B(_0428_),
    .Y(_0467_));
 sky130_fd_sc_hd__and3_4 _5242_ (.A(_0299_),
    .B(_0300_),
    .C(_0364_),
    .X(_0468_));
 sky130_fd_sc_hd__nor2_4 _5243_ (.A(_0289_),
    .B(net86),
    .Y(_0469_));
 sky130_fd_sc_hd__nor2_4 _5244_ (.A(_0326_),
    .B(net82),
    .Y(_0470_));
 sky130_fd_sc_hd__xor2_4 _5245_ (.A(_0423_),
    .B(_0469_),
    .X(_0471_));
 sky130_fd_sc_hd__a22o_4 _5246_ (.A1(_0423_),
    .A2(_0469_),
    .B1(_0470_),
    .B2(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__and3_2 _5247_ (.A(_0114_),
    .B(_0280_),
    .C(_0281_),
    .X(_0473_));
 sky130_fd_sc_hd__nor2_8 _5248_ (.A(_0282_),
    .B(_0473_),
    .Y(_0474_));
 sky130_fd_sc_hd__nand2_4 _5249_ (.A(_3464_),
    .B(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__nor2_1 _5250_ (.A(_0418_),
    .B(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__or2_2 _5251_ (.A(net66),
    .B(_0410_),
    .X(_0477_));
 sky130_fd_sc_hd__a32o_1 _5252_ (.A1(_3464_),
    .A2(_0414_),
    .A3(_0415_),
    .B1(net48),
    .B2(net199),
    .X(_0478_));
 sky130_fd_sc_hd__o21a_2 _5253_ (.A1(_0418_),
    .A2(_0475_),
    .B1(_0478_),
    .X(_0479_));
 sky130_fd_sc_hd__a31o_4 _5254_ (.A1(net65),
    .A2(_0411_),
    .A3(_0479_),
    .B1(_0476_),
    .X(_0480_));
 sky130_fd_sc_hd__xor2_4 _5255_ (.A(_0425_),
    .B(_0426_),
    .X(_0481_));
 sky130_fd_sc_hd__nand2_1 _5256_ (.A(_0480_),
    .B(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__xor2_4 _5257_ (.A(_0480_),
    .B(_0481_),
    .X(_0483_));
 sky130_fd_sc_hd__xor2_4 _5258_ (.A(_0472_),
    .B(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__xnor2_4 _5259_ (.A(_0418_),
    .B(_0419_),
    .Y(_0485_));
 sky130_fd_sc_hd__and2_2 _5260_ (.A(_0484_),
    .B(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__and2b_1 _5261_ (.A_N(_0467_),
    .B(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__xnor2_4 _5262_ (.A(_0467_),
    .B(_0486_),
    .Y(_0488_));
 sky130_fd_sc_hd__a21boi_4 _5263_ (.A1(_0472_),
    .A2(_0483_),
    .B1_N(_0482_),
    .Y(_0489_));
 sky130_fd_sc_hd__or3_1 _5264_ (.A(_0365_),
    .B(_0376_),
    .C(_0432_),
    .X(_0490_));
 sky130_fd_sc_hd__nand2_1 _5265_ (.A(_0434_),
    .B(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__a21o_2 _5266_ (.A1(_0365_),
    .A2(_0376_),
    .B1(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__xor2_4 _5267_ (.A(_0489_),
    .B(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__and2_2 _5268_ (.A(_1715_),
    .B(_0312_),
    .X(_0494_));
 sky130_fd_sc_hd__a31oi_4 _5269_ (.A1(net167),
    .A2(_0309_),
    .A3(_0310_),
    .B1(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__a31o_4 _5270_ (.A1(net167),
    .A2(_0309_),
    .A3(_0310_),
    .B1(_0494_),
    .X(_0496_));
 sky130_fd_sc_hd__nor2_1 _5271_ (.A(net173),
    .B(_0495_),
    .Y(_0497_));
 sky130_fd_sc_hd__nand2_8 _5272_ (.A(net171),
    .B(_0496_),
    .Y(_0498_));
 sky130_fd_sc_hd__or2_4 _5273_ (.A(net42),
    .B(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__nor2_4 _5274_ (.A(net211),
    .B(net75),
    .Y(_0500_));
 sky130_fd_sc_hd__and3_4 _5275_ (.A(_0376_),
    .B(_0432_),
    .C(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__xor2_4 _5276_ (.A(_0493_),
    .B(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__a21oi_2 _5277_ (.A1(_0488_),
    .A2(_0502_),
    .B1(_0487_),
    .Y(_0503_));
 sky130_fd_sc_hd__nor2_2 _5278_ (.A(_0466_),
    .B(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__a2bb2o_4 _5279_ (.A1_N(_0489_),
    .A2_N(_0492_),
    .B1(_0493_),
    .B2(_0501_),
    .X(_0505_));
 sky130_fd_sc_hd__nand2_2 _5280_ (.A(_0466_),
    .B(_0503_),
    .Y(_0506_));
 sky130_fd_sc_hd__and2b_2 _5281_ (.A_N(_0504_),
    .B(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__a21oi_4 _5282_ (.A1(_0505_),
    .A2(_0506_),
    .B1(_0504_),
    .Y(_0508_));
 sky130_fd_sc_hd__nor2_1 _5283_ (.A(_0465_),
    .B(_0508_),
    .Y(_0509_));
 sky130_fd_sc_hd__nand2_1 _5284_ (.A(_0405_),
    .B(_0447_),
    .Y(_0510_));
 sky130_fd_sc_hd__and2_1 _5285_ (.A(_0448_),
    .B(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__nand2_1 _5286_ (.A(_0509_),
    .B(_0511_),
    .Y(_0512_));
 sky130_fd_sc_hd__or2_1 _5287_ (.A(_0509_),
    .B(_0511_),
    .X(_0513_));
 sky130_fd_sc_hd__nand2_1 _5288_ (.A(_0512_),
    .B(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__o31a_2 _5289_ (.A1(_0171_),
    .A2(_0205_),
    .A3(_0278_),
    .B1(_0170_),
    .X(_0515_));
 sky130_fd_sc_hd__xnor2_4 _5290_ (.A(_0141_),
    .B(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__nor2_8 _5291_ (.A(net66),
    .B(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__or2_4 _5292_ (.A(net85),
    .B(_0416_),
    .X(_0518_));
 sky130_fd_sc_hd__nand2_8 _5293_ (.A(net87),
    .B(_0474_),
    .Y(_0519_));
 sky130_fd_sc_hd__xor2_4 _5294_ (.A(_0518_),
    .B(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__nor2_4 _5295_ (.A(net81),
    .B(net46),
    .Y(_0521_));
 sky130_fd_sc_hd__xor2_4 _5296_ (.A(_0520_),
    .B(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__nand2_2 _5297_ (.A(_0517_),
    .B(_0522_),
    .Y(_0523_));
 sky130_fd_sc_hd__xnor2_4 _5298_ (.A(_0517_),
    .B(_0522_),
    .Y(_0524_));
 sky130_fd_sc_hd__and2_1 _5299_ (.A(_0235_),
    .B(_0273_),
    .X(_0525_));
 sky130_fd_sc_hd__a21bo_2 _5300_ (.A1(_0255_),
    .A2(_0525_),
    .B1_N(_0274_),
    .X(_0526_));
 sky130_fd_sc_hd__nor2_4 _5301_ (.A(net84),
    .B(net54),
    .Y(_0527_));
 sky130_fd_sc_hd__nor2_8 _5302_ (.A(net202),
    .B(_0516_),
    .Y(_0528_));
 sky130_fd_sc_hd__nor2_4 _5303_ (.A(net202),
    .B(net54),
    .Y(_0529_));
 sky130_fd_sc_hd__nand2_2 _5304_ (.A(_0527_),
    .B(_0528_),
    .Y(_0530_));
 sky130_fd_sc_hd__nor2_1 _5305_ (.A(net89),
    .B(net53),
    .Y(_0531_));
 sky130_fd_sc_hd__mux2_8 _5306_ (.A0(net89),
    .A1(_0531_),
    .S(_0530_),
    .X(_0532_));
 sky130_fd_sc_hd__o2bb2a_2 _5307_ (.A1_N(_0364_),
    .A2_N(net48),
    .B1(_0416_),
    .B2(net81),
    .X(_0533_));
 sky130_fd_sc_hd__nand2_8 _5308_ (.A(_0372_),
    .B(net48),
    .Y(_0534_));
 sky130_fd_sc_hd__o21ba_2 _5309_ (.A1(_0518_),
    .A2(_0534_),
    .B1_N(_0533_),
    .X(_0535_));
 sky130_fd_sc_hd__or2_4 _5310_ (.A(net46),
    .B(net78),
    .X(_0536_));
 sky130_fd_sc_hd__xnor2_4 _5311_ (.A(_0535_),
    .B(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__o2bb2a_4 _5312_ (.A1_N(_0532_),
    .A2_N(_0537_),
    .B1(net89),
    .B2(_0530_),
    .X(_0538_));
 sky130_fd_sc_hd__nor2_1 _5313_ (.A(_0524_),
    .B(_0538_),
    .Y(_0539_));
 sky130_fd_sc_hd__xor2_4 _5314_ (.A(_0524_),
    .B(_0538_),
    .X(_0540_));
 sky130_fd_sc_hd__and4_1 _5315_ (.A(net170),
    .B(net168),
    .C(_0360_),
    .D(_0361_),
    .X(_0541_));
 sky130_fd_sc_hd__nand4_4 _5316_ (.A(net171),
    .B(net168),
    .C(_0360_),
    .D(_0361_),
    .Y(_0542_));
 sky130_fd_sc_hd__and3_2 _5317_ (.A(_0299_),
    .B(_0300_),
    .C(net112),
    .X(_0543_));
 sky130_fd_sc_hd__or2_4 _5318_ (.A(net47),
    .B(net74),
    .X(_0544_));
 sky130_fd_sc_hd__or2_4 _5319_ (.A(net47),
    .B(net111),
    .X(_0545_));
 sky130_fd_sc_hd__nand3_4 _5320_ (.A(_0299_),
    .B(_0300_),
    .C(net77),
    .Y(_0546_));
 sky130_fd_sc_hd__or2_1 _5321_ (.A(_0545_),
    .B(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__nor2_8 _5322_ (.A(net172),
    .B(_3462_),
    .Y(_0548_));
 sky130_fd_sc_hd__a211o_2 _5323_ (.A1(_3458_),
    .A2(_3461_),
    .B1(net172),
    .C1(_1715_),
    .X(_0549_));
 sky130_fd_sc_hd__nor2_2 _5324_ (.A(net43),
    .B(net109),
    .Y(_0550_));
 sky130_fd_sc_hd__xnor2_4 _5325_ (.A(_0545_),
    .B(_0546_),
    .Y(_0551_));
 sky130_fd_sc_hd__o31a_4 _5326_ (.A1(net43),
    .A2(net109),
    .A3(_0551_),
    .B1(_0547_),
    .X(_0552_));
 sky130_fd_sc_hd__o22ai_4 _5327_ (.A1(_0518_),
    .A2(_0534_),
    .B1(_0536_),
    .B2(_0533_),
    .Y(_0553_));
 sky130_fd_sc_hd__or2_4 _5328_ (.A(net47),
    .B(net78),
    .X(_0554_));
 sky130_fd_sc_hd__and3_4 _5329_ (.A(_0299_),
    .B(_0300_),
    .C(net80),
    .X(_0555_));
 sky130_fd_sc_hd__xnor2_4 _5330_ (.A(_0544_),
    .B(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__nor2_4 _5331_ (.A(net43),
    .B(net111),
    .Y(_0557_));
 sky130_fd_sc_hd__xor2_4 _5332_ (.A(_0556_),
    .B(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__nand2_1 _5333_ (.A(_0553_),
    .B(_0558_),
    .Y(_0559_));
 sky130_fd_sc_hd__nor2_1 _5334_ (.A(_0553_),
    .B(_0558_),
    .Y(_0560_));
 sky130_fd_sc_hd__xor2_4 _5335_ (.A(_0553_),
    .B(_0558_),
    .X(_0561_));
 sky130_fd_sc_hd__xnor2_4 _5336_ (.A(_0552_),
    .B(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__a21oi_4 _5337_ (.A1(_0540_),
    .A2(_0562_),
    .B1(_0539_),
    .Y(_0563_));
 sky130_fd_sc_hd__nand2_1 _5338_ (.A(net65),
    .B(_0474_),
    .Y(_0564_));
 sky130_fd_sc_hd__o21ai_1 _5339_ (.A1(net89),
    .A2(_0416_),
    .B1(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__or2_4 _5340_ (.A(net66),
    .B(_0416_),
    .X(_0566_));
 sky130_fd_sc_hd__o21a_4 _5341_ (.A1(_0519_),
    .A2(_0566_),
    .B1(_0565_),
    .X(_0567_));
 sky130_fd_sc_hd__nor2_4 _5342_ (.A(net85),
    .B(_0410_),
    .Y(_0568_));
 sky130_fd_sc_hd__xor2_4 _5343_ (.A(_0567_),
    .B(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__nor2_8 _5344_ (.A(net70),
    .B(_0516_),
    .Y(_0570_));
 sky130_fd_sc_hd__nand2_2 _5345_ (.A(_0569_),
    .B(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__xor2_4 _5346_ (.A(_0569_),
    .B(_0570_),
    .X(_0572_));
 sky130_fd_sc_hd__xnor2_4 _5347_ (.A(_0523_),
    .B(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__a2bb2o_4 _5348_ (.A1_N(_0546_),
    .A2_N(_0554_),
    .B1(_0556_),
    .B2(_0557_),
    .X(_0574_));
 sky130_fd_sc_hd__a2bb2oi_4 _5349_ (.A1_N(_0518_),
    .A2_N(_0519_),
    .B1(_0520_),
    .B2(_0521_),
    .Y(_0575_));
 sky130_fd_sc_hd__nor2_4 _5350_ (.A(net43),
    .B(net74),
    .Y(_0576_));
 sky130_fd_sc_hd__nor2_8 _5351_ (.A(net47),
    .B(net81),
    .Y(_0577_));
 sky130_fd_sc_hd__and3_2 _5352_ (.A(_0299_),
    .B(_0300_),
    .C(net83),
    .X(_0578_));
 sky130_fd_sc_hd__xnor2_4 _5353_ (.A(_0554_),
    .B(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__xor2_4 _5354_ (.A(_0576_),
    .B(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__nand2b_1 _5355_ (.A_N(_0575_),
    .B(_0580_),
    .Y(_0581_));
 sky130_fd_sc_hd__xnor2_4 _5356_ (.A(_0575_),
    .B(_0580_),
    .Y(_0582_));
 sky130_fd_sc_hd__xor2_4 _5357_ (.A(_0574_),
    .B(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__xnor2_4 _5358_ (.A(_0573_),
    .B(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__nor2_1 _5359_ (.A(_0563_),
    .B(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__xor2_4 _5360_ (.A(_0563_),
    .B(_0584_),
    .X(_0586_));
 sky130_fd_sc_hd__and2_4 _5361_ (.A(net170),
    .B(_0293_),
    .X(_0587_));
 sky130_fd_sc_hd__nand2_2 _5362_ (.A(net170),
    .B(_0293_),
    .Y(_0588_));
 sky130_fd_sc_hd__o21ai_1 _5363_ (.A1(_0205_),
    .A2(_0278_),
    .B1(_0171_),
    .Y(_0589_));
 sky130_fd_sc_hd__nand2_2 _5364_ (.A(_0279_),
    .B(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__or2_4 _5365_ (.A(net103),
    .B(net50),
    .X(_0591_));
 sky130_fd_sc_hd__inv_2 _5366_ (.A(_0591_),
    .Y(_0592_));
 sky130_fd_sc_hd__or2_4 _5367_ (.A(net66),
    .B(net52),
    .X(_0593_));
 sky130_fd_sc_hd__nor2_4 _5368_ (.A(net42),
    .B(net102),
    .Y(_0594_));
 sky130_fd_sc_hd__nand2_4 _5369_ (.A(_0356_),
    .B(_0592_),
    .Y(_0595_));
 sky130_fd_sc_hd__nor2_8 _5370_ (.A(net211),
    .B(net107),
    .Y(_0596_));
 sky130_fd_sc_hd__nor2_8 _5371_ (.A(_3507_),
    .B(net102),
    .Y(_0597_));
 sky130_fd_sc_hd__o21a_4 _5372_ (.A1(_0347_),
    .A2(_0348_),
    .B1(net73),
    .X(_0598_));
 sky130_fd_sc_hd__xor2_4 _5373_ (.A(_0597_),
    .B(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__nor2_4 _5374_ (.A(net70),
    .B(net52),
    .Y(_0600_));
 sky130_fd_sc_hd__xnor2_4 _5375_ (.A(_0599_),
    .B(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__nor2_1 _5376_ (.A(_0595_),
    .B(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__xor2_4 _5377_ (.A(_0595_),
    .B(_0601_),
    .X(_0603_));
 sky130_fd_sc_hd__and3_1 _5378_ (.A(_0233_),
    .B(_0275_),
    .C(_0276_),
    .X(_0604_));
 sky130_fd_sc_hd__or2_4 _5379_ (.A(_0277_),
    .B(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__nor2_4 _5380_ (.A(net202),
    .B(net49),
    .Y(_0606_));
 sky130_fd_sc_hd__a21o_4 _5381_ (.A1(_0603_),
    .A2(_0606_),
    .B1(_0602_),
    .X(_0607_));
 sky130_fd_sc_hd__o21a_4 _5382_ (.A1(_0552_),
    .A2(_0560_),
    .B1(_0559_),
    .X(_0608_));
 sky130_fd_sc_hd__a22o_4 _5383_ (.A1(_0594_),
    .A2(_0596_),
    .B1(_0599_),
    .B2(_0600_),
    .X(_0609_));
 sky130_fd_sc_hd__or2_4 _5384_ (.A(net202),
    .B(net50),
    .X(_0610_));
 sky130_fd_sc_hd__nor2_8 _5385_ (.A(net211),
    .B(net110),
    .Y(_0611_));
 sky130_fd_sc_hd__nor2_4 _5386_ (.A(net42),
    .B(net111),
    .Y(_0612_));
 sky130_fd_sc_hd__nor2_1 _5387_ (.A(_0596_),
    .B(_0612_),
    .Y(_0613_));
 sky130_fd_sc_hd__xor2_4 _5388_ (.A(_0596_),
    .B(_0612_),
    .X(_0614_));
 sky130_fd_sc_hd__xnor2_4 _5389_ (.A(_0610_),
    .B(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hd__nand2_4 _5390_ (.A(_0609_),
    .B(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__xnor2_4 _5391_ (.A(_0609_),
    .B(_0615_),
    .Y(_0617_));
 sky130_fd_sc_hd__nor2_1 _5392_ (.A(_0608_),
    .B(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__nand2_1 _5393_ (.A(_0608_),
    .B(_0617_),
    .Y(_0619_));
 sky130_fd_sc_hd__xnor2_4 _5394_ (.A(_0608_),
    .B(_0617_),
    .Y(_0620_));
 sky130_fd_sc_hd__xnor2_4 _5395_ (.A(_0607_),
    .B(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__a21oi_4 _5396_ (.A1(_0586_),
    .A2(_0621_),
    .B1(_0585_),
    .Y(_0622_));
 sky130_fd_sc_hd__a32oi_4 _5397_ (.A1(_0517_),
    .A2(_0522_),
    .A3(_0572_),
    .B1(_0573_),
    .B2(_0583_),
    .Y(_0623_));
 sky130_fd_sc_hd__and2_1 _5398_ (.A(_0475_),
    .B(_0566_),
    .X(_0624_));
 sky130_fd_sc_hd__xor2_4 _5399_ (.A(_0475_),
    .B(_0566_),
    .X(_0625_));
 sky130_fd_sc_hd__or2_4 _5400_ (.A(net89),
    .B(net46),
    .X(_0626_));
 sky130_fd_sc_hd__xnor2_4 _5401_ (.A(_0625_),
    .B(_0626_),
    .Y(_0627_));
 sky130_fd_sc_hd__xor2_4 _5402_ (.A(_0528_),
    .B(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__xnor2_4 _5403_ (.A(_0571_),
    .B(_0628_),
    .Y(_0629_));
 sky130_fd_sc_hd__a22oi_4 _5404_ (.A1(_0555_),
    .A2(_0577_),
    .B1(_0579_),
    .B2(_0576_),
    .Y(_0630_));
 sky130_fd_sc_hd__a2bb2o_4 _5405_ (.A1_N(_0519_),
    .A2_N(_0566_),
    .B1(_0567_),
    .B2(_0568_),
    .X(_0631_));
 sky130_fd_sc_hd__nor2_4 _5406_ (.A(net43),
    .B(net78),
    .Y(_0632_));
 sky130_fd_sc_hd__xor2_4 _5407_ (.A(_0468_),
    .B(_0577_),
    .X(_0633_));
 sky130_fd_sc_hd__xor2_4 _5408_ (.A(_0632_),
    .B(_0633_),
    .X(_0634_));
 sky130_fd_sc_hd__nand2_1 _5409_ (.A(_0631_),
    .B(_0634_),
    .Y(_0636_));
 sky130_fd_sc_hd__xnor2_4 _5410_ (.A(_0631_),
    .B(_0634_),
    .Y(_0637_));
 sky130_fd_sc_hd__xor2_4 _5411_ (.A(_0630_),
    .B(_0637_),
    .X(_0638_));
 sky130_fd_sc_hd__xnor2_4 _5412_ (.A(_0629_),
    .B(_0638_),
    .Y(_0639_));
 sky130_fd_sc_hd__nor2_1 _5413_ (.A(_0623_),
    .B(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__xor2_4 _5414_ (.A(_0623_),
    .B(_0639_),
    .X(_0641_));
 sky130_fd_sc_hd__a21bo_4 _5415_ (.A1(_0574_),
    .A2(_0582_),
    .B1_N(_0581_),
    .X(_0642_));
 sky130_fd_sc_hd__o2bb2a_4 _5416_ (.A1_N(_0598_),
    .A2_N(_0611_),
    .B1(_0613_),
    .B2(_0610_),
    .X(_0643_));
 sky130_fd_sc_hd__xor2_4 _5417_ (.A(_0499_),
    .B(_0611_),
    .X(_0644_));
 sky130_fd_sc_hd__nor2_4 _5418_ (.A(_0643_),
    .B(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__xnor2_4 _5419_ (.A(_0643_),
    .B(_0644_),
    .Y(_0647_));
 sky130_fd_sc_hd__nand2b_1 _5420_ (.A_N(_0647_),
    .B(_0642_),
    .Y(_0648_));
 sky130_fd_sc_hd__xor2_4 _5421_ (.A(_0642_),
    .B(_0647_),
    .X(_0649_));
 sky130_fd_sc_hd__xor2_4 _5422_ (.A(_0616_),
    .B(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__xnor2_2 _5423_ (.A(_0641_),
    .B(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__or2_1 _5424_ (.A(_0622_),
    .B(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__a21o_1 _5425_ (.A1(_0607_),
    .A2(_0619_),
    .B1(_0618_),
    .X(_0653_));
 sky130_fd_sc_hd__xor2_2 _5426_ (.A(_0622_),
    .B(_0651_),
    .X(_0654_));
 sky130_fd_sc_hd__nand2_1 _5427_ (.A(_0653_),
    .B(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__o21ai_2 _5428_ (.A1(_0616_),
    .A2(_0649_),
    .B1(_0648_),
    .Y(_0656_));
 sky130_fd_sc_hd__a21o_1 _5429_ (.A1(_0641_),
    .A2(_0650_),
    .B1(_0640_),
    .X(_0658_));
 sky130_fd_sc_hd__a32oi_4 _5430_ (.A1(_0569_),
    .A2(_0570_),
    .A3(_0628_),
    .B1(_0629_),
    .B2(_0638_),
    .Y(_0659_));
 sky130_fd_sc_hd__xnor2_2 _5431_ (.A(_0477_),
    .B(_0479_),
    .Y(_0660_));
 sky130_fd_sc_hd__and3_2 _5432_ (.A(_0528_),
    .B(_0627_),
    .C(_0660_),
    .X(_0661_));
 sky130_fd_sc_hd__a21oi_2 _5433_ (.A1(_0528_),
    .A2(_0627_),
    .B1(_0660_),
    .Y(_0662_));
 sky130_fd_sc_hd__nor2_4 _5434_ (.A(_0661_),
    .B(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__a22o_4 _5435_ (.A1(_0468_),
    .A2(_0577_),
    .B1(_0632_),
    .B2(_0633_),
    .X(_0664_));
 sky130_fd_sc_hd__o22a_4 _5436_ (.A1(_0417_),
    .A2(_0564_),
    .B1(_0624_),
    .B2(_0626_),
    .X(_0665_));
 sky130_fd_sc_hd__xor2_4 _5437_ (.A(_0470_),
    .B(_0471_),
    .X(_0666_));
 sky130_fd_sc_hd__and2b_1 _5438_ (.A_N(_0665_),
    .B(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__xnor2_4 _5439_ (.A(_0665_),
    .B(_0666_),
    .Y(_0669_));
 sky130_fd_sc_hd__xor2_4 _5440_ (.A(_0664_),
    .B(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__xnor2_4 _5441_ (.A(_0663_),
    .B(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__nor2_1 _5442_ (.A(_0659_),
    .B(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__xor2_4 _5443_ (.A(_0659_),
    .B(_0671_),
    .X(_0673_));
 sky130_fd_sc_hd__o21a_4 _5444_ (.A1(_0630_),
    .A2(_0637_),
    .B1(_0636_),
    .X(_0674_));
 sky130_fd_sc_hd__or4_4 _5445_ (.A(net211),
    .B(net80),
    .C(_0499_),
    .D(net111),
    .X(_0675_));
 sky130_fd_sc_hd__or3_1 _5446_ (.A(_0433_),
    .B(_0499_),
    .C(_0611_),
    .X(_0676_));
 sky130_fd_sc_hd__o211a_4 _5447_ (.A1(_0432_),
    .A2(_0500_),
    .B1(_0675_),
    .C1(_0676_),
    .X(_0677_));
 sky130_fd_sc_hd__nand2b_1 _5448_ (.A_N(_0674_),
    .B(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__xnor2_4 _5449_ (.A(_0674_),
    .B(_0677_),
    .Y(_0680_));
 sky130_fd_sc_hd__xor2_4 _5450_ (.A(_0645_),
    .B(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__xor2_2 _5451_ (.A(_0673_),
    .B(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__nand2_1 _5452_ (.A(_0658_),
    .B(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__xnor2_1 _5453_ (.A(_0658_),
    .B(_0682_),
    .Y(_0684_));
 sky130_fd_sc_hd__nand2b_1 _5454_ (.A_N(_0684_),
    .B(_0656_),
    .Y(_0685_));
 sky130_fd_sc_hd__xor2_1 _5455_ (.A(_0656_),
    .B(_0684_),
    .X(_0686_));
 sky130_fd_sc_hd__a21o_2 _5456_ (.A1(_0652_),
    .A2(_0655_),
    .B1(_0686_),
    .X(_0687_));
 sky130_fd_sc_hd__a21bo_4 _5457_ (.A1(_0645_),
    .A2(_0680_),
    .B1_N(_0678_),
    .X(_0688_));
 sky130_fd_sc_hd__a21o_2 _5458_ (.A1(_0673_),
    .A2(_0681_),
    .B1(_0672_),
    .X(_0689_));
 sky130_fd_sc_hd__xnor2_4 _5459_ (.A(_0484_),
    .B(_0485_),
    .Y(_0691_));
 sky130_fd_sc_hd__a21o_4 _5460_ (.A1(_0663_),
    .A2(_0670_),
    .B1(_0661_),
    .X(_0692_));
 sky130_fd_sc_hd__and2b_1 _5461_ (.A_N(_0691_),
    .B(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__xnor2_4 _5462_ (.A(_0691_),
    .B(_0692_),
    .Y(_0694_));
 sky130_fd_sc_hd__a21o_4 _5463_ (.A1(_0664_),
    .A2(_0669_),
    .B1(_0667_),
    .X(_0695_));
 sky130_fd_sc_hd__and3b_1 _5464_ (.A_N(_0500_),
    .B(_0432_),
    .C(_0375_),
    .X(_0696_));
 sky130_fd_sc_hd__nand2_2 _5465_ (.A(_0374_),
    .B(_0433_),
    .Y(_0697_));
 sky130_fd_sc_hd__nor2_2 _5466_ (.A(_0501_),
    .B(_0696_),
    .Y(_0698_));
 sky130_fd_sc_hd__nand2_2 _5467_ (.A(_0697_),
    .B(_0698_),
    .Y(_0699_));
 sky130_fd_sc_hd__xnor2_4 _5468_ (.A(_0695_),
    .B(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hd__and2b_1 _5469_ (.A_N(_0675_),
    .B(_0700_),
    .X(_0702_));
 sky130_fd_sc_hd__xnor2_4 _5470_ (.A(_0675_),
    .B(_0700_),
    .Y(_0703_));
 sky130_fd_sc_hd__xnor2_4 _5471_ (.A(_0694_),
    .B(_0703_),
    .Y(_0704_));
 sky130_fd_sc_hd__and2b_1 _5472_ (.A_N(_0704_),
    .B(_0689_),
    .X(_0705_));
 sky130_fd_sc_hd__xnor2_4 _5473_ (.A(_0689_),
    .B(_0704_),
    .Y(_0706_));
 sky130_fd_sc_hd__xnor2_2 _5474_ (.A(_0688_),
    .B(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__a21o_4 _5475_ (.A1(_0683_),
    .A2(_0685_),
    .B1(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__inv_2 _5476_ (.A(_0708_),
    .Y(_0709_));
 sky130_fd_sc_hd__nand3_1 _5477_ (.A(_0683_),
    .B(_0685_),
    .C(_0707_),
    .Y(_0710_));
 sky130_fd_sc_hd__and2_1 _5478_ (.A(_0708_),
    .B(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__and2b_1 _5479_ (.A_N(_0687_),
    .B(_0711_),
    .X(_0713_));
 sky130_fd_sc_hd__xor2_2 _5480_ (.A(_0687_),
    .B(_0711_),
    .X(_0714_));
 sky130_fd_sc_hd__a31o_4 _5481_ (.A1(_0695_),
    .A2(_0697_),
    .A3(_0698_),
    .B1(_0702_),
    .X(_0715_));
 sky130_fd_sc_hd__xnor2_2 _5482_ (.A(_0488_),
    .B(_0502_),
    .Y(_0716_));
 sky130_fd_sc_hd__a21oi_2 _5483_ (.A1(_0694_),
    .A2(_0703_),
    .B1(_0693_),
    .Y(_0717_));
 sky130_fd_sc_hd__nor2_2 _5484_ (.A(_0716_),
    .B(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__nand2_2 _5485_ (.A(_0716_),
    .B(_0717_),
    .Y(_0719_));
 sky130_fd_sc_hd__and2b_2 _5486_ (.A_N(_0718_),
    .B(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__xnor2_4 _5487_ (.A(_0715_),
    .B(_0720_),
    .Y(_0721_));
 sky130_fd_sc_hd__a21oi_4 _5488_ (.A1(_0688_),
    .A2(_0706_),
    .B1(_0705_),
    .Y(_0722_));
 sky130_fd_sc_hd__nor2_2 _5489_ (.A(_0721_),
    .B(_0722_),
    .Y(_0724_));
 sky130_fd_sc_hd__xor2_4 _5490_ (.A(_0721_),
    .B(_0722_),
    .X(_0725_));
 sky130_fd_sc_hd__xnor2_4 _5491_ (.A(_0708_),
    .B(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__xnor2_4 _5492_ (.A(_0505_),
    .B(_0507_),
    .Y(_0727_));
 sky130_fd_sc_hd__a21oi_4 _5493_ (.A1(_0715_),
    .A2(_0719_),
    .B1(_0718_),
    .Y(_0728_));
 sky130_fd_sc_hd__or2_4 _5494_ (.A(_0727_),
    .B(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__xor2_4 _5495_ (.A(_0727_),
    .B(_0728_),
    .X(_0730_));
 sky130_fd_sc_hd__nand2_1 _5496_ (.A(_0724_),
    .B(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__xnor2_2 _5497_ (.A(_0724_),
    .B(_0730_),
    .Y(_0732_));
 sky130_fd_sc_hd__xnor2_4 _5498_ (.A(_0465_),
    .B(_0508_),
    .Y(_0733_));
 sky130_fd_sc_hd__xnor2_4 _5499_ (.A(_0729_),
    .B(_0733_),
    .Y(_0735_));
 sky130_fd_sc_hd__or2_1 _5500_ (.A(_0732_),
    .B(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__nand2b_1 _5501_ (.A_N(_0714_),
    .B(_0726_),
    .Y(_0737_));
 sky130_fd_sc_hd__or2_1 _5502_ (.A(_0736_),
    .B(_0737_),
    .X(_0738_));
 sky130_fd_sc_hd__xnor2_4 _5503_ (.A(_0540_),
    .B(_0562_),
    .Y(_0739_));
 sky130_fd_sc_hd__xnor2_4 _5504_ (.A(_0532_),
    .B(_0537_),
    .Y(_0740_));
 sky130_fd_sc_hd__o21ba_1 _5505_ (.A1(net85),
    .A2(net53),
    .B1_N(_0529_),
    .X(_0741_));
 sky130_fd_sc_hd__a21o_1 _5506_ (.A1(_0527_),
    .A2(_0528_),
    .B1(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__o21ai_4 _5507_ (.A1(_0271_),
    .A2(_0272_),
    .B1(_0256_),
    .Y(_0743_));
 sky130_fd_sc_hd__and2_4 _5508_ (.A(_0273_),
    .B(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__and3_4 _5509_ (.A(_3464_),
    .B(_0273_),
    .C(_0743_),
    .X(_0745_));
 sky130_fd_sc_hd__nor2_2 _5510_ (.A(net81),
    .B(net53),
    .Y(_0746_));
 sky130_fd_sc_hd__o2bb2a_2 _5511_ (.A1_N(_0744_),
    .A2_N(net199),
    .B1(net70),
    .B2(net54),
    .X(_0747_));
 sky130_fd_sc_hd__a21oi_4 _5512_ (.A1(_0529_),
    .A2(_0745_),
    .B1(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__a22oi_4 _5513_ (.A1(_0529_),
    .A2(_0745_),
    .B1(_0746_),
    .B2(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__nor2_4 _5514_ (.A(_0742_),
    .B(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__and3_2 _5515_ (.A(_0414_),
    .B(_0415_),
    .C(net80),
    .X(_0751_));
 sky130_fd_sc_hd__or2_2 _5516_ (.A(_0416_),
    .B(net78),
    .X(_0752_));
 sky130_fd_sc_hd__nand2_2 _5517_ (.A(net80),
    .B(net48),
    .Y(_0753_));
 sky130_fd_sc_hd__xnor2_4 _5518_ (.A(_0534_),
    .B(_0751_),
    .Y(_0754_));
 sky130_fd_sc_hd__nor2_4 _5519_ (.A(net46),
    .B(net74),
    .Y(_0755_));
 sky130_fd_sc_hd__nand2_1 _5520_ (.A(_0754_),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__xor2_4 _5521_ (.A(_0754_),
    .B(_0755_),
    .X(_0757_));
 sky130_fd_sc_hd__and2_1 _5522_ (.A(_0742_),
    .B(_0749_),
    .X(_0758_));
 sky130_fd_sc_hd__nor2_4 _5523_ (.A(_0750_),
    .B(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__a21oi_4 _5524_ (.A1(_0757_),
    .A2(_0759_),
    .B1(_0750_),
    .Y(_0760_));
 sky130_fd_sc_hd__nor2_2 _5525_ (.A(_0740_),
    .B(_0760_),
    .Y(_0761_));
 sky130_fd_sc_hd__xor2_4 _5526_ (.A(_0740_),
    .B(_0760_),
    .X(_0762_));
 sky130_fd_sc_hd__or2_4 _5527_ (.A(_0301_),
    .B(net108),
    .X(_0763_));
 sky130_fd_sc_hd__or2_4 _5528_ (.A(net47),
    .B(net108),
    .X(_0764_));
 sky130_fd_sc_hd__nor2_1 _5529_ (.A(net43),
    .B(net102),
    .Y(_0765_));
 sky130_fd_sc_hd__or2_4 _5530_ (.A(net43),
    .B(net102),
    .X(_0766_));
 sky130_fd_sc_hd__xnor2_4 _5531_ (.A(_0543_),
    .B(_0764_),
    .Y(_0767_));
 sky130_fd_sc_hd__a2bb2oi_4 _5532_ (.A1_N(_0545_),
    .A2_N(_0763_),
    .B1(_0765_),
    .B2(_0767_),
    .Y(_0768_));
 sky130_fd_sc_hd__o21ai_4 _5533_ (.A1(_0534_),
    .A2(_0752_),
    .B1(_0756_),
    .Y(_0769_));
 sky130_fd_sc_hd__xnor2_4 _5534_ (.A(_0550_),
    .B(_0551_),
    .Y(_0770_));
 sky130_fd_sc_hd__nand2_1 _5535_ (.A(_0769_),
    .B(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__nor2_1 _5536_ (.A(_0769_),
    .B(_0770_),
    .Y(_0772_));
 sky130_fd_sc_hd__xor2_4 _5537_ (.A(_0769_),
    .B(_0770_),
    .X(_0773_));
 sky130_fd_sc_hd__xnor2_4 _5538_ (.A(_0768_),
    .B(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__a21oi_4 _5539_ (.A1(_0762_),
    .A2(_0774_),
    .B1(_0761_),
    .Y(_0776_));
 sky130_fd_sc_hd__nor2_1 _5540_ (.A(_0739_),
    .B(_0776_),
    .Y(_0777_));
 sky130_fd_sc_hd__or2_4 _5541_ (.A(net70),
    .B(net49),
    .X(_0778_));
 sky130_fd_sc_hd__xnor2_4 _5542_ (.A(_0593_),
    .B(_0594_),
    .Y(_0779_));
 sky130_fd_sc_hd__nand2b_2 _5543_ (.A_N(_0778_),
    .B(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__o21ai_4 _5544_ (.A1(_0768_),
    .A2(_0772_),
    .B1(_0771_),
    .Y(_0781_));
 sky130_fd_sc_hd__xor2_4 _5545_ (.A(_0603_),
    .B(_0606_),
    .X(_0782_));
 sky130_fd_sc_hd__nand2_1 _5546_ (.A(_0781_),
    .B(_0782_),
    .Y(_0783_));
 sky130_fd_sc_hd__xnor2_4 _5547_ (.A(_0781_),
    .B(_0782_),
    .Y(_0784_));
 sky130_fd_sc_hd__xor2_2 _5548_ (.A(_0780_),
    .B(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__xor2_2 _5549_ (.A(_0739_),
    .B(_0776_),
    .X(_0787_));
 sky130_fd_sc_hd__a21o_1 _5550_ (.A1(_0785_),
    .A2(_0787_),
    .B1(_0777_),
    .X(_0788_));
 sky130_fd_sc_hd__xnor2_2 _5551_ (.A(_0586_),
    .B(_0621_),
    .Y(_0789_));
 sky130_fd_sc_hd__nand2b_1 _5552_ (.A_N(_0789_),
    .B(_0788_),
    .Y(_0790_));
 sky130_fd_sc_hd__o21ai_2 _5553_ (.A1(_0780_),
    .A2(_0784_),
    .B1(_0783_),
    .Y(_0791_));
 sky130_fd_sc_hd__xnor2_1 _5554_ (.A(_0788_),
    .B(_0789_),
    .Y(_0792_));
 sky130_fd_sc_hd__nand2_2 _5555_ (.A(_0791_),
    .B(_0792_),
    .Y(_0793_));
 sky130_fd_sc_hd__xnor2_1 _5556_ (.A(_0653_),
    .B(_0654_),
    .Y(_0794_));
 sky130_fd_sc_hd__a21o_2 _5557_ (.A1(_0790_),
    .A2(_0793_),
    .B1(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__nand3_1 _5558_ (.A(_0790_),
    .B(_0793_),
    .C(_0794_),
    .Y(_0796_));
 sky130_fd_sc_hd__and2_2 _5559_ (.A(_0795_),
    .B(_0796_),
    .X(_0798_));
 sky130_fd_sc_hd__xnor2_1 _5560_ (.A(_0785_),
    .B(_0787_),
    .Y(_0799_));
 sky130_fd_sc_hd__xnor2_4 _5561_ (.A(_0762_),
    .B(_0774_),
    .Y(_0800_));
 sky130_fd_sc_hd__xnor2_2 _5562_ (.A(_0757_),
    .B(_0759_),
    .Y(_0801_));
 sky130_fd_sc_hd__xnor2_1 _5563_ (.A(_0746_),
    .B(_0748_),
    .Y(_0802_));
 sky130_fd_sc_hd__nor2_8 _5564_ (.A(net66),
    .B(net54),
    .Y(_0803_));
 sky130_fd_sc_hd__nor2_4 _5565_ (.A(net78),
    .B(net53),
    .Y(_0804_));
 sky130_fd_sc_hd__xor2_4 _5566_ (.A(_0745_),
    .B(_0803_),
    .X(_0805_));
 sky130_fd_sc_hd__a22o_1 _5567_ (.A1(_0745_),
    .A2(_0803_),
    .B1(_0804_),
    .B2(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__and2b_2 _5568_ (.A_N(_0802_),
    .B(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__and2b_1 _5569_ (.A_N(_0806_),
    .B(_0802_),
    .X(_0809_));
 sky130_fd_sc_hd__nor2_4 _5570_ (.A(_0807_),
    .B(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__or2_4 _5571_ (.A(net46),
    .B(net111),
    .X(_0811_));
 sky130_fd_sc_hd__and3_2 _5572_ (.A(_0414_),
    .B(_0415_),
    .C(net76),
    .X(_0812_));
 sky130_fd_sc_hd__nand2_4 _5573_ (.A(net48),
    .B(net76),
    .Y(_0813_));
 sky130_fd_sc_hd__nor2_1 _5574_ (.A(_0752_),
    .B(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__xnor2_4 _5575_ (.A(_0753_),
    .B(_0812_),
    .Y(_0815_));
 sky130_fd_sc_hd__xnor2_4 _5576_ (.A(_0811_),
    .B(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__a21oi_2 _5577_ (.A1(_0810_),
    .A2(_0816_),
    .B1(_0807_),
    .Y(_0817_));
 sky130_fd_sc_hd__nor2_2 _5578_ (.A(_0801_),
    .B(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__and2_1 _5579_ (.A(_0801_),
    .B(_0817_),
    .X(_0819_));
 sky130_fd_sc_hd__nor2_4 _5580_ (.A(_0818_),
    .B(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__nor2_2 _5581_ (.A(_0301_),
    .B(net102),
    .Y(_0821_));
 sky130_fd_sc_hd__or2_4 _5582_ (.A(net47),
    .B(net102),
    .X(_0822_));
 sky130_fd_sc_hd__or2_4 _5583_ (.A(_0763_),
    .B(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__a31o_4 _5584_ (.A1(_0411_),
    .A2(net112),
    .A3(_0815_),
    .B1(_0814_),
    .X(_0824_));
 sky130_fd_sc_hd__xnor2_4 _5585_ (.A(_0766_),
    .B(_0767_),
    .Y(_0825_));
 sky130_fd_sc_hd__nand2_1 _5586_ (.A(_0824_),
    .B(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__nor2_1 _5587_ (.A(_0824_),
    .B(_0825_),
    .Y(_0827_));
 sky130_fd_sc_hd__xor2_4 _5588_ (.A(_0824_),
    .B(_0825_),
    .X(_0828_));
 sky130_fd_sc_hd__xnor2_4 _5589_ (.A(_0823_),
    .B(_0828_),
    .Y(_0829_));
 sky130_fd_sc_hd__a21o_2 _5590_ (.A1(_0820_),
    .A2(_0829_),
    .B1(_0818_),
    .X(_0830_));
 sky130_fd_sc_hd__nand2b_1 _5591_ (.A_N(_0800_),
    .B(_0830_),
    .Y(_0831_));
 sky130_fd_sc_hd__or2_4 _5592_ (.A(net89),
    .B(net49),
    .X(_0832_));
 sky130_fd_sc_hd__or2_1 _5593_ (.A(net89),
    .B(net52),
    .X(_0833_));
 sky130_fd_sc_hd__or2_4 _5594_ (.A(_0593_),
    .B(_0832_),
    .X(_0834_));
 sky130_fd_sc_hd__o21ai_4 _5595_ (.A1(_0823_),
    .A2(_0827_),
    .B1(_0826_),
    .Y(_0835_));
 sky130_fd_sc_hd__xnor2_4 _5596_ (.A(_0778_),
    .B(_0779_),
    .Y(_0836_));
 sky130_fd_sc_hd__xor2_4 _5597_ (.A(_0835_),
    .B(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__nand2b_1 _5598_ (.A_N(_0834_),
    .B(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__xnor2_4 _5599_ (.A(_0834_),
    .B(_0837_),
    .Y(_0839_));
 sky130_fd_sc_hd__xnor2_4 _5600_ (.A(_0800_),
    .B(_0830_),
    .Y(_0840_));
 sky130_fd_sc_hd__a21boi_2 _5601_ (.A1(_0839_),
    .A2(_0840_),
    .B1_N(_0831_),
    .Y(_0841_));
 sky130_fd_sc_hd__or2_4 _5602_ (.A(_0799_),
    .B(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__a21bo_4 _5603_ (.A1(_0835_),
    .A2(_0836_),
    .B1_N(_0838_),
    .X(_0843_));
 sky130_fd_sc_hd__nand2_1 _5604_ (.A(_0799_),
    .B(_0841_),
    .Y(_0844_));
 sky130_fd_sc_hd__nand2_2 _5605_ (.A(_0842_),
    .B(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__nand2b_2 _5606_ (.A_N(_0845_),
    .B(_0843_),
    .Y(_0846_));
 sky130_fd_sc_hd__or2_1 _5607_ (.A(_0791_),
    .B(_0792_),
    .X(_0847_));
 sky130_fd_sc_hd__nand2_2 _5608_ (.A(_0793_),
    .B(_0847_),
    .Y(_0848_));
 sky130_fd_sc_hd__a21oi_4 _5609_ (.A1(_0842_),
    .A2(_0846_),
    .B1(_0848_),
    .Y(_0849_));
 sky130_fd_sc_hd__nand2_1 _5610_ (.A(_0798_),
    .B(_0849_),
    .Y(_0850_));
 sky130_fd_sc_hd__xnor2_4 _5611_ (.A(_0798_),
    .B(_0849_),
    .Y(_0851_));
 sky130_fd_sc_hd__nand3_1 _5612_ (.A(_0652_),
    .B(_0655_),
    .C(_0686_),
    .Y(_0852_));
 sky130_fd_sc_hd__nand2_2 _5613_ (.A(_0687_),
    .B(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__xnor2_2 _5614_ (.A(_0795_),
    .B(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__nor2_2 _5615_ (.A(_0851_),
    .B(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__and3_1 _5616_ (.A(_0842_),
    .B(_0846_),
    .C(_0848_),
    .X(_0856_));
 sky130_fd_sc_hd__nor2_4 _5617_ (.A(_0849_),
    .B(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__xnor2_4 _5618_ (.A(_0839_),
    .B(_0840_),
    .Y(_0858_));
 sky130_fd_sc_hd__xnor2_4 _5619_ (.A(_0804_),
    .B(_0805_),
    .Y(_0859_));
 sky130_fd_sc_hd__and3_2 _5620_ (.A(_0273_),
    .B(net88),
    .C(_0743_),
    .X(_0860_));
 sky130_fd_sc_hd__nor2_1 _5621_ (.A(net89),
    .B(net54),
    .Y(_0861_));
 sky130_fd_sc_hd__nor2_1 _5622_ (.A(net74),
    .B(net53),
    .Y(_0862_));
 sky130_fd_sc_hd__a21oi_1 _5623_ (.A1(net64),
    .A2(_0744_),
    .B1(_0861_),
    .Y(_0863_));
 sky130_fd_sc_hd__a21oi_2 _5624_ (.A1(_0803_),
    .A2(_0860_),
    .B1(_0863_),
    .Y(_0864_));
 sky130_fd_sc_hd__a22o_4 _5625_ (.A1(_0803_),
    .A2(_0860_),
    .B1(_0862_),
    .B2(_0864_),
    .X(_0865_));
 sky130_fd_sc_hd__and2b_1 _5626_ (.A_N(_0859_),
    .B(_0865_),
    .X(_0866_));
 sky130_fd_sc_hd__xnor2_4 _5627_ (.A(_0859_),
    .B(_0865_),
    .Y(_0867_));
 sky130_fd_sc_hd__or2_4 _5628_ (.A(net46),
    .B(net108),
    .X(_0868_));
 sky130_fd_sc_hd__and3_2 _5629_ (.A(_0414_),
    .B(_0415_),
    .C(net112),
    .X(_0869_));
 sky130_fd_sc_hd__nand2_4 _5630_ (.A(net48),
    .B(net112),
    .Y(_0870_));
 sky130_fd_sc_hd__and3_1 _5631_ (.A(net48),
    .B(net112),
    .C(_0812_),
    .X(_0871_));
 sky130_fd_sc_hd__xnor2_4 _5632_ (.A(_0813_),
    .B(_0869_),
    .Y(_0872_));
 sky130_fd_sc_hd__xnor2_4 _5633_ (.A(_0868_),
    .B(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__a21o_4 _5634_ (.A1(_0867_),
    .A2(_0873_),
    .B1(_0866_),
    .X(_0874_));
 sky130_fd_sc_hd__xor2_4 _5635_ (.A(_0810_),
    .B(_0816_),
    .X(_0875_));
 sky130_fd_sc_hd__nand2_1 _5636_ (.A(_0874_),
    .B(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__xor2_4 _5637_ (.A(_0874_),
    .B(_0875_),
    .X(_0877_));
 sky130_fd_sc_hd__a31oi_4 _5638_ (.A1(_0411_),
    .A2(net73),
    .A3(_0872_),
    .B1(_0871_),
    .Y(_0878_));
 sky130_fd_sc_hd__xnor2_4 _5639_ (.A(_0763_),
    .B(_0822_),
    .Y(_0879_));
 sky130_fd_sc_hd__or2_4 _5640_ (.A(_0878_),
    .B(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__xor2_4 _5641_ (.A(_0878_),
    .B(_0879_),
    .X(_0881_));
 sky130_fd_sc_hd__a21bo_4 _5642_ (.A1(_0877_),
    .A2(_0881_),
    .B1_N(_0876_),
    .X(_0882_));
 sky130_fd_sc_hd__xnor2_4 _5643_ (.A(_0820_),
    .B(_0829_),
    .Y(_0883_));
 sky130_fd_sc_hd__and2b_1 _5644_ (.A_N(_0883_),
    .B(_0882_),
    .X(_0884_));
 sky130_fd_sc_hd__xnor2_4 _5645_ (.A(_0882_),
    .B(_0883_),
    .Y(_0885_));
 sky130_fd_sc_hd__or2_2 _5646_ (.A(net85),
    .B(net49),
    .X(_0886_));
 sky130_fd_sc_hd__nor2_8 _5647_ (.A(net85),
    .B(net52),
    .Y(_0887_));
 sky130_fd_sc_hd__or2_4 _5648_ (.A(_0833_),
    .B(_0886_),
    .X(_0888_));
 sky130_fd_sc_hd__o21ai_1 _5649_ (.A1(net67),
    .A2(net49),
    .B1(_0833_),
    .Y(_0889_));
 sky130_fd_sc_hd__and2_2 _5650_ (.A(_0834_),
    .B(_0889_),
    .X(_0890_));
 sky130_fd_sc_hd__inv_2 _5651_ (.A(_0890_),
    .Y(_0891_));
 sky130_fd_sc_hd__xnor2_4 _5652_ (.A(_0880_),
    .B(_0890_),
    .Y(_0892_));
 sky130_fd_sc_hd__nand2b_1 _5653_ (.A_N(_0888_),
    .B(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__xnor2_4 _5654_ (.A(_0888_),
    .B(_0892_),
    .Y(_0894_));
 sky130_fd_sc_hd__a21oi_4 _5655_ (.A1(_0885_),
    .A2(_0894_),
    .B1(_0884_),
    .Y(_0895_));
 sky130_fd_sc_hd__o21ai_4 _5656_ (.A1(_0880_),
    .A2(_0891_),
    .B1(_0893_),
    .Y(_0896_));
 sky130_fd_sc_hd__xnor2_4 _5657_ (.A(_0858_),
    .B(_0895_),
    .Y(_0897_));
 sky130_fd_sc_hd__nand2b_1 _5658_ (.A_N(_0897_),
    .B(_0896_),
    .Y(_0898_));
 sky130_fd_sc_hd__o21ai_4 _5659_ (.A1(_0858_),
    .A2(_0895_),
    .B1(_0898_),
    .Y(_0899_));
 sky130_fd_sc_hd__xor2_4 _5660_ (.A(_0843_),
    .B(_0845_),
    .X(_0900_));
 sky130_fd_sc_hd__and2b_2 _5661_ (.A_N(_0900_),
    .B(_0899_),
    .X(_0901_));
 sky130_fd_sc_hd__xor2_4 _5662_ (.A(_0896_),
    .B(_0897_),
    .X(_0902_));
 sky130_fd_sc_hd__xnor2_1 _5663_ (.A(_0862_),
    .B(_0864_),
    .Y(_0903_));
 sky130_fd_sc_hd__and3_1 _5664_ (.A(_0273_),
    .B(_0364_),
    .C(_0743_),
    .X(_0904_));
 sky130_fd_sc_hd__or2_4 _5665_ (.A(net53),
    .B(net110),
    .X(_0905_));
 sky130_fd_sc_hd__nor2_1 _5666_ (.A(_0527_),
    .B(_0860_),
    .Y(_0906_));
 sky130_fd_sc_hd__a21o_2 _5667_ (.A1(_0861_),
    .A2(_0904_),
    .B1(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__o2bb2ai_1 _5668_ (.A1_N(_0527_),
    .A2_N(_0860_),
    .B1(_0905_),
    .B2(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__and2b_2 _5669_ (.A_N(_0903_),
    .B(_0908_),
    .X(_0909_));
 sky130_fd_sc_hd__and2b_1 _5670_ (.A_N(_0908_),
    .B(_0903_),
    .X(_0910_));
 sky130_fd_sc_hd__nor2_4 _5671_ (.A(_0909_),
    .B(_0910_),
    .Y(_0911_));
 sky130_fd_sc_hd__nor2_2 _5672_ (.A(net46),
    .B(net102),
    .Y(_0912_));
 sky130_fd_sc_hd__nand3_4 _5673_ (.A(_0414_),
    .B(_0415_),
    .C(net73),
    .Y(_0913_));
 sky130_fd_sc_hd__nand2_2 _5674_ (.A(net48),
    .B(net73),
    .Y(_0914_));
 sky130_fd_sc_hd__or2_1 _5675_ (.A(_0870_),
    .B(_0913_),
    .X(_0915_));
 sky130_fd_sc_hd__xnor2_4 _5676_ (.A(_0870_),
    .B(_0913_),
    .Y(_0916_));
 sky130_fd_sc_hd__xnor2_4 _5677_ (.A(_0912_),
    .B(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__a21oi_4 _5678_ (.A1(_0911_),
    .A2(_0917_),
    .B1(_0909_),
    .Y(_0918_));
 sky130_fd_sc_hd__xnor2_4 _5679_ (.A(_0867_),
    .B(_0873_),
    .Y(_0919_));
 sky130_fd_sc_hd__nor2_1 _5680_ (.A(_0918_),
    .B(_0919_),
    .Y(_0920_));
 sky130_fd_sc_hd__xor2_4 _5681_ (.A(_0918_),
    .B(_0919_),
    .X(_0921_));
 sky130_fd_sc_hd__o31a_4 _5682_ (.A1(net46),
    .A2(net102),
    .A3(_0916_),
    .B1(_0915_),
    .X(_0922_));
 sky130_fd_sc_hd__or3_4 _5683_ (.A(_0301_),
    .B(net102),
    .C(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__xnor2_4 _5684_ (.A(_0821_),
    .B(_0922_),
    .Y(_0924_));
 sky130_fd_sc_hd__a21o_4 _5685_ (.A1(_0921_),
    .A2(_0924_),
    .B1(_0920_),
    .X(_0925_));
 sky130_fd_sc_hd__xor2_4 _5686_ (.A(_0877_),
    .B(_0881_),
    .X(_0926_));
 sky130_fd_sc_hd__nand2_1 _5687_ (.A(_0925_),
    .B(_0926_),
    .Y(_0927_));
 sky130_fd_sc_hd__xor2_4 _5688_ (.A(_0925_),
    .B(_0926_),
    .X(_0928_));
 sky130_fd_sc_hd__nor2_4 _5689_ (.A(net81),
    .B(net49),
    .Y(_0929_));
 sky130_fd_sc_hd__nor2_1 _5690_ (.A(net81),
    .B(net51),
    .Y(_0930_));
 sky130_fd_sc_hd__nand2_4 _5691_ (.A(_0887_),
    .B(_0929_),
    .Y(_0931_));
 sky130_fd_sc_hd__xnor2_4 _5692_ (.A(_0832_),
    .B(_0887_),
    .Y(_0932_));
 sky130_fd_sc_hd__and2b_1 _5693_ (.A_N(_0923_),
    .B(_0932_),
    .X(_0933_));
 sky130_fd_sc_hd__xnor2_4 _5694_ (.A(_0923_),
    .B(_0932_),
    .Y(_0934_));
 sky130_fd_sc_hd__xnor2_4 _5695_ (.A(_0931_),
    .B(_0934_),
    .Y(_0935_));
 sky130_fd_sc_hd__a21bo_4 _5696_ (.A1(_0928_),
    .A2(_0935_),
    .B1_N(_0927_),
    .X(_0936_));
 sky130_fd_sc_hd__xnor2_4 _5697_ (.A(_0885_),
    .B(_0894_),
    .Y(_0937_));
 sky130_fd_sc_hd__nand2b_1 _5698_ (.A_N(_0937_),
    .B(_0936_),
    .Y(_0938_));
 sky130_fd_sc_hd__a31o_4 _5699_ (.A1(_0887_),
    .A2(_0929_),
    .A3(_0934_),
    .B1(_0933_),
    .X(_0939_));
 sky130_fd_sc_hd__xnor2_4 _5700_ (.A(_0936_),
    .B(_0937_),
    .Y(_0940_));
 sky130_fd_sc_hd__a21boi_4 _5701_ (.A1(_0939_),
    .A2(_0940_),
    .B1_N(_0938_),
    .Y(_0941_));
 sky130_fd_sc_hd__nor2_1 _5702_ (.A(_0902_),
    .B(_0941_),
    .Y(_0942_));
 sky130_fd_sc_hd__nand2_4 _5703_ (.A(_0234_),
    .B(_0274_),
    .Y(_0943_));
 sky130_fd_sc_hd__and2_4 _5704_ (.A(_0275_),
    .B(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__and3_2 _5705_ (.A(_0275_),
    .B(net199),
    .C(_0943_),
    .X(_0945_));
 sky130_fd_sc_hd__xor2_4 _5706_ (.A(_0902_),
    .B(_0941_),
    .X(_0946_));
 sky130_fd_sc_hd__a21o_1 _5707_ (.A1(_0945_),
    .A2(_0946_),
    .B1(_0942_),
    .X(_0947_));
 sky130_fd_sc_hd__xor2_1 _5708_ (.A(_0899_),
    .B(_0900_),
    .X(_0948_));
 sky130_fd_sc_hd__and2b_1 _5709_ (.A_N(_0948_),
    .B(_0947_),
    .X(_0949_));
 sky130_fd_sc_hd__o21a_1 _5710_ (.A1(_0901_),
    .A2(_0949_),
    .B1(_0857_),
    .X(_0950_));
 sky130_fd_sc_hd__a21oi_1 _5711_ (.A1(_0795_),
    .A2(_0850_),
    .B1(_0853_),
    .Y(_0951_));
 sky130_fd_sc_hd__a21o_2 _5712_ (.A1(_0855_),
    .A2(_0950_),
    .B1(_0951_),
    .X(_0952_));
 sky130_fd_sc_hd__xnor2_4 _5713_ (.A(_0905_),
    .B(_0907_),
    .Y(_0953_));
 sky130_fd_sc_hd__and3_1 _5714_ (.A(_0273_),
    .B(net83),
    .C(_0743_),
    .X(_0954_));
 sky130_fd_sc_hd__or2_2 _5715_ (.A(net81),
    .B(net54),
    .X(_0955_));
 sky130_fd_sc_hd__xnor2_1 _5716_ (.A(_0904_),
    .B(_0955_),
    .Y(_0956_));
 sky130_fd_sc_hd__or3b_4 _5717_ (.A(net53),
    .B(net108),
    .C_N(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__a21bo_2 _5718_ (.A1(_0527_),
    .A2(_0954_),
    .B1_N(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__and2b_1 _5719_ (.A_N(_0953_),
    .B(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__xnor2_4 _5720_ (.A(_0953_),
    .B(_0958_),
    .Y(_0960_));
 sky130_fd_sc_hd__and2_2 _5721_ (.A(net48),
    .B(_0587_),
    .X(_0961_));
 sky130_fd_sc_hd__and3_2 _5722_ (.A(_0414_),
    .B(_0415_),
    .C(_0587_),
    .X(_0962_));
 sky130_fd_sc_hd__and3_4 _5723_ (.A(net48),
    .B(net73),
    .C(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__xnor2_4 _5724_ (.A(_0914_),
    .B(_0962_),
    .Y(_0964_));
 sky130_fd_sc_hd__a21o_2 _5725_ (.A1(_0960_),
    .A2(_0964_),
    .B1(_0959_),
    .X(_0965_));
 sky130_fd_sc_hd__xor2_4 _5726_ (.A(_0911_),
    .B(_0917_),
    .X(_0966_));
 sky130_fd_sc_hd__and2_1 _5727_ (.A(_0965_),
    .B(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__xor2_4 _5728_ (.A(_0965_),
    .B(_0966_),
    .X(_0968_));
 sky130_fd_sc_hd__a21oi_4 _5729_ (.A1(_0963_),
    .A2(_0968_),
    .B1(_0967_),
    .Y(_0969_));
 sky130_fd_sc_hd__xnor2_4 _5730_ (.A(_0921_),
    .B(_0924_),
    .Y(_0970_));
 sky130_fd_sc_hd__nor2_1 _5731_ (.A(_0969_),
    .B(_0970_),
    .Y(_0971_));
 sky130_fd_sc_hd__xor2_4 _5732_ (.A(_0969_),
    .B(_0970_),
    .X(_0972_));
 sky130_fd_sc_hd__o21ai_1 _5733_ (.A1(net81),
    .A2(net51),
    .B1(_0886_),
    .Y(_0973_));
 sky130_fd_sc_hd__nor2_1 _5734_ (.A(net78),
    .B(_0605_),
    .Y(_0974_));
 sky130_fd_sc_hd__nand2_1 _5735_ (.A(_0930_),
    .B(_0974_),
    .Y(_0975_));
 sky130_fd_sc_hd__and3_4 _5736_ (.A(_0886_),
    .B(_0930_),
    .C(_0974_),
    .X(_0976_));
 sky130_fd_sc_hd__a21boi_2 _5737_ (.A1(_0931_),
    .A2(_0973_),
    .B1_N(_0975_),
    .Y(_0977_));
 sky130_fd_sc_hd__nor2_4 _5738_ (.A(_0976_),
    .B(_0977_),
    .Y(_0978_));
 sky130_fd_sc_hd__a21o_4 _5739_ (.A1(_0972_),
    .A2(_0978_),
    .B1(_0971_),
    .X(_0980_));
 sky130_fd_sc_hd__xor2_4 _5740_ (.A(_0928_),
    .B(_0935_),
    .X(_0981_));
 sky130_fd_sc_hd__xor2_4 _5741_ (.A(_0980_),
    .B(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__a22o_4 _5742_ (.A1(_0980_),
    .A2(_0981_),
    .B1(_0982_),
    .B2(_0976_),
    .X(_0983_));
 sky130_fd_sc_hd__xnor2_4 _5743_ (.A(_0939_),
    .B(_0940_),
    .Y(_0984_));
 sky130_fd_sc_hd__and2b_1 _5744_ (.A_N(_0984_),
    .B(_0983_),
    .X(_0985_));
 sky130_fd_sc_hd__and3_4 _5745_ (.A(_3464_),
    .B(_0275_),
    .C(_0943_),
    .X(_0986_));
 sky130_fd_sc_hd__xnor2_4 _5746_ (.A(_0983_),
    .B(_0984_),
    .Y(_0987_));
 sky130_fd_sc_hd__and2_1 _5747_ (.A(_0986_),
    .B(_0987_),
    .X(_0988_));
 sky130_fd_sc_hd__xor2_2 _5748_ (.A(_0945_),
    .B(_0946_),
    .X(_0989_));
 sky130_fd_sc_hd__o21a_1 _5749_ (.A1(_0985_),
    .A2(_0988_),
    .B1(_0989_),
    .X(_0990_));
 sky130_fd_sc_hd__or3_1 _5750_ (.A(_0985_),
    .B(_0988_),
    .C(_0989_),
    .X(_0991_));
 sky130_fd_sc_hd__xnor2_4 _5751_ (.A(_0986_),
    .B(_0987_),
    .Y(_0992_));
 sky130_fd_sc_hd__o21bai_4 _5752_ (.A1(net53),
    .A2(net108),
    .B1_N(_0956_),
    .Y(_0993_));
 sky130_fd_sc_hd__nand2_2 _5753_ (.A(net80),
    .B(_0744_),
    .Y(_0994_));
 sky130_fd_sc_hd__or2_2 _5754_ (.A(_0955_),
    .B(_0994_),
    .X(_0995_));
 sky130_fd_sc_hd__or2_4 _5755_ (.A(net53),
    .B(net103),
    .X(_0996_));
 sky130_fd_sc_hd__o21ba_2 _5756_ (.A1(net78),
    .A2(net54),
    .B1_N(_0954_),
    .X(_0997_));
 sky130_fd_sc_hd__o21ba_2 _5757_ (.A1(_0955_),
    .A2(_0994_),
    .B1_N(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__o31ai_4 _5758_ (.A1(net53),
    .A2(net103),
    .A3(_0997_),
    .B1(_0995_),
    .Y(_0999_));
 sky130_fd_sc_hd__nand3_4 _5759_ (.A(_0957_),
    .B(_0993_),
    .C(_0999_),
    .Y(_1001_));
 sky130_fd_sc_hd__a21o_2 _5760_ (.A1(_0957_),
    .A2(_0993_),
    .B1(_0999_),
    .X(_1002_));
 sky130_fd_sc_hd__nand3_4 _5761_ (.A(_0961_),
    .B(_1001_),
    .C(_1002_),
    .Y(_1003_));
 sky130_fd_sc_hd__nand2_4 _5762_ (.A(_1001_),
    .B(_1003_),
    .Y(_1004_));
 sky130_fd_sc_hd__xnor2_4 _5763_ (.A(_0960_),
    .B(_0964_),
    .Y(_1005_));
 sky130_fd_sc_hd__nand2b_4 _5764_ (.A_N(_1005_),
    .B(_1004_),
    .Y(_1006_));
 sky130_fd_sc_hd__xor2_4 _5765_ (.A(_0963_),
    .B(_0968_),
    .X(_1007_));
 sky130_fd_sc_hd__nand2b_1 _5766_ (.A_N(_1006_),
    .B(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__xor2_4 _5767_ (.A(_1006_),
    .B(_1007_),
    .X(_1009_));
 sky130_fd_sc_hd__nor2_1 _5768_ (.A(net78),
    .B(net51),
    .Y(_1010_));
 sky130_fd_sc_hd__or2_1 _5769_ (.A(net74),
    .B(net49),
    .X(_1012_));
 sky130_fd_sc_hd__or3_2 _5770_ (.A(net78),
    .B(net51),
    .C(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__and2b_4 _5771_ (.A_N(_1013_),
    .B(_0975_),
    .X(_1014_));
 sky130_fd_sc_hd__o21ai_1 _5772_ (.A1(_0929_),
    .A2(_1010_),
    .B1(_0975_),
    .Y(_1015_));
 sky130_fd_sc_hd__a21oi_1 _5773_ (.A1(_1013_),
    .A2(_1015_),
    .B1(_1014_),
    .Y(_1016_));
 sky130_fd_sc_hd__inv_2 _5774_ (.A(_1016_),
    .Y(_1017_));
 sky130_fd_sc_hd__o21a_4 _5775_ (.A1(_1009_),
    .A2(_1017_),
    .B1(_1008_),
    .X(_1018_));
 sky130_fd_sc_hd__xnor2_4 _5776_ (.A(_0972_),
    .B(_0978_),
    .Y(_1019_));
 sky130_fd_sc_hd__xor2_4 _5777_ (.A(_1018_),
    .B(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__a2bb2o_4 _5778_ (.A1_N(_1018_),
    .A2_N(_1019_),
    .B1(_1020_),
    .B2(_1014_),
    .X(_1021_));
 sky130_fd_sc_hd__xor2_4 _5779_ (.A(_0976_),
    .B(_0982_),
    .X(_1023_));
 sky130_fd_sc_hd__nand2_1 _5780_ (.A(net65),
    .B(_0944_),
    .Y(_1024_));
 sky130_fd_sc_hd__xor2_2 _5781_ (.A(_1021_),
    .B(_1023_),
    .X(_1025_));
 sky130_fd_sc_hd__and3_1 _5782_ (.A(net65),
    .B(_0944_),
    .C(_1025_),
    .X(_1026_));
 sky130_fd_sc_hd__a21oi_4 _5783_ (.A1(_1021_),
    .A2(_1023_),
    .B1(_1026_),
    .Y(_1027_));
 sky130_fd_sc_hd__nor2_8 _5784_ (.A(_0992_),
    .B(_1027_),
    .Y(_1028_));
 sky130_fd_sc_hd__o21a_2 _5785_ (.A1(_0990_),
    .A2(_1028_),
    .B1(_0991_),
    .X(_1029_));
 sky130_fd_sc_hd__and2_2 _5786_ (.A(_0992_),
    .B(_1027_),
    .X(_1030_));
 sky130_fd_sc_hd__nor2_8 _5787_ (.A(_1028_),
    .B(_1030_),
    .Y(_1031_));
 sky130_fd_sc_hd__xor2_4 _5788_ (.A(_1004_),
    .B(_1005_),
    .X(_1032_));
 sky130_fd_sc_hd__a21o_1 _5789_ (.A1(_1001_),
    .A2(_1002_),
    .B1(_0961_),
    .X(_1034_));
 sky130_fd_sc_hd__xnor2_4 _5790_ (.A(_0996_),
    .B(_0998_),
    .Y(_1035_));
 sky130_fd_sc_hd__or2_2 _5791_ (.A(net74),
    .B(net54),
    .X(_1036_));
 sky130_fd_sc_hd__nor2_4 _5792_ (.A(_0994_),
    .B(_1036_),
    .Y(_1037_));
 sky130_fd_sc_hd__and2_2 _5793_ (.A(_1035_),
    .B(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__nand3_4 _5794_ (.A(_1003_),
    .B(_1034_),
    .C(_1038_),
    .Y(_1039_));
 sky130_fd_sc_hd__xor2_2 _5795_ (.A(_1032_),
    .B(_1039_),
    .X(_1040_));
 sky130_fd_sc_hd__nor2_1 _5796_ (.A(net74),
    .B(net51),
    .Y(_1041_));
 sky130_fd_sc_hd__or2_4 _5797_ (.A(net111),
    .B(net49),
    .X(_1042_));
 sky130_fd_sc_hd__and3b_4 _5798_ (.A_N(_1042_),
    .B(_1013_),
    .C(_1041_),
    .X(_1043_));
 sky130_fd_sc_hd__inv_2 _5799_ (.A(_1043_),
    .Y(_1045_));
 sky130_fd_sc_hd__or4_1 _5800_ (.A(net78),
    .B(net112),
    .C(net50),
    .D(_1012_),
    .X(_1046_));
 sky130_fd_sc_hd__o211a_1 _5801_ (.A1(_0974_),
    .A2(_1041_),
    .B1(_1045_),
    .C1(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__nand2_2 _5802_ (.A(_1040_),
    .B(_1047_),
    .Y(_1048_));
 sky130_fd_sc_hd__o21ai_4 _5803_ (.A1(_1032_),
    .A2(_1039_),
    .B1(_1048_),
    .Y(_1049_));
 sky130_fd_sc_hd__xnor2_4 _5804_ (.A(_1009_),
    .B(_1017_),
    .Y(_1050_));
 sky130_fd_sc_hd__nand2b_1 _5805_ (.A_N(_1050_),
    .B(_1049_),
    .Y(_1051_));
 sky130_fd_sc_hd__xnor2_4 _5806_ (.A(_1049_),
    .B(_1050_),
    .Y(_1052_));
 sky130_fd_sc_hd__a21boi_4 _5807_ (.A1(_1043_),
    .A2(_1052_),
    .B1_N(_1051_),
    .Y(_1053_));
 sky130_fd_sc_hd__xnor2_4 _5808_ (.A(_1014_),
    .B(_1020_),
    .Y(_1054_));
 sky130_fd_sc_hd__or2_1 _5809_ (.A(_1053_),
    .B(_1054_),
    .X(_1056_));
 sky130_fd_sc_hd__nand2_2 _5810_ (.A(net87),
    .B(_0944_),
    .Y(_1057_));
 sky130_fd_sc_hd__xor2_4 _5811_ (.A(_1053_),
    .B(_1054_),
    .X(_1058_));
 sky130_fd_sc_hd__nand2b_1 _5812_ (.A_N(_1057_),
    .B(_1058_),
    .Y(_1059_));
 sky130_fd_sc_hd__xor2_1 _5813_ (.A(_1024_),
    .B(_1025_),
    .X(_1060_));
 sky130_fd_sc_hd__a21o_1 _5814_ (.A1(_1056_),
    .A2(_1059_),
    .B1(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__and3_1 _5815_ (.A(_1056_),
    .B(_1059_),
    .C(_1060_),
    .X(_1062_));
 sky130_fd_sc_hd__inv_2 _5816_ (.A(_1062_),
    .Y(_1063_));
 sky130_fd_sc_hd__xor2_2 _5817_ (.A(_1057_),
    .B(_1058_),
    .X(_1064_));
 sky130_fd_sc_hd__a21o_1 _5818_ (.A1(_1003_),
    .A2(_1034_),
    .B1(_1038_),
    .X(_1065_));
 sky130_fd_sc_hd__nand2_1 _5819_ (.A(net112),
    .B(_0744_),
    .Y(_1067_));
 sky130_fd_sc_hd__or2_1 _5820_ (.A(net54),
    .B(net110),
    .X(_1068_));
 sky130_fd_sc_hd__or2_1 _5821_ (.A(_1036_),
    .B(_1067_),
    .X(_1069_));
 sky130_fd_sc_hd__and2_1 _5822_ (.A(_0994_),
    .B(_1036_),
    .X(_1070_));
 sky130_fd_sc_hd__or2_2 _5823_ (.A(_1037_),
    .B(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__xnor2_4 _5824_ (.A(_1035_),
    .B(_1037_),
    .Y(_1072_));
 sky130_fd_sc_hd__nor3_2 _5825_ (.A(_1069_),
    .B(_1071_),
    .C(_1072_),
    .Y(_1073_));
 sky130_fd_sc_hd__nand3_1 _5826_ (.A(_1039_),
    .B(_1065_),
    .C(_1073_),
    .Y(_1074_));
 sky130_fd_sc_hd__a21o_1 _5827_ (.A1(_1039_),
    .A2(_1065_),
    .B1(_1073_),
    .X(_1075_));
 sky130_fd_sc_hd__nor2_4 _5828_ (.A(net108),
    .B(net49),
    .Y(_1076_));
 sky130_fd_sc_hd__nor4_1 _5829_ (.A(net77),
    .B(net108),
    .C(net50),
    .D(_1042_),
    .Y(_1078_));
 sky130_fd_sc_hd__or4_4 _5830_ (.A(net76),
    .B(net108),
    .C(net50),
    .D(_1042_),
    .X(_1079_));
 sky130_fd_sc_hd__o21ai_1 _5831_ (.A1(net111),
    .A2(net50),
    .B1(_1012_),
    .Y(_1080_));
 sky130_fd_sc_hd__or4_1 _5832_ (.A(net74),
    .B(net73),
    .C(net50),
    .D(_1042_),
    .X(_1081_));
 sky130_fd_sc_hd__and3_1 _5833_ (.A(_1079_),
    .B(_1080_),
    .C(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__and3_2 _5834_ (.A(_1074_),
    .B(_1075_),
    .C(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__a31o_4 _5835_ (.A1(_1039_),
    .A2(_1065_),
    .A3(_1073_),
    .B1(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__or2_1 _5836_ (.A(_1040_),
    .B(_1047_),
    .X(_1085_));
 sky130_fd_sc_hd__nand2_2 _5837_ (.A(_1048_),
    .B(_1085_),
    .Y(_1086_));
 sky130_fd_sc_hd__xnor2_4 _5838_ (.A(_1084_),
    .B(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__a32o_2 _5839_ (.A1(_1048_),
    .A2(_1084_),
    .A3(_1085_),
    .B1(_1087_),
    .B2(_1078_),
    .X(_1089_));
 sky130_fd_sc_hd__xnor2_2 _5840_ (.A(_1043_),
    .B(_1052_),
    .Y(_1090_));
 sky130_fd_sc_hd__and2b_1 _5841_ (.A_N(_1090_),
    .B(_1089_),
    .X(_1091_));
 sky130_fd_sc_hd__and3_1 _5842_ (.A(_0275_),
    .B(_0364_),
    .C(_0943_),
    .X(_1092_));
 sky130_fd_sc_hd__xnor2_2 _5843_ (.A(_1089_),
    .B(_1090_),
    .Y(_1093_));
 sky130_fd_sc_hd__a21oi_2 _5844_ (.A1(_1092_),
    .A2(_1093_),
    .B1(_1091_),
    .Y(_1094_));
 sky130_fd_sc_hd__or2_1 _5845_ (.A(_1064_),
    .B(_1094_),
    .X(_1095_));
 sky130_fd_sc_hd__a21oi_1 _5846_ (.A1(_1061_),
    .A2(_1095_),
    .B1(_1062_),
    .Y(_1096_));
 sky130_fd_sc_hd__nand2_1 _5847_ (.A(_1061_),
    .B(_1063_),
    .Y(_1097_));
 sky130_fd_sc_hd__xnor2_1 _5848_ (.A(_1064_),
    .B(_1094_),
    .Y(_1098_));
 sky130_fd_sc_hd__inv_2 _5849_ (.A(_1098_),
    .Y(_1100_));
 sky130_fd_sc_hd__xnor2_1 _5850_ (.A(_1092_),
    .B(_1093_),
    .Y(_1101_));
 sky130_fd_sc_hd__xor2_4 _5851_ (.A(_1079_),
    .B(_1087_),
    .X(_1102_));
 sky130_fd_sc_hd__a21oi_2 _5852_ (.A1(_1074_),
    .A2(_1075_),
    .B1(_1082_),
    .Y(_1103_));
 sky130_fd_sc_hd__nor2_1 _5853_ (.A(net103),
    .B(net49),
    .Y(_1104_));
 sky130_fd_sc_hd__o211a_1 _5854_ (.A1(net111),
    .A2(net50),
    .B1(_0592_),
    .C1(_1076_),
    .X(_1105_));
 sky130_fd_sc_hd__or4_1 _5855_ (.A(net108),
    .B(net50),
    .C(_1042_),
    .D(_1104_),
    .X(_1106_));
 sky130_fd_sc_hd__o31ai_1 _5856_ (.A1(net108),
    .A2(net50),
    .A3(_1104_),
    .B1(_1042_),
    .Y(_1107_));
 sky130_fd_sc_hd__nand2_1 _5857_ (.A(_1106_),
    .B(_1107_),
    .Y(_1108_));
 sky130_fd_sc_hd__nand2_1 _5858_ (.A(net73),
    .B(_0744_),
    .Y(_1109_));
 sky130_fd_sc_hd__nor2_1 _5859_ (.A(_1068_),
    .B(_1109_),
    .Y(_1111_));
 sky130_fd_sc_hd__o21a_1 _5860_ (.A1(_1068_),
    .A2(_1109_),
    .B1(_1069_),
    .X(_1112_));
 sky130_fd_sc_hd__nor2_2 _5861_ (.A(_1071_),
    .B(_1112_),
    .Y(_1113_));
 sky130_fd_sc_hd__xnor2_2 _5862_ (.A(_1072_),
    .B(_1113_),
    .Y(_1114_));
 sky130_fd_sc_hd__nand2b_1 _5863_ (.A_N(_1108_),
    .B(_1114_),
    .Y(_1115_));
 sky130_fd_sc_hd__nand2_1 _5864_ (.A(net74),
    .B(_1111_),
    .Y(_1116_));
 sky130_fd_sc_hd__o31a_1 _5865_ (.A1(_1071_),
    .A2(_1072_),
    .A3(_1116_),
    .B1(_1115_),
    .X(_1117_));
 sky130_fd_sc_hd__or3_2 _5866_ (.A(_1083_),
    .B(_1103_),
    .C(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__o21ai_2 _5867_ (.A1(_1083_),
    .A2(_1103_),
    .B1(_1117_),
    .Y(_1119_));
 sky130_fd_sc_hd__nand3_2 _5868_ (.A(_1105_),
    .B(_1118_),
    .C(_1119_),
    .Y(_1120_));
 sky130_fd_sc_hd__and2_2 _5869_ (.A(_1118_),
    .B(_1120_),
    .X(_1122_));
 sky130_fd_sc_hd__nand2_1 _5870_ (.A(_0372_),
    .B(_0944_),
    .Y(_1123_));
 sky130_fd_sc_hd__xor2_2 _5871_ (.A(_1102_),
    .B(_1122_),
    .X(_1124_));
 sky130_fd_sc_hd__nand2b_1 _5872_ (.A_N(_1123_),
    .B(_1124_),
    .Y(_1125_));
 sky130_fd_sc_hd__o21a_1 _5873_ (.A1(_1102_),
    .A2(_1122_),
    .B1(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__nor2_1 _5874_ (.A(_1101_),
    .B(_1126_),
    .Y(_1127_));
 sky130_fd_sc_hd__nand2_1 _5875_ (.A(_1101_),
    .B(_1126_),
    .Y(_1128_));
 sky130_fd_sc_hd__nand2b_2 _5876_ (.A_N(_1127_),
    .B(_1128_),
    .Y(_1129_));
 sky130_fd_sc_hd__xor2_1 _5877_ (.A(_1123_),
    .B(_1124_),
    .X(_1130_));
 sky130_fd_sc_hd__a21o_1 _5878_ (.A1(_1118_),
    .A2(_1119_),
    .B1(_1105_),
    .X(_1131_));
 sky130_fd_sc_hd__xor2_1 _5879_ (.A(_1108_),
    .B(_1114_),
    .X(_1133_));
 sky130_fd_sc_hd__nor2_1 _5880_ (.A(net54),
    .B(net103),
    .Y(_1134_));
 sky130_fd_sc_hd__or4_2 _5881_ (.A(_0526_),
    .B(net112),
    .C(net102),
    .D(_1109_),
    .X(_1135_));
 sky130_fd_sc_hd__a21boi_1 _5882_ (.A1(net76),
    .A2(_0744_),
    .B1_N(_1068_),
    .Y(_1136_));
 sky130_fd_sc_hd__a21oi_1 _5883_ (.A1(net76),
    .A2(_1111_),
    .B1(_1112_),
    .Y(_1137_));
 sky130_fd_sc_hd__or3_4 _5884_ (.A(_1135_),
    .B(_1136_),
    .C(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__and2_1 _5885_ (.A(_1071_),
    .B(_1112_),
    .X(_1139_));
 sky130_fd_sc_hd__or2_4 _5886_ (.A(_1113_),
    .B(_1139_),
    .X(_1140_));
 sky130_fd_sc_hd__nor2_1 _5887_ (.A(_1138_),
    .B(_1140_),
    .Y(_1141_));
 sky130_fd_sc_hd__xor2_4 _5888_ (.A(_1138_),
    .B(_1140_),
    .X(_1142_));
 sky130_fd_sc_hd__xnor2_4 _5889_ (.A(_0591_),
    .B(_1076_),
    .Y(_1144_));
 sky130_fd_sc_hd__a21oi_1 _5890_ (.A1(_1142_),
    .A2(_1144_),
    .B1(_1141_),
    .Y(_1145_));
 sky130_fd_sc_hd__nor2_1 _5891_ (.A(_1133_),
    .B(_1145_),
    .Y(_1146_));
 sky130_fd_sc_hd__and3_1 _5892_ (.A(_1120_),
    .B(_1131_),
    .C(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__nand3_1 _5893_ (.A(_1120_),
    .B(_1131_),
    .C(_1146_),
    .Y(_1148_));
 sky130_fd_sc_hd__nand2_1 _5894_ (.A(net80),
    .B(_0944_),
    .Y(_1149_));
 sky130_fd_sc_hd__a21oi_1 _5895_ (.A1(_1120_),
    .A2(_1131_),
    .B1(_1146_),
    .Y(_1150_));
 sky130_fd_sc_hd__or3_2 _5896_ (.A(_1147_),
    .B(_1149_),
    .C(_1150_),
    .X(_1151_));
 sky130_fd_sc_hd__nand3_1 _5897_ (.A(_1130_),
    .B(_1148_),
    .C(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hd__a21o_1 _5898_ (.A1(_1148_),
    .A2(_1151_),
    .B1(_1130_),
    .X(_1153_));
 sky130_fd_sc_hd__o21ai_1 _5899_ (.A1(_1147_),
    .A2(_1150_),
    .B1(_1149_),
    .Y(_1155_));
 sky130_fd_sc_hd__and2_1 _5900_ (.A(_1133_),
    .B(_1145_),
    .X(_1156_));
 sky130_fd_sc_hd__or2_1 _5901_ (.A(_1146_),
    .B(_1156_),
    .X(_1157_));
 sky130_fd_sc_hd__xor2_2 _5902_ (.A(_1142_),
    .B(_1144_),
    .X(_1158_));
 sky130_fd_sc_hd__o21ai_1 _5903_ (.A1(_1136_),
    .A2(_1137_),
    .B1(_1135_),
    .Y(_1159_));
 sky130_fd_sc_hd__and2_1 _5904_ (.A(_1138_),
    .B(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__and2_1 _5905_ (.A(_1104_),
    .B(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__and2_1 _5906_ (.A(_1158_),
    .B(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__nand2_1 _5907_ (.A(_1158_),
    .B(_1161_),
    .Y(_1163_));
 sky130_fd_sc_hd__and3_1 _5908_ (.A(_0275_),
    .B(net77),
    .C(_0943_),
    .X(_1164_));
 sky130_fd_sc_hd__xnor2_1 _5909_ (.A(_1157_),
    .B(_1162_),
    .Y(_1166_));
 sky130_fd_sc_hd__nand2_1 _5910_ (.A(_1164_),
    .B(_1166_),
    .Y(_1167_));
 sky130_fd_sc_hd__o21ai_1 _5911_ (.A1(_1157_),
    .A2(_1163_),
    .B1(_1167_),
    .Y(_1168_));
 sky130_fd_sc_hd__and3_1 _5912_ (.A(_1151_),
    .B(_1155_),
    .C(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__a21oi_1 _5913_ (.A1(_1151_),
    .A2(_1155_),
    .B1(_1168_),
    .Y(_1170_));
 sky130_fd_sc_hd__nor2_1 _5914_ (.A(_1169_),
    .B(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__or2_1 _5915_ (.A(_1164_),
    .B(_1166_),
    .X(_1172_));
 sky130_fd_sc_hd__nand2_1 _5916_ (.A(_1167_),
    .B(_1172_),
    .Y(_1173_));
 sky130_fd_sc_hd__nor2_1 _5917_ (.A(_1158_),
    .B(_1161_),
    .Y(_1174_));
 sky130_fd_sc_hd__nor2_1 _5918_ (.A(_1162_),
    .B(_1174_),
    .Y(_1175_));
 sky130_fd_sc_hd__and3_1 _5919_ (.A(net112),
    .B(_0944_),
    .C(_1175_),
    .X(_1177_));
 sky130_fd_sc_hd__a21oi_1 _5920_ (.A1(net112),
    .A2(_0944_),
    .B1(_1175_),
    .Y(_1178_));
 sky130_fd_sc_hd__nor2_1 _5921_ (.A(_1104_),
    .B(_1160_),
    .Y(_1179_));
 sky130_fd_sc_hd__or2_1 _5922_ (.A(_1161_),
    .B(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__nand2_1 _5923_ (.A(_0548_),
    .B(_0944_),
    .Y(_1181_));
 sky130_fd_sc_hd__xor2_1 _5924_ (.A(_1180_),
    .B(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__nand2_1 _5925_ (.A(net103),
    .B(_1111_),
    .Y(_1183_));
 sky130_fd_sc_hd__o21ai_1 _5926_ (.A1(_0526_),
    .A2(net107),
    .B1(_1067_),
    .Y(_1184_));
 sky130_fd_sc_hd__and4_1 _5927_ (.A(_0587_),
    .B(_0944_),
    .C(_1135_),
    .D(_1184_),
    .X(_1185_));
 sky130_fd_sc_hd__and2_1 _5928_ (.A(_1182_),
    .B(_1185_),
    .X(_1186_));
 sky130_fd_sc_hd__o21ba_1 _5929_ (.A1(_1180_),
    .A2(_1181_),
    .B1_N(_1186_),
    .X(_1188_));
 sky130_fd_sc_hd__o21ba_1 _5930_ (.A1(_1178_),
    .A2(_1188_),
    .B1_N(_1177_),
    .X(_1189_));
 sky130_fd_sc_hd__nor2_1 _5931_ (.A(_1173_),
    .B(_1189_),
    .Y(_1190_));
 sky130_fd_sc_hd__a21o_1 _5932_ (.A1(_1171_),
    .A2(_1190_),
    .B1(_1169_),
    .X(_1191_));
 sky130_fd_sc_hd__and2b_1 _5933_ (.A_N(_1191_),
    .B(_1153_),
    .X(_1192_));
 sky130_fd_sc_hd__a21bo_1 _5934_ (.A1(_1152_),
    .A2(_1191_),
    .B1_N(_1153_),
    .X(_1193_));
 sky130_fd_sc_hd__a21o_4 _5935_ (.A1(_1128_),
    .A2(_1193_),
    .B1(_1127_),
    .X(_1194_));
 sky130_fd_sc_hd__nand2_1 _5936_ (.A(_1100_),
    .B(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__a41o_4 _5937_ (.A1(_1061_),
    .A2(_1063_),
    .A3(_1100_),
    .A4(_1194_),
    .B1(_1096_),
    .X(_1196_));
 sky130_fd_sc_hd__and2b_4 _5938_ (.A_N(_0990_),
    .B(_0991_),
    .X(_1197_));
 sky130_fd_sc_hd__a31oi_4 _5939_ (.A1(_1031_),
    .A2(_1196_),
    .A3(_1197_),
    .B1(_1029_),
    .Y(_1199_));
 sky130_fd_sc_hd__a31o_2 _5940_ (.A1(_1031_),
    .A2(_1196_),
    .A3(_1197_),
    .B1(_1029_),
    .X(_1200_));
 sky130_fd_sc_hd__and2b_1 _5941_ (.A_N(_0947_),
    .B(_0948_),
    .X(_1201_));
 sky130_fd_sc_hd__or2_4 _5942_ (.A(_0949_),
    .B(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__xnor2_4 _5943_ (.A(_0857_),
    .B(_0901_),
    .Y(_1203_));
 sky130_fd_sc_hd__nor2_2 _5944_ (.A(_1202_),
    .B(_1203_),
    .Y(_1204_));
 sky130_fd_sc_hd__a31oi_4 _5945_ (.A1(_0855_),
    .A2(_1200_),
    .A3(_1204_),
    .B1(_0952_),
    .Y(_1205_));
 sky130_fd_sc_hd__nand2b_1 _5946_ (.A_N(_0738_),
    .B(_0952_),
    .Y(_1206_));
 sky130_fd_sc_hd__or4bb_2 _5947_ (.A(_0738_),
    .B(_1199_),
    .C_N(_1204_),
    .D_N(_0855_),
    .X(_1207_));
 sky130_fd_sc_hd__o21ai_1 _5948_ (.A1(_0709_),
    .A2(_0713_),
    .B1(_0725_),
    .Y(_1208_));
 sky130_fd_sc_hd__a21o_1 _5949_ (.A1(_0729_),
    .A2(_0731_),
    .B1(_0733_),
    .X(_1210_));
 sky130_fd_sc_hd__o21a_1 _5950_ (.A1(_0736_),
    .A2(_1208_),
    .B1(_1210_),
    .X(_1211_));
 sky130_fd_sc_hd__and3_1 _5951_ (.A(_1206_),
    .B(_1207_),
    .C(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__a311o_2 _5952_ (.A1(_1206_),
    .A2(_1207_),
    .A3(_1211_),
    .B1(_0514_),
    .C1(_0464_),
    .X(_1213_));
 sky130_fd_sc_hd__a21bo_1 _5953_ (.A1(_0448_),
    .A2(_0512_),
    .B1_N(_0463_),
    .X(_1214_));
 sky130_fd_sc_hd__nor2_8 _5954_ (.A(net212),
    .B(net201),
    .Y(_1215_));
 sky130_fd_sc_hd__or2_4 _5955_ (.A(net212),
    .B(net201),
    .X(_1216_));
 sky130_fd_sc_hd__nand2_1 _5956_ (.A(_0389_),
    .B(_1215_),
    .Y(_1217_));
 sky130_fd_sc_hd__xor2_1 _5957_ (.A(_0451_),
    .B(_1217_),
    .X(_1218_));
 sky130_fd_sc_hd__a21o_1 _5958_ (.A1(_0455_),
    .A2(_0457_),
    .B1(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__nand3_1 _5959_ (.A(_0455_),
    .B(_0457_),
    .C(_1218_),
    .Y(_1221_));
 sky130_fd_sc_hd__nand2_2 _5960_ (.A(_1219_),
    .B(_1221_),
    .Y(_1222_));
 sky130_fd_sc_hd__xnor2_2 _5961_ (.A(_0461_),
    .B(_1222_),
    .Y(_1223_));
 sky130_fd_sc_hd__a21oi_1 _5962_ (.A1(_1213_),
    .A2(_1214_),
    .B1(_1223_),
    .Y(_1224_));
 sky130_fd_sc_hd__a21o_1 _5963_ (.A1(_1213_),
    .A2(_1214_),
    .B1(_1223_),
    .X(_1225_));
 sky130_fd_sc_hd__o211a_1 _5964_ (.A1(_0452_),
    .A2(_1216_),
    .B1(_1219_),
    .C1(_0389_),
    .X(_1226_));
 sky130_fd_sc_hd__o21a_1 _5965_ (.A1(_0461_),
    .A2(_1222_),
    .B1(_1226_),
    .X(_1227_));
 sky130_fd_sc_hd__and2_4 _5966_ (.A(_1225_),
    .B(_1227_),
    .X(_1228_));
 sky130_fd_sc_hd__and4_2 _5967_ (.A(net127),
    .B(net134),
    .C(net123),
    .D(net175),
    .X(_1229_));
 sky130_fd_sc_hd__and3b_4 _5968_ (.A_N(_3515_),
    .B(_3562_),
    .C(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__nand3b_4 _5969_ (.A_N(_3515_),
    .B(_3562_),
    .C(_1229_),
    .Y(_1232_));
 sky130_fd_sc_hd__and3_4 _5970_ (.A(_1225_),
    .B(_1227_),
    .C(net101),
    .X(_1233_));
 sky130_fd_sc_hd__nand2_2 _5971_ (.A(_1228_),
    .B(net101),
    .Y(_1234_));
 sky130_fd_sc_hd__nor2_1 _5972_ (.A(_3446_),
    .B(_1233_),
    .Y(_1235_));
 sky130_fd_sc_hd__a21oi_4 _5973_ (.A1(_0357_),
    .A2(_0358_),
    .B1(net169),
    .Y(_1236_));
 sky130_fd_sc_hd__o211a_1 _5974_ (.A1(_1209_),
    .A2(_1891_),
    .B1(_2056_),
    .C1(net131),
    .X(_1237_));
 sky130_fd_sc_hd__o211a_1 _5975_ (.A1(_1121_),
    .A2(_1891_),
    .B1(_2001_),
    .C1(net133),
    .X(_1238_));
 sky130_fd_sc_hd__o31ai_4 _5976_ (.A1(_1715_),
    .A2(_1237_),
    .A3(_1238_),
    .B1(net171),
    .Y(_1239_));
 sky130_fd_sc_hd__nand4_4 _5977_ (.A(net173),
    .B(net167),
    .C(_0360_),
    .D(_0361_),
    .Y(_1240_));
 sky130_fd_sc_hd__o21ai_4 _5978_ (.A1(_1236_),
    .A2(_1239_),
    .B1(_1240_),
    .Y(_1241_));
 sky130_fd_sc_hd__xnor2_4 _5979_ (.A(_3445_),
    .B(_1233_),
    .Y(_1243_));
 sky130_fd_sc_hd__a21oi_4 _5980_ (.A1(_1241_),
    .A2(_1243_),
    .B1(_1235_),
    .Y(_1244_));
 sky130_fd_sc_hd__a211o_1 _5981_ (.A1(_1242_),
    .A2(net129),
    .B1(_3452_),
    .C1(net131),
    .X(_1245_));
 sky130_fd_sc_hd__o21a_1 _5982_ (.A1(_1407_),
    .A2(net133),
    .B1(net169),
    .X(_1246_));
 sky130_fd_sc_hd__a32oi_4 _5983_ (.A1(_1715_),
    .A2(_0306_),
    .A3(_0307_),
    .B1(_1245_),
    .B2(_1246_),
    .Y(_1247_));
 sky130_fd_sc_hd__nand2_1 _5984_ (.A(net171),
    .B(_1247_),
    .Y(_1248_));
 sky130_fd_sc_hd__o21a_2 _5985_ (.A1(net171),
    .A2(_0496_),
    .B1(_1248_),
    .X(_1249_));
 sky130_fd_sc_hd__mux2_8 _5986_ (.A0(_0495_),
    .A1(_1247_),
    .S(net171),
    .X(_1250_));
 sky130_fd_sc_hd__xnor2_4 _5987_ (.A(_3434_),
    .B(_1244_),
    .Y(_1251_));
 sky130_fd_sc_hd__a2bb2o_4 _5988_ (.A1_N(_3435_),
    .A2_N(_1244_),
    .B1(_1249_),
    .B2(_1251_),
    .X(_1252_));
 sky130_fd_sc_hd__xnor2_4 _5989_ (.A(_2221_),
    .B(net190),
    .Y(_1254_));
 sky130_fd_sc_hd__xnor2_2 _5990_ (.A(net216),
    .B(net190),
    .Y(_1255_));
 sky130_fd_sc_hd__a211o_2 _5991_ (.A1(_1363_),
    .A2(_1880_),
    .B1(net205),
    .C1(_1319_),
    .X(_1256_));
 sky130_fd_sc_hd__inv_2 _5992_ (.A(_1256_),
    .Y(_1257_));
 sky130_fd_sc_hd__nand2_2 _5993_ (.A(net203),
    .B(net129),
    .Y(_1258_));
 sky130_fd_sc_hd__and2_4 _5994_ (.A(_1256_),
    .B(_1258_),
    .X(_1259_));
 sky130_fd_sc_hd__nand2_1 _5995_ (.A(_1256_),
    .B(_1258_),
    .Y(_1260_));
 sky130_fd_sc_hd__nor2_2 _5996_ (.A(_1255_),
    .B(_1260_),
    .Y(_1261_));
 sky130_fd_sc_hd__nand2_1 _5997_ (.A(_1254_),
    .B(_1259_),
    .Y(_1262_));
 sky130_fd_sc_hd__nor2_4 _5998_ (.A(_1254_),
    .B(_1259_),
    .Y(_1263_));
 sky130_fd_sc_hd__nor2_4 _5999_ (.A(_1261_),
    .B(_1263_),
    .Y(_1265_));
 sky130_fd_sc_hd__or2_4 _6000_ (.A(_1261_),
    .B(_1263_),
    .X(_1266_));
 sky130_fd_sc_hd__and2_1 _6001_ (.A(_2100_),
    .B(_3384_),
    .X(_1267_));
 sky130_fd_sc_hd__a211o_4 _6002_ (.A1(_3394_),
    .A2(_1252_),
    .B1(_1265_),
    .C1(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__a21oi_2 _6003_ (.A1(_3394_),
    .A2(_1252_),
    .B1(_1267_),
    .Y(_1269_));
 sky130_fd_sc_hd__o21a_4 _6004_ (.A1(_1266_),
    .A2(_1269_),
    .B1(_1268_),
    .X(_1270_));
 sky130_fd_sc_hd__nand2b_1 _6005_ (.A_N(_2100_),
    .B(_3384_),
    .Y(_1271_));
 sky130_fd_sc_hd__and2b_2 _6006_ (.A_N(_3384_),
    .B(_2100_),
    .X(_1272_));
 sky130_fd_sc_hd__xor2_4 _6007_ (.A(_2100_),
    .B(_3384_),
    .X(_1273_));
 sky130_fd_sc_hd__xnor2_1 _6008_ (.A(_1252_),
    .B(_1273_),
    .Y(_1274_));
 sky130_fd_sc_hd__xor2_4 _6009_ (.A(_1252_),
    .B(_1273_),
    .X(_1276_));
 sky130_fd_sc_hd__xor2_4 _6010_ (.A(_1241_),
    .B(_1243_),
    .X(_1277_));
 sky130_fd_sc_hd__xnor2_4 _6011_ (.A(_1250_),
    .B(_1251_),
    .Y(_1278_));
 sky130_fd_sc_hd__nor2_1 _6012_ (.A(_1277_),
    .B(_1278_),
    .Y(_1279_));
 sky130_fd_sc_hd__o2111a_4 _6013_ (.A1(_1266_),
    .A2(_1269_),
    .B1(_1274_),
    .C1(_1279_),
    .D1(_1268_),
    .X(_1280_));
 sky130_fd_sc_hd__nor2_2 _6014_ (.A(_2221_),
    .B(net212),
    .Y(_1281_));
 sky130_fd_sc_hd__or3_4 _6015_ (.A(_1088_),
    .B(net201),
    .C(_1281_),
    .X(_1282_));
 sky130_fd_sc_hd__clkinv_4 _6016_ (.A(_1282_),
    .Y(_1283_));
 sky130_fd_sc_hd__xnor2_2 _6017_ (.A(net192),
    .B(_1254_),
    .Y(_1284_));
 sky130_fd_sc_hd__nand2_4 _6018_ (.A(_1770_),
    .B(_1257_),
    .Y(_1285_));
 sky130_fd_sc_hd__o21a_2 _6019_ (.A1(net132),
    .A2(_1257_),
    .B1(_1285_),
    .X(_1287_));
 sky130_fd_sc_hd__inv_2 _6020_ (.A(_1287_),
    .Y(_1288_));
 sky130_fd_sc_hd__mux2_1 _6021_ (.A0(net132),
    .A1(_1288_),
    .S(_1258_),
    .X(_1289_));
 sky130_fd_sc_hd__and2b_1 _6022_ (.A_N(_1284_),
    .B(_1289_),
    .X(_1290_));
 sky130_fd_sc_hd__or2_4 _6023_ (.A(_1284_),
    .B(_1289_),
    .X(_1291_));
 sky130_fd_sc_hd__nand2_1 _6024_ (.A(_1284_),
    .B(_1289_),
    .Y(_1292_));
 sky130_fd_sc_hd__and2_4 _6025_ (.A(_1291_),
    .B(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__a21o_2 _6026_ (.A1(_1255_),
    .A2(_1259_),
    .B1(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__nand2_1 _6027_ (.A(_1259_),
    .B(_1293_),
    .Y(_1295_));
 sky130_fd_sc_hd__o21a_4 _6028_ (.A1(_1254_),
    .A2(_1295_),
    .B1(_1294_),
    .X(_1296_));
 sky130_fd_sc_hd__a21o_2 _6029_ (.A1(_1770_),
    .A2(_1891_),
    .B1(_1088_),
    .X(_1298_));
 sky130_fd_sc_hd__xnor2_4 _6030_ (.A(_1726_),
    .B(_1285_),
    .Y(_1299_));
 sky130_fd_sc_hd__xnor2_2 _6031_ (.A(_1298_),
    .B(_1299_),
    .Y(_1300_));
 sky130_fd_sc_hd__nand2_1 _6032_ (.A(net216),
    .B(_3403_),
    .Y(_1301_));
 sky130_fd_sc_hd__or2_4 _6033_ (.A(net216),
    .B(_3403_),
    .X(_1302_));
 sky130_fd_sc_hd__xnor2_4 _6034_ (.A(_2859_),
    .B(_1302_),
    .Y(_1303_));
 sky130_fd_sc_hd__mux2_2 _6035_ (.A0(net197),
    .A1(_1303_),
    .S(_1301_),
    .X(_1304_));
 sky130_fd_sc_hd__nor2_2 _6036_ (.A(_1300_),
    .B(_1304_),
    .Y(_1305_));
 sky130_fd_sc_hd__and2_1 _6037_ (.A(_1300_),
    .B(_1304_),
    .X(_1306_));
 sky130_fd_sc_hd__and2b_1 _6038_ (.A_N(_1304_),
    .B(_1300_),
    .X(_1307_));
 sky130_fd_sc_hd__nor2_4 _6039_ (.A(_1305_),
    .B(_1306_),
    .Y(_1309_));
 sky130_fd_sc_hd__inv_2 _6040_ (.A(_1309_),
    .Y(_1310_));
 sky130_fd_sc_hd__nand2_2 _6041_ (.A(_1291_),
    .B(_1309_),
    .Y(_1311_));
 sky130_fd_sc_hd__inv_2 _6042_ (.A(_1311_),
    .Y(_1312_));
 sky130_fd_sc_hd__nor2_4 _6043_ (.A(_1291_),
    .B(_1309_),
    .Y(_1313_));
 sky130_fd_sc_hd__nor2_4 _6044_ (.A(_1312_),
    .B(_1313_),
    .Y(_1314_));
 sky130_fd_sc_hd__and2_4 _6045_ (.A(_1296_),
    .B(_1314_),
    .X(_1315_));
 sky130_fd_sc_hd__a31o_1 _6046_ (.A1(_2859_),
    .A2(net192),
    .A3(net188),
    .B1(_2221_),
    .X(_1316_));
 sky130_fd_sc_hd__a21o_2 _6047_ (.A1(_2221_),
    .A2(_2617_),
    .B1(net185),
    .X(_1317_));
 sky130_fd_sc_hd__mux2_2 _6048_ (.A0(net187),
    .A1(_1317_),
    .S(_1316_),
    .X(_1318_));
 sky130_fd_sc_hd__a21o_1 _6049_ (.A1(_1298_),
    .A2(_1299_),
    .B1(_1088_),
    .X(_1320_));
 sky130_fd_sc_hd__o21ai_2 _6050_ (.A1(net204),
    .A2(_1561_),
    .B1(_1451_),
    .Y(_1321_));
 sky130_fd_sc_hd__mux2_1 _6051_ (.A0(_1451_),
    .A1(_1321_),
    .S(_1320_),
    .X(_1322_));
 sky130_fd_sc_hd__and2b_1 _6052_ (.A_N(_1318_),
    .B(_1322_),
    .X(_1323_));
 sky130_fd_sc_hd__nor2_1 _6053_ (.A(_1318_),
    .B(_1322_),
    .Y(_1324_));
 sky130_fd_sc_hd__and2_1 _6054_ (.A(_1318_),
    .B(_1322_),
    .X(_1325_));
 sky130_fd_sc_hd__or2_4 _6055_ (.A(_1324_),
    .B(_1325_),
    .X(_1326_));
 sky130_fd_sc_hd__clkinv_4 _6056_ (.A(_1326_),
    .Y(_1327_));
 sky130_fd_sc_hd__nor2_1 _6057_ (.A(_1307_),
    .B(_1326_),
    .Y(_1328_));
 sky130_fd_sc_hd__and2_1 _6058_ (.A(_1307_),
    .B(_1326_),
    .X(_1329_));
 sky130_fd_sc_hd__or2_4 _6059_ (.A(_1328_),
    .B(_1329_),
    .X(_1331_));
 sky130_fd_sc_hd__nor2_2 _6060_ (.A(_1088_),
    .B(_2221_),
    .Y(_1332_));
 sky130_fd_sc_hd__nand2_4 _6061_ (.A(net205),
    .B(net216),
    .Y(_1333_));
 sky130_fd_sc_hd__nor2_1 _6062_ (.A(_1216_),
    .B(_1333_),
    .Y(_1334_));
 sky130_fd_sc_hd__a21oi_4 _6063_ (.A1(net204),
    .A2(net199),
    .B1(_1281_),
    .Y(_1335_));
 sky130_fd_sc_hd__nor2_2 _6064_ (.A(_1334_),
    .B(_1335_),
    .Y(_1336_));
 sky130_fd_sc_hd__or2_2 _6065_ (.A(_1334_),
    .B(_1335_),
    .X(_1337_));
 sky130_fd_sc_hd__or2_2 _6066_ (.A(_1323_),
    .B(_1337_),
    .X(_1338_));
 sky130_fd_sc_hd__nand2_2 _6067_ (.A(_1323_),
    .B(_1337_),
    .Y(_1339_));
 sky130_fd_sc_hd__nand2_4 _6068_ (.A(_1338_),
    .B(_1339_),
    .Y(_1340_));
 sky130_fd_sc_hd__nor2_2 _6069_ (.A(_1331_),
    .B(_1340_),
    .Y(_1342_));
 sky130_fd_sc_hd__a21oi_4 _6070_ (.A1(_1294_),
    .A2(_1311_),
    .B1(_1313_),
    .Y(_1343_));
 sky130_fd_sc_hd__inv_2 _6071_ (.A(_1343_),
    .Y(_1344_));
 sky130_fd_sc_hd__o21ai_1 _6072_ (.A1(_1329_),
    .A2(_1344_),
    .B1(_1338_),
    .Y(_1345_));
 sky130_fd_sc_hd__o21a_2 _6073_ (.A1(_1328_),
    .A2(_1345_),
    .B1(_1339_),
    .X(_1346_));
 sky130_fd_sc_hd__a31oi_4 _6074_ (.A1(_1268_),
    .A2(_1315_),
    .A3(_1342_),
    .B1(_1346_),
    .Y(_1347_));
 sky130_fd_sc_hd__a31o_4 _6075_ (.A1(_1268_),
    .A2(_1315_),
    .A3(_1342_),
    .B1(_1346_),
    .X(_1348_));
 sky130_fd_sc_hd__nor2_4 _6076_ (.A(_1283_),
    .B(_1347_),
    .Y(_1349_));
 sky130_fd_sc_hd__nand2_8 _6077_ (.A(_1282_),
    .B(_1348_),
    .Y(_1350_));
 sky130_fd_sc_hd__or3_4 _6078_ (.A(_1270_),
    .B(_1283_),
    .C(_1347_),
    .X(_1351_));
 sky130_fd_sc_hd__o21ai_4 _6079_ (.A1(_1283_),
    .A2(_1347_),
    .B1(_1270_),
    .Y(_1353_));
 sky130_fd_sc_hd__and2_1 _6080_ (.A(_1351_),
    .B(_1353_),
    .X(_1354_));
 sky130_fd_sc_hd__nand2_4 _6081_ (.A(_1351_),
    .B(_1353_),
    .Y(_1355_));
 sky130_fd_sc_hd__a21o_4 _6082_ (.A1(_1351_),
    .A2(_1353_),
    .B1(_1280_),
    .X(_1356_));
 sky130_fd_sc_hd__a21oi_4 _6083_ (.A1(_1282_),
    .A2(_1348_),
    .B1(_1280_),
    .Y(_1357_));
 sky130_fd_sc_hd__xor2_4 _6084_ (.A(_1268_),
    .B(_1296_),
    .X(_1358_));
 sky130_fd_sc_hd__xor2_4 _6085_ (.A(_1357_),
    .B(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__xnor2_4 _6086_ (.A(_1357_),
    .B(_1358_),
    .Y(_1360_));
 sky130_fd_sc_hd__nor2_2 _6087_ (.A(_1356_),
    .B(_1360_),
    .Y(_1361_));
 sky130_fd_sc_hd__nand2_2 _6088_ (.A(_1280_),
    .B(_1296_),
    .Y(_1362_));
 sky130_fd_sc_hd__o2bb2a_4 _6089_ (.A1_N(_1280_),
    .A2_N(_1296_),
    .B1(_1347_),
    .B2(_1283_),
    .X(_1364_));
 sky130_fd_sc_hd__a21boi_4 _6090_ (.A1(_1268_),
    .A2(_1296_),
    .B1_N(_1294_),
    .Y(_1365_));
 sky130_fd_sc_hd__xnor2_4 _6091_ (.A(_1314_),
    .B(_1365_),
    .Y(_1366_));
 sky130_fd_sc_hd__xnor2_4 _6092_ (.A(_1364_),
    .B(_1366_),
    .Y(_1367_));
 sky130_fd_sc_hd__or3_1 _6093_ (.A(_1356_),
    .B(_1360_),
    .C(_1367_),
    .X(_1368_));
 sky130_fd_sc_hd__a21oi_4 _6094_ (.A1(_1268_),
    .A2(_1315_),
    .B1(_1343_),
    .Y(_1369_));
 sky130_fd_sc_hd__xor2_4 _6095_ (.A(_1331_),
    .B(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__xnor2_4 _6096_ (.A(_1331_),
    .B(_1369_),
    .Y(_1371_));
 sky130_fd_sc_hd__o211ai_4 _6097_ (.A1(_1362_),
    .A2(_1366_),
    .B1(_1371_),
    .C1(_1350_),
    .Y(_1372_));
 sky130_fd_sc_hd__a211o_4 _6098_ (.A1(_1350_),
    .A2(_1366_),
    .B1(_1371_),
    .C1(_1364_),
    .X(_1373_));
 sky130_fd_sc_hd__nand2_1 _6099_ (.A(_1372_),
    .B(_1373_),
    .Y(_1375_));
 sky130_fd_sc_hd__o31a_4 _6100_ (.A1(_1362_),
    .A2(_1366_),
    .A3(_1370_),
    .B1(_1350_),
    .X(_1376_));
 sky130_fd_sc_hd__o21ba_2 _6101_ (.A1(_1329_),
    .A2(_1369_),
    .B1_N(_1328_),
    .X(_1377_));
 sky130_fd_sc_hd__xnor2_4 _6102_ (.A(_1340_),
    .B(_1377_),
    .Y(_1378_));
 sky130_fd_sc_hd__xor2_4 _6103_ (.A(_1376_),
    .B(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__xnor2_4 _6104_ (.A(_1376_),
    .B(_1378_),
    .Y(_1380_));
 sky130_fd_sc_hd__a2111oi_4 _6105_ (.A1(_1372_),
    .A2(_1373_),
    .B1(_1356_),
    .C1(_1360_),
    .D1(_1367_),
    .Y(_1381_));
 sky130_fd_sc_hd__a2111o_4 _6106_ (.A1(_1372_),
    .A2(_1373_),
    .B1(_1356_),
    .C1(_1360_),
    .D1(_1367_),
    .X(_1382_));
 sky130_fd_sc_hd__or3b_1 _6107_ (.A(_1375_),
    .B(_1380_),
    .C_N(_1368_),
    .X(_1383_));
 sky130_fd_sc_hd__clkinv_8 _6108_ (.A(net14),
    .Y(_1384_));
 sky130_fd_sc_hd__nand2_4 _6109_ (.A(_1379_),
    .B(_1382_),
    .Y(_1386_));
 sky130_fd_sc_hd__xnor2_2 _6110_ (.A(_1356_),
    .B(_1359_),
    .Y(_1387_));
 sky130_fd_sc_hd__and3b_2 _6111_ (.A_N(_1387_),
    .B(_1379_),
    .C(_1382_),
    .X(_1388_));
 sky130_fd_sc_hd__or3_1 _6112_ (.A(_1380_),
    .B(_1381_),
    .C(_1387_),
    .X(_1389_));
 sky130_fd_sc_hd__or3_2 _6113_ (.A(_1354_),
    .B(_1380_),
    .C(_1381_),
    .X(_1390_));
 sky130_fd_sc_hd__o21bai_4 _6114_ (.A1(_1199_),
    .A2(_1202_),
    .B1_N(_0949_),
    .Y(_1391_));
 sky130_fd_sc_hd__xor2_4 _6115_ (.A(_1203_),
    .B(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__a21oi_2 _6116_ (.A1(_1200_),
    .A2(_1204_),
    .B1(_0950_),
    .Y(_1393_));
 sky130_fd_sc_hd__or2_1 _6117_ (.A(_0851_),
    .B(_1393_),
    .X(_1394_));
 sky130_fd_sc_hd__nand2_1 _6118_ (.A(_0851_),
    .B(_1393_),
    .Y(_1395_));
 sky130_fd_sc_hd__a21oi_2 _6119_ (.A1(_1394_),
    .A2(_1395_),
    .B1(_1230_),
    .Y(_1397_));
 sky130_fd_sc_hd__and2b_1 _6120_ (.A_N(_1228_),
    .B(_1397_),
    .X(_1398_));
 sky130_fd_sc_hd__a221oi_4 _6121_ (.A1(net109),
    .A2(_1230_),
    .B1(_1233_),
    .B2(_1392_),
    .C1(_1398_),
    .Y(_1399_));
 sky130_fd_sc_hd__o21ai_1 _6122_ (.A1(_0851_),
    .A2(_1393_),
    .B1(_0850_),
    .Y(_1400_));
 sky130_fd_sc_hd__nand2_1 _6123_ (.A(_0854_),
    .B(_1400_),
    .Y(_1401_));
 sky130_fd_sc_hd__o211a_1 _6124_ (.A1(_0854_),
    .A2(_1400_),
    .B1(_1401_),
    .C1(net101),
    .X(_1402_));
 sky130_fd_sc_hd__mux2_1 _6125_ (.A0(_1402_),
    .A1(_1397_),
    .S(_1228_),
    .X(_1403_));
 sky130_fd_sc_hd__or2_4 _6126_ (.A(_1228_),
    .B(_1230_),
    .X(_1404_));
 sky130_fd_sc_hd__clkinv_4 _6127_ (.A(_1404_),
    .Y(_1405_));
 sky130_fd_sc_hd__a21oi_2 _6128_ (.A1(net111),
    .A2(_1230_),
    .B1(_1403_),
    .Y(_1406_));
 sky130_fd_sc_hd__a31o_1 _6129_ (.A1(_1355_),
    .A2(_1379_),
    .A3(_1382_),
    .B1(_1406_),
    .X(_1408_));
 sky130_fd_sc_hd__o21ai_1 _6130_ (.A1(net9),
    .A2(_1399_),
    .B1(_1408_),
    .Y(_1409_));
 sky130_fd_sc_hd__o21a_1 _6131_ (.A1(net9),
    .A2(_1399_),
    .B1(_1408_),
    .X(_1410_));
 sky130_fd_sc_hd__xnor2_4 _6132_ (.A(_1361_),
    .B(_1367_),
    .Y(_1411_));
 sky130_fd_sc_hd__nor2_8 _6133_ (.A(_1386_),
    .B(_1411_),
    .Y(_1412_));
 sky130_fd_sc_hd__or2_1 _6134_ (.A(_1386_),
    .B(_1411_),
    .X(_1413_));
 sky130_fd_sc_hd__xnor2_4 _6135_ (.A(_1199_),
    .B(_1202_),
    .Y(_1414_));
 sky130_fd_sc_hd__a21oi_4 _6136_ (.A1(_1031_),
    .A2(_1196_),
    .B1(_1028_),
    .Y(_1415_));
 sky130_fd_sc_hd__xor2_4 _6137_ (.A(_1197_),
    .B(_1415_),
    .X(_1416_));
 sky130_fd_sc_hd__o22ai_2 _6138_ (.A1(_1404_),
    .A2(_1414_),
    .B1(_1416_),
    .B2(_1234_),
    .Y(_1417_));
 sky130_fd_sc_hd__nor2_2 _6139_ (.A(_0587_),
    .B(net101),
    .Y(_1419_));
 sky130_fd_sc_hd__a221oi_4 _6140_ (.A1(_1392_),
    .A2(_1405_),
    .B1(_1414_),
    .B2(_1233_),
    .C1(_1419_),
    .Y(_1420_));
 sky130_fd_sc_hd__mux2_1 _6141_ (.A0(_1417_),
    .A1(_1420_),
    .S(net10),
    .X(_1421_));
 sky130_fd_sc_hd__mux2_1 _6142_ (.A0(_1410_),
    .A1(_1421_),
    .S(net13),
    .X(_1422_));
 sky130_fd_sc_hd__nor2_2 _6143_ (.A(_0714_),
    .B(_1205_),
    .Y(_1423_));
 sky130_fd_sc_hd__and2_1 _6144_ (.A(_0714_),
    .B(_1205_),
    .X(_1424_));
 sky130_fd_sc_hd__nor2_1 _6145_ (.A(_1423_),
    .B(_1424_),
    .Y(_1425_));
 sky130_fd_sc_hd__or2_1 _6146_ (.A(_1234_),
    .B(_1425_),
    .X(_1426_));
 sky130_fd_sc_hd__nor2_1 _6147_ (.A(_0713_),
    .B(_1423_),
    .Y(_1427_));
 sky130_fd_sc_hd__xnor2_2 _6148_ (.A(_0726_),
    .B(_1427_),
    .Y(_1428_));
 sky130_fd_sc_hd__o221a_2 _6149_ (.A1(_0430_),
    .A2(net101),
    .B1(_1404_),
    .B2(_1428_),
    .C1(_1426_),
    .X(_1430_));
 sky130_fd_sc_hd__nand2_1 _6150_ (.A(_1228_),
    .B(_1402_),
    .Y(_1431_));
 sky130_fd_sc_hd__o221a_1 _6151_ (.A1(net77),
    .A2(net101),
    .B1(_1404_),
    .B2(_1425_),
    .C1(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__a31o_1 _6152_ (.A1(_1355_),
    .A2(_1379_),
    .A3(_1382_),
    .B1(_1430_),
    .X(_1433_));
 sky130_fd_sc_hd__o21ai_1 _6153_ (.A1(net9),
    .A2(_1432_),
    .B1(_1433_),
    .Y(_1434_));
 sky130_fd_sc_hd__a21boi_2 _6154_ (.A1(_0726_),
    .A2(_1423_),
    .B1_N(_1208_),
    .Y(_1435_));
 sky130_fd_sc_hd__xnor2_1 _6155_ (.A(_0732_),
    .B(_1435_),
    .Y(_1436_));
 sky130_fd_sc_hd__nand2_1 _6156_ (.A(_1405_),
    .B(_1436_),
    .Y(_1437_));
 sky130_fd_sc_hd__o221a_1 _6157_ (.A1(net83),
    .A2(_1232_),
    .B1(_1234_),
    .B2(_1428_),
    .C1(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__o21a_2 _6158_ (.A1(_0732_),
    .A2(_1435_),
    .B1(_0731_),
    .X(_1439_));
 sky130_fd_sc_hd__xnor2_4 _6159_ (.A(_0735_),
    .B(_1439_),
    .Y(_1441_));
 sky130_fd_sc_hd__and2_1 _6160_ (.A(_1233_),
    .B(_1436_),
    .X(_1442_));
 sky130_fd_sc_hd__a221oi_4 _6161_ (.A1(net86),
    .A2(_1230_),
    .B1(_1405_),
    .B2(_1441_),
    .C1(_1442_),
    .Y(_1443_));
 sky130_fd_sc_hd__a31o_1 _6162_ (.A1(_1355_),
    .A2(_1379_),
    .A3(_1382_),
    .B1(_1443_),
    .X(_1444_));
 sky130_fd_sc_hd__or4_1 _6163_ (.A(_1354_),
    .B(_1380_),
    .C(_1381_),
    .D(_1438_),
    .X(_1445_));
 sky130_fd_sc_hd__a21oi_1 _6164_ (.A1(_1444_),
    .A2(_1445_),
    .B1(net13),
    .Y(_1446_));
 sky130_fd_sc_hd__a21oi_1 _6165_ (.A1(net13),
    .A2(_1434_),
    .B1(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__mux2_2 _6166_ (.A0(_1422_),
    .A1(_1447_),
    .S(net8),
    .X(_1448_));
 sky130_fd_sc_hd__a31o_1 _6167_ (.A1(_1355_),
    .A2(_1379_),
    .A3(_1382_),
    .B1(_1276_),
    .X(_1449_));
 sky130_fd_sc_hd__o21a_1 _6168_ (.A1(_1278_),
    .A2(net10),
    .B1(_1449_),
    .X(_1450_));
 sky130_fd_sc_hd__a2bb2o_1 _6169_ (.A1_N(_1353_),
    .A2_N(_1386_),
    .B1(net10),
    .B2(_1349_),
    .X(_1452_));
 sky130_fd_sc_hd__mux2_2 _6170_ (.A0(_1450_),
    .A1(_1452_),
    .S(net11),
    .X(_1453_));
 sky130_fd_sc_hd__o21a_1 _6171_ (.A1(_0514_),
    .A2(_1212_),
    .B1(_0512_),
    .X(_1454_));
 sky130_fd_sc_hd__xor2_2 _6172_ (.A(_0464_),
    .B(_1454_),
    .X(_1455_));
 sky130_fd_sc_hd__xor2_1 _6173_ (.A(_0514_),
    .B(_1212_),
    .X(_1456_));
 sky130_fd_sc_hd__or2_1 _6174_ (.A(_1230_),
    .B(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__or3b_1 _6175_ (.A(_1457_),
    .B(_1224_),
    .C_N(_1227_),
    .X(_1458_));
 sky130_fd_sc_hd__o221a_1 _6176_ (.A1(net65),
    .A2(net101),
    .B1(_1404_),
    .B2(_1455_),
    .C1(_1458_),
    .X(_1459_));
 sky130_fd_sc_hd__nand2_1 _6177_ (.A(_1233_),
    .B(_1441_),
    .Y(_1460_));
 sky130_fd_sc_hd__o221a_1 _6178_ (.A1(net87),
    .A2(net101),
    .B1(_1457_),
    .B2(_1228_),
    .C1(_1460_),
    .X(_1461_));
 sky130_fd_sc_hd__mux2_1 _6179_ (.A0(_1461_),
    .A1(_1459_),
    .S(net9),
    .X(_1463_));
 sky130_fd_sc_hd__and3_1 _6180_ (.A(_1213_),
    .B(_1214_),
    .C(_1223_),
    .X(_1464_));
 sky130_fd_sc_hd__o21ai_1 _6181_ (.A1(_1224_),
    .A2(_1464_),
    .B1(_1405_),
    .Y(_1465_));
 sky130_fd_sc_hd__o221a_1 _6182_ (.A1(_3464_),
    .A2(net101),
    .B1(_1234_),
    .B2(_1455_),
    .C1(_1465_),
    .X(_1466_));
 sky130_fd_sc_hd__mux2_1 _6183_ (.A0(_1466_),
    .A1(_1277_),
    .S(net9),
    .X(_1467_));
 sky130_fd_sc_hd__mux2_1 _6184_ (.A0(_1463_),
    .A1(_1467_),
    .S(net12),
    .X(_1468_));
 sky130_fd_sc_hd__mux2_2 _6185_ (.A0(_1453_),
    .A1(_1468_),
    .S(_1412_),
    .X(_1469_));
 sky130_fd_sc_hd__mux2_8 _6186_ (.A0(_1448_),
    .A1(_1469_),
    .S(net14),
    .X(_1470_));
 sky130_fd_sc_hd__xor2_4 _6187_ (.A(net234),
    .B(net231),
    .X(_1471_));
 sky130_fd_sc_hd__xnor2_4 _6188_ (.A(net234),
    .B(net231),
    .Y(_1472_));
 sky130_fd_sc_hd__a31o_1 _6189_ (.A1(_1355_),
    .A2(_1379_),
    .A3(_1382_),
    .B1(_1438_),
    .X(_1474_));
 sky130_fd_sc_hd__o21a_1 _6190_ (.A1(_1390_),
    .A2(_1430_),
    .B1(_1474_),
    .X(_1475_));
 sky130_fd_sc_hd__a31o_1 _6191_ (.A1(_1355_),
    .A2(_1379_),
    .A3(_1382_),
    .B1(_1432_),
    .X(_1476_));
 sky130_fd_sc_hd__or4_1 _6192_ (.A(_1354_),
    .B(_1380_),
    .C(_1381_),
    .D(_1406_),
    .X(_1477_));
 sky130_fd_sc_hd__and3_1 _6193_ (.A(_1388_),
    .B(_1476_),
    .C(_1477_),
    .X(_1478_));
 sky130_fd_sc_hd__mux2_1 _6194_ (.A0(_1443_),
    .A1(_1461_),
    .S(net9),
    .X(_1479_));
 sky130_fd_sc_hd__mux2_1 _6195_ (.A0(_1459_),
    .A1(_1466_),
    .S(net9),
    .X(_1480_));
 sky130_fd_sc_hd__mux2_2 _6196_ (.A0(_1479_),
    .A1(_1480_),
    .S(net12),
    .X(_1481_));
 sky130_fd_sc_hd__a211o_1 _6197_ (.A1(net12),
    .A2(_1475_),
    .B1(_1478_),
    .C1(net7),
    .X(_1482_));
 sky130_fd_sc_hd__o21ai_2 _6198_ (.A1(_1412_),
    .A2(_1481_),
    .B1(_1482_),
    .Y(_1483_));
 sky130_fd_sc_hd__mux2_2 _6199_ (.A0(_1420_),
    .A1(_1399_),
    .S(net9),
    .X(_1485_));
 sky130_fd_sc_hd__and3_1 _6200_ (.A(net12),
    .B(_1476_),
    .C(_1477_),
    .X(_1486_));
 sky130_fd_sc_hd__a21oi_2 _6201_ (.A1(_1388_),
    .A2(_1485_),
    .B1(_1486_),
    .Y(_1487_));
 sky130_fd_sc_hd__o211a_1 _6202_ (.A1(net9),
    .A2(_1430_),
    .B1(_1474_),
    .C1(net13),
    .X(_1488_));
 sky130_fd_sc_hd__a21oi_1 _6203_ (.A1(net12),
    .A2(_1479_),
    .B1(_1488_),
    .Y(_1489_));
 sky130_fd_sc_hd__mux2_2 _6204_ (.A0(_1487_),
    .A1(_1489_),
    .S(net7),
    .X(_1490_));
 sky130_fd_sc_hd__xor2_4 _6205_ (.A(_1031_),
    .B(_1196_),
    .X(_1491_));
 sky130_fd_sc_hd__a2bb2o_1 _6206_ (.A1_N(_1404_),
    .A2_N(_1416_),
    .B1(_1491_),
    .B2(_1233_),
    .X(_1492_));
 sky130_fd_sc_hd__a31o_1 _6207_ (.A1(_1355_),
    .A2(_1379_),
    .A3(_1382_),
    .B1(_1417_),
    .X(_1493_));
 sky130_fd_sc_hd__o21a_1 _6208_ (.A1(net10),
    .A2(_1492_),
    .B1(_1493_),
    .X(_1494_));
 sky130_fd_sc_hd__o211a_1 _6209_ (.A1(net10),
    .A2(_1492_),
    .B1(_1493_),
    .C1(net13),
    .X(_1496_));
 sky130_fd_sc_hd__a21o_1 _6210_ (.A1(net11),
    .A2(_1485_),
    .B1(_1496_),
    .X(_1497_));
 sky130_fd_sc_hd__a211o_1 _6211_ (.A1(net12),
    .A2(_1475_),
    .B1(_1478_),
    .C1(_1412_),
    .X(_1498_));
 sky130_fd_sc_hd__a211o_1 _6212_ (.A1(net12),
    .A2(_1485_),
    .B1(_1496_),
    .C1(net8),
    .X(_1499_));
 sky130_fd_sc_hd__a31o_1 _6213_ (.A1(_1355_),
    .A2(_1379_),
    .A3(_1382_),
    .B1(_1278_),
    .X(_1500_));
 sky130_fd_sc_hd__o21a_1 _6214_ (.A1(_1277_),
    .A2(net10),
    .B1(_1500_),
    .X(_1501_));
 sky130_fd_sc_hd__o211a_1 _6215_ (.A1(_1277_),
    .A2(net9),
    .B1(_1500_),
    .C1(net12),
    .X(_1502_));
 sky130_fd_sc_hd__a21o_1 _6216_ (.A1(net13),
    .A2(_1480_),
    .B1(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__a21oi_1 _6217_ (.A1(net13),
    .A2(_1480_),
    .B1(_1502_),
    .Y(_1504_));
 sky130_fd_sc_hd__mux2_2 _6218_ (.A0(_1489_),
    .A1(_1504_),
    .S(net7),
    .X(_1505_));
 sky130_fd_sc_hd__and3_1 _6219_ (.A(net13),
    .B(_1444_),
    .C(_1445_),
    .X(_1507_));
 sky130_fd_sc_hd__a21oi_1 _6220_ (.A1(net12),
    .A2(_1463_),
    .B1(_1507_),
    .Y(_1508_));
 sky130_fd_sc_hd__o211a_1 _6221_ (.A1(_1278_),
    .A2(net10),
    .B1(_1449_),
    .C1(net11),
    .X(_1509_));
 sky130_fd_sc_hd__a21oi_2 _6222_ (.A1(net13),
    .A2(_1467_),
    .B1(_1509_),
    .Y(_1510_));
 sky130_fd_sc_hd__mux2_1 _6223_ (.A0(_1508_),
    .A1(_1510_),
    .S(net7),
    .X(_1511_));
 sky130_fd_sc_hd__mux2_1 _6224_ (.A0(_1409_),
    .A1(_1434_),
    .S(net12),
    .X(_1512_));
 sky130_fd_sc_hd__mux2_1 _6225_ (.A0(_1508_),
    .A1(_1512_),
    .S(_1412_),
    .X(_1513_));
 sky130_fd_sc_hd__mux2_2 _6226_ (.A0(_1447_),
    .A1(_1468_),
    .S(net7),
    .X(_1514_));
 sky130_fd_sc_hd__xnor2_4 _6227_ (.A(_1100_),
    .B(_1194_),
    .Y(_1515_));
 sky130_fd_sc_hd__and2_1 _6228_ (.A(_1095_),
    .B(_1195_),
    .X(_1516_));
 sky130_fd_sc_hd__a21oi_1 _6229_ (.A1(_1097_),
    .A2(_1516_),
    .B1(_1230_),
    .Y(_1518_));
 sky130_fd_sc_hd__o21a_2 _6230_ (.A1(_1097_),
    .A2(_1516_),
    .B1(_1518_),
    .X(_1519_));
 sky130_fd_sc_hd__inv_2 _6231_ (.A(_1519_),
    .Y(_1520_));
 sky130_fd_sc_hd__o22ai_2 _6232_ (.A1(_1234_),
    .A2(_1515_),
    .B1(_1520_),
    .B2(_1228_),
    .Y(_1521_));
 sky130_fd_sc_hd__a32o_1 _6233_ (.A1(_1135_),
    .A2(_1183_),
    .A3(_1184_),
    .B1(_0944_),
    .B2(_0587_),
    .X(_1522_));
 sky130_fd_sc_hd__o21ba_1 _6234_ (.A1(_1182_),
    .A2(_1522_),
    .B1_N(_1186_),
    .X(_1523_));
 sky130_fd_sc_hd__o22a_1 _6235_ (.A1(_0548_),
    .A2(_0587_),
    .B1(_0744_),
    .B2(_1134_),
    .X(_1524_));
 sky130_fd_sc_hd__and2_1 _6236_ (.A(_1173_),
    .B(_1178_),
    .X(_1525_));
 sky130_fd_sc_hd__mux2_1 _6237_ (.A0(_1525_),
    .A1(_1190_),
    .S(_1171_),
    .X(_1526_));
 sky130_fd_sc_hd__or3b_1 _6238_ (.A(_1523_),
    .B(_1524_),
    .C_N(_1526_),
    .X(_1527_));
 sky130_fd_sc_hd__xnor2_1 _6239_ (.A(_1129_),
    .B(_1192_),
    .Y(_1529_));
 sky130_fd_sc_hd__nand2_1 _6240_ (.A(_1515_),
    .B(_1529_),
    .Y(_1530_));
 sky130_fd_sc_hd__xnor2_1 _6241_ (.A(_1129_),
    .B(_1193_),
    .Y(_1531_));
 sky130_fd_sc_hd__mux2_1 _6242_ (.A0(_1530_),
    .A1(_1531_),
    .S(_1228_),
    .X(_1532_));
 sky130_fd_sc_hd__a211o_2 _6243_ (.A1(_1152_),
    .A2(_1192_),
    .B1(_1527_),
    .C1(_1532_),
    .X(_1533_));
 sky130_fd_sc_hd__a22o_1 _6244_ (.A1(net10),
    .A2(_1521_),
    .B1(_1533_),
    .B2(net101),
    .X(_1534_));
 sky130_fd_sc_hd__or3_1 _6245_ (.A(net11),
    .B(_1421_),
    .C(_1534_),
    .X(_1535_));
 sky130_fd_sc_hd__a22o_1 _6246_ (.A1(_1405_),
    .A2(_1491_),
    .B1(_1519_),
    .B2(_1228_),
    .X(_1536_));
 sky130_fd_sc_hd__mux2_1 _6247_ (.A0(_1521_),
    .A1(_1492_),
    .S(net10),
    .X(_1537_));
 sky130_fd_sc_hd__or2_2 _6248_ (.A(_1536_),
    .B(_1537_),
    .X(_1538_));
 sky130_fd_sc_hd__o41a_1 _6249_ (.A1(net13),
    .A2(_1410_),
    .A3(_1412_),
    .A4(_1538_),
    .B1(_1535_),
    .X(_1540_));
 sky130_fd_sc_hd__nand2_1 _6250_ (.A(_1487_),
    .B(_1512_),
    .Y(_1541_));
 sky130_fd_sc_hd__a211o_1 _6251_ (.A1(_1387_),
    .A2(_1538_),
    .B1(_1534_),
    .C1(net8),
    .X(_1542_));
 sky130_fd_sc_hd__o31a_1 _6252_ (.A1(_1497_),
    .A2(_1540_),
    .A3(_1541_),
    .B1(_1542_),
    .X(_1543_));
 sky130_fd_sc_hd__a211o_1 _6253_ (.A1(net8),
    .A2(_1534_),
    .B1(_1494_),
    .C1(_1421_),
    .X(_1544_));
 sky130_fd_sc_hd__mux2_1 _6254_ (.A0(_1538_),
    .A1(_1544_),
    .S(net11),
    .X(_1545_));
 sky130_fd_sc_hd__nand4_1 _6255_ (.A(_1483_),
    .B(_1490_),
    .C(_1505_),
    .D(_1511_),
    .Y(_1546_));
 sky130_fd_sc_hd__a21bo_1 _6256_ (.A1(_1498_),
    .A2(_1499_),
    .B1_N(_1513_),
    .X(_1547_));
 sky130_fd_sc_hd__o41a_1 _6257_ (.A1(_1448_),
    .A2(_1514_),
    .A3(_1546_),
    .A4(_1547_),
    .B1(net14),
    .X(_1548_));
 sky130_fd_sc_hd__or4_1 _6258_ (.A(_1470_),
    .B(_1543_),
    .C(_1545_),
    .D(_1548_),
    .X(_1549_));
 sky130_fd_sc_hd__and3_1 _6259_ (.A(_1354_),
    .B(_1359_),
    .C(_1375_),
    .X(_1551_));
 sky130_fd_sc_hd__a21oi_2 _6260_ (.A1(net15),
    .A2(net6),
    .B1(_1551_),
    .Y(_1552_));
 sky130_fd_sc_hd__a21o_1 _6261_ (.A1(_1549_),
    .A2(_1552_),
    .B1(net225),
    .X(_1553_));
 sky130_fd_sc_hd__mux2_1 _6262_ (.A0(_1276_),
    .A1(_1350_),
    .S(net10),
    .X(_1554_));
 sky130_fd_sc_hd__mux2_1 _6263_ (.A0(_1501_),
    .A1(_1554_),
    .S(net11),
    .X(_1555_));
 sky130_fd_sc_hd__mux2_2 _6264_ (.A0(_1481_),
    .A1(_1555_),
    .S(net6),
    .X(_1556_));
 sky130_fd_sc_hd__a21o_1 _6265_ (.A1(_1498_),
    .A2(_1499_),
    .B1(net14),
    .X(_1557_));
 sky130_fd_sc_hd__o21a_1 _6266_ (.A1(_1384_),
    .A2(_1556_),
    .B1(_1557_),
    .X(_1558_));
 sky130_fd_sc_hd__and3_1 _6267_ (.A(_1470_),
    .B(_1553_),
    .C(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__and3b_4 _6268_ (.A_N(\cmd[6] ),
    .B(_1215_),
    .C(\cmd[7] ),
    .X(_1560_));
 sky130_fd_sc_hd__or3b_4 _6269_ (.A(\cmd[6] ),
    .B(_1216_),
    .C_N(\cmd[7] ),
    .X(_1562_));
 sky130_fd_sc_hd__a21oi_1 _6270_ (.A1(_1553_),
    .A2(_1558_),
    .B1(_1470_),
    .Y(_1563_));
 sky130_fd_sc_hd__nand2_1 _6271_ (.A(net203),
    .B(_2221_),
    .Y(_1564_));
 sky130_fd_sc_hd__nor2_1 _6272_ (.A(net203),
    .B(_2221_),
    .Y(_1565_));
 sky130_fd_sc_hd__or2_1 _6273_ (.A(_1330_),
    .B(_2342_),
    .X(_1566_));
 sky130_fd_sc_hd__nor2_1 _6274_ (.A(_1561_),
    .B(_2617_),
    .Y(_1567_));
 sky130_fd_sc_hd__a211o_1 _6275_ (.A1(\posit_add.in1[1] ),
    .A2(_2914_),
    .B1(_0657_),
    .C1(net235),
    .X(_1568_));
 sky130_fd_sc_hd__o221a_1 _6276_ (.A1(_1484_),
    .A2(_2804_),
    .B1(_2914_),
    .B2(_1517_),
    .C1(_1568_),
    .X(_1569_));
 sky130_fd_sc_hd__a22o_1 _6277_ (.A1(_1671_),
    .A2(_2749_),
    .B1(_2804_),
    .B2(_1484_),
    .X(_1570_));
 sky130_fd_sc_hd__or2_1 _6278_ (.A(_1671_),
    .B(_2749_),
    .X(_1571_));
 sky130_fd_sc_hd__o221a_1 _6279_ (.A1(_1638_),
    .A2(_2705_),
    .B1(_1569_),
    .B2(_1570_),
    .C1(_1571_),
    .X(_1573_));
 sky130_fd_sc_hd__a22o_1 _6280_ (.A1(_1594_),
    .A2(_2661_),
    .B1(_2705_),
    .B2(_1638_),
    .X(_1574_));
 sky130_fd_sc_hd__o22a_1 _6281_ (.A1(_1594_),
    .A2(_2661_),
    .B1(_1573_),
    .B2(_1574_),
    .X(_1575_));
 sky130_fd_sc_hd__a21oi_1 _6282_ (.A1(_1561_),
    .A2(_2617_),
    .B1(_1575_),
    .Y(_1576_));
 sky130_fd_sc_hd__o22a_1 _6283_ (.A1(_1154_),
    .A2(_2529_),
    .B1(_1567_),
    .B2(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__a221o_1 _6284_ (.A1(_1154_),
    .A2(_2529_),
    .B1(_2551_),
    .B2(_1110_),
    .C1(_1577_),
    .X(_1578_));
 sky130_fd_sc_hd__o2bb2a_1 _6285_ (.A1_N(_1242_),
    .A2_N(_2430_),
    .B1(_2551_),
    .B2(_1110_),
    .X(_1579_));
 sky130_fd_sc_hd__o22ai_1 _6286_ (.A1(_1209_),
    .A2(_2397_),
    .B1(_2430_),
    .B2(_1242_),
    .Y(_1580_));
 sky130_fd_sc_hd__a21oi_1 _6287_ (.A1(_1578_),
    .A2(_1579_),
    .B1(_1580_),
    .Y(_1581_));
 sky130_fd_sc_hd__a22o_1 _6288_ (.A1(_1407_),
    .A2(_2287_),
    .B1(_2397_),
    .B2(_1209_),
    .X(_1582_));
 sky130_fd_sc_hd__or2_1 _6289_ (.A(_1363_),
    .B(_2243_),
    .X(_1584_));
 sky130_fd_sc_hd__o221a_1 _6290_ (.A1(_1407_),
    .A2(_2287_),
    .B1(_1581_),
    .B2(_1582_),
    .C1(_1584_),
    .X(_1585_));
 sky130_fd_sc_hd__a221o_1 _6291_ (.A1(_1363_),
    .A2(_2243_),
    .B1(_2342_),
    .B2(_1330_),
    .C1(_1585_),
    .X(_1586_));
 sky130_fd_sc_hd__a31o_4 _6292_ (.A1(_1564_),
    .A2(_1566_),
    .A3(_1586_),
    .B1(_1565_),
    .X(_1587_));
 sky130_fd_sc_hd__mux2_4 _6293_ (.A0(_1303_),
    .A1(_1299_),
    .S(net97),
    .X(_1588_));
 sky130_fd_sc_hd__mux2_8 _6294_ (.A0(_1254_),
    .A1(_1259_),
    .S(net98),
    .X(_1589_));
 sky130_fd_sc_hd__a21o_1 _6295_ (.A1(_2221_),
    .A2(net189),
    .B1(net192),
    .X(_1590_));
 sky130_fd_sc_hd__and2_2 _6296_ (.A(_1302_),
    .B(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__mux2_8 _6297_ (.A0(_1591_),
    .A1(_1287_),
    .S(net98),
    .X(_1592_));
 sky130_fd_sc_hd__a21o_2 _6298_ (.A1(_1589_),
    .A2(_1592_),
    .B1(_1333_),
    .X(_1593_));
 sky130_fd_sc_hd__xnor2_4 _6299_ (.A(_1588_),
    .B(_1593_),
    .Y(_1595_));
 sky130_fd_sc_hd__a31o_4 _6300_ (.A1(_1588_),
    .A2(_1589_),
    .A3(_1592_),
    .B1(_1333_),
    .X(_1596_));
 sky130_fd_sc_hd__mux2_8 _6301_ (.A0(_1317_),
    .A1(_1321_),
    .S(net98),
    .X(_1597_));
 sky130_fd_sc_hd__xor2_4 _6302_ (.A(_1596_),
    .B(_1597_),
    .X(_1598_));
 sky130_fd_sc_hd__xnor2_1 _6303_ (.A(_1595_),
    .B(_1598_),
    .Y(_1599_));
 sky130_fd_sc_hd__or2_4 _6304_ (.A(_1333_),
    .B(_1589_),
    .X(_1600_));
 sky130_fd_sc_hd__xnor2_4 _6305_ (.A(_1592_),
    .B(_1600_),
    .Y(_1601_));
 sky130_fd_sc_hd__inv_2 _6306_ (.A(_1601_),
    .Y(_1602_));
 sky130_fd_sc_hd__nand2_1 _6307_ (.A(_1595_),
    .B(_1602_),
    .Y(_1603_));
 sky130_fd_sc_hd__xnor2_2 _6308_ (.A(_1595_),
    .B(_1601_),
    .Y(_1604_));
 sky130_fd_sc_hd__nor2_1 _6309_ (.A(_3434_),
    .B(_1250_),
    .Y(_1606_));
 sky130_fd_sc_hd__xnor2_4 _6310_ (.A(_3435_),
    .B(_1250_),
    .Y(_1607_));
 sky130_fd_sc_hd__nor2_1 _6311_ (.A(_3445_),
    .B(net97),
    .Y(_1608_));
 sky130_fd_sc_hd__a21o_2 _6312_ (.A1(_1241_),
    .A2(net97),
    .B1(_1608_),
    .X(_1609_));
 sky130_fd_sc_hd__o211a_1 _6313_ (.A1(_1236_),
    .A2(_1239_),
    .B1(_1240_),
    .C1(_3445_),
    .X(_1610_));
 sky130_fd_sc_hd__a211o_4 _6314_ (.A1(_1241_),
    .A2(net97),
    .B1(_1608_),
    .C1(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__xnor2_1 _6315_ (.A(_3434_),
    .B(net97),
    .Y(_1612_));
 sky130_fd_sc_hd__mux2_8 _6316_ (.A0(_1611_),
    .A1(_1612_),
    .S(_1607_),
    .X(_1613_));
 sky130_fd_sc_hd__nor2_1 _6317_ (.A(_3384_),
    .B(net97),
    .Y(_1614_));
 sky130_fd_sc_hd__a21oi_4 _6318_ (.A1(_2100_),
    .A2(net97),
    .B1(_1614_),
    .Y(_1615_));
 sky130_fd_sc_hd__o2bb2ai_4 _6319_ (.A1_N(_1273_),
    .A2_N(_1613_),
    .B1(_1615_),
    .B2(_1272_),
    .Y(_1617_));
 sky130_fd_sc_hd__xnor2_4 _6320_ (.A(_1265_),
    .B(_1617_),
    .Y(_1618_));
 sky130_fd_sc_hd__inv_2 _6321_ (.A(_1618_),
    .Y(_1619_));
 sky130_fd_sc_hd__xnor2_4 _6322_ (.A(_1273_),
    .B(_1613_),
    .Y(_1620_));
 sky130_fd_sc_hd__mux2_2 _6323_ (.A0(_1260_),
    .A1(_1255_),
    .S(net97),
    .X(_1621_));
 sky130_fd_sc_hd__a2bb2o_2 _6324_ (.A1_N(_1589_),
    .A2_N(_1621_),
    .B1(_1617_),
    .B2(_1266_),
    .X(_1622_));
 sky130_fd_sc_hd__nand2_1 _6325_ (.A(_1293_),
    .B(_1622_),
    .Y(_1623_));
 sky130_fd_sc_hd__nor2_1 _6326_ (.A(net204),
    .B(net216),
    .Y(_1624_));
 sky130_fd_sc_hd__nand2b_1 _6327_ (.A_N(_1624_),
    .B(_1621_),
    .Y(_1625_));
 sky130_fd_sc_hd__mux2_2 _6328_ (.A0(_1287_),
    .A1(_1591_),
    .S(net98),
    .X(_1626_));
 sky130_fd_sc_hd__inv_2 _6329_ (.A(_1626_),
    .Y(_1628_));
 sky130_fd_sc_hd__xnor2_1 _6330_ (.A(_1625_),
    .B(_1626_),
    .Y(_1629_));
 sky130_fd_sc_hd__a22o_1 _6331_ (.A1(_1293_),
    .A2(_1622_),
    .B1(_1629_),
    .B2(_1602_),
    .X(_1630_));
 sky130_fd_sc_hd__o21ba_1 _6332_ (.A1(_1621_),
    .A2(_1628_),
    .B1_N(_1624_),
    .X(_1631_));
 sky130_fd_sc_hd__mux2_1 _6333_ (.A0(_1299_),
    .A1(_1303_),
    .S(net98),
    .X(_1632_));
 sky130_fd_sc_hd__xnor2_1 _6334_ (.A(_1631_),
    .B(_1632_),
    .Y(_1633_));
 sky130_fd_sc_hd__a2bb2o_2 _6335_ (.A1_N(_1595_),
    .A2_N(_1633_),
    .B1(_1630_),
    .B2(_1310_),
    .X(_1634_));
 sky130_fd_sc_hd__nor2_1 _6336_ (.A(_1624_),
    .B(_1632_),
    .Y(_1635_));
 sky130_fd_sc_hd__mux2_1 _6337_ (.A0(_1321_),
    .A1(_1317_),
    .S(net98),
    .X(_1636_));
 sky130_fd_sc_hd__or3_1 _6338_ (.A(_1631_),
    .B(_1635_),
    .C(_1636_),
    .X(_1637_));
 sky130_fd_sc_hd__o21ai_1 _6339_ (.A1(_1631_),
    .A2(_1635_),
    .B1(_1636_),
    .Y(_1639_));
 sky130_fd_sc_hd__a32o_2 _6340_ (.A1(_1598_),
    .A2(_1637_),
    .A3(_1639_),
    .B1(_1634_),
    .B2(_1326_),
    .X(_1640_));
 sky130_fd_sc_hd__xnor2_2 _6341_ (.A(_1327_),
    .B(_1634_),
    .Y(_1641_));
 sky130_fd_sc_hd__or2_1 _6342_ (.A(_1293_),
    .B(_1622_),
    .X(_1642_));
 sky130_fd_sc_hd__xnor2_1 _6343_ (.A(_1309_),
    .B(_1630_),
    .Y(_1643_));
 sky130_fd_sc_hd__a21o_1 _6344_ (.A1(_1623_),
    .A2(_1642_),
    .B1(_1643_),
    .X(_1644_));
 sky130_fd_sc_hd__a211oi_4 _6345_ (.A1(_1336_),
    .A2(_1640_),
    .B1(_1641_),
    .C1(_1644_),
    .Y(_1645_));
 sky130_fd_sc_hd__and2_4 _6346_ (.A(_1620_),
    .B(_1645_),
    .X(_1646_));
 sky130_fd_sc_hd__nand2_1 _6347_ (.A(_1620_),
    .B(_1645_),
    .Y(_1647_));
 sky130_fd_sc_hd__xor2_4 _6348_ (.A(_1607_),
    .B(_1611_),
    .X(_1648_));
 sky130_fd_sc_hd__and2_1 _6349_ (.A(_3446_),
    .B(_1241_),
    .X(_1650_));
 sky130_fd_sc_hd__or2_4 _6350_ (.A(_1610_),
    .B(_1650_),
    .X(_1651_));
 sky130_fd_sc_hd__inv_2 _6351_ (.A(_1651_),
    .Y(_1652_));
 sky130_fd_sc_hd__and2_2 _6352_ (.A(_1645_),
    .B(_1651_),
    .X(_1653_));
 sky130_fd_sc_hd__nand2_1 _6353_ (.A(_1215_),
    .B(net62),
    .Y(_1654_));
 sky130_fd_sc_hd__and3_1 _6354_ (.A(_1215_),
    .B(_1648_),
    .C(net62),
    .X(_1655_));
 sky130_fd_sc_hd__or3b_4 _6355_ (.A(_1618_),
    .B(net63),
    .C_N(_1655_),
    .X(_1656_));
 sky130_fd_sc_hd__and2_2 _6356_ (.A(_1619_),
    .B(_1645_),
    .X(_1657_));
 sky130_fd_sc_hd__nand2_2 _6357_ (.A(_1619_),
    .B(_1645_),
    .Y(_1658_));
 sky130_fd_sc_hd__and2_4 _6358_ (.A(_1645_),
    .B(_1648_),
    .X(_1659_));
 sky130_fd_sc_hd__nand2_4 _6359_ (.A(_1645_),
    .B(_1648_),
    .Y(_1661_));
 sky130_fd_sc_hd__mux2_1 _6360_ (.A0(_3464_),
    .A1(net128),
    .S(net100),
    .X(_1662_));
 sky130_fd_sc_hd__mux2_2 _6361_ (.A0(_1215_),
    .A1(_1662_),
    .S(net62),
    .X(_1663_));
 sky130_fd_sc_hd__nand2_1 _6362_ (.A(_1659_),
    .B(_1663_),
    .Y(_1664_));
 sky130_fd_sc_hd__and3_1 _6363_ (.A(_1620_),
    .B(_1659_),
    .C(_1663_),
    .X(_1665_));
 sky130_fd_sc_hd__nand2_1 _6364_ (.A(_1657_),
    .B(_1665_),
    .Y(_1666_));
 sky130_fd_sc_hd__mux2_4 _6365_ (.A0(_3476_),
    .A1(net69),
    .S(net99),
    .X(_1667_));
 sky130_fd_sc_hd__nor2_2 _6366_ (.A(_1666_),
    .B(_1667_),
    .Y(_1668_));
 sky130_fd_sc_hd__mux2_1 _6367_ (.A0(net64),
    .A1(net162),
    .S(net100),
    .X(_1669_));
 sky130_fd_sc_hd__or3b_1 _6368_ (.A(_1652_),
    .B(_1669_),
    .C_N(_1645_),
    .X(_1670_));
 sky130_fd_sc_hd__o21ai_1 _6369_ (.A1(net62),
    .A2(_1662_),
    .B1(_1670_),
    .Y(_1672_));
 sky130_fd_sc_hd__o22a_1 _6370_ (.A1(_1648_),
    .A2(_1654_),
    .B1(_1661_),
    .B2(_1672_),
    .X(_1673_));
 sky130_fd_sc_hd__or2_4 _6371_ (.A(net63),
    .B(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__mux2_2 _6372_ (.A0(net162),
    .A1(net64),
    .S(net99),
    .X(_1675_));
 sky130_fd_sc_hd__or3b_2 _6373_ (.A(_1618_),
    .B(_1674_),
    .C_N(_1675_),
    .X(_1676_));
 sky130_fd_sc_hd__or3_2 _6374_ (.A(_1618_),
    .B(_1674_),
    .C(_1675_),
    .X(_1677_));
 sky130_fd_sc_hd__o21a_1 _6375_ (.A1(_1618_),
    .A2(_1674_),
    .B1(_1675_),
    .X(_1678_));
 sky130_fd_sc_hd__inv_2 _6376_ (.A(_1678_),
    .Y(_1679_));
 sky130_fd_sc_hd__nand2_4 _6377_ (.A(_1677_),
    .B(_1679_),
    .Y(_1680_));
 sky130_fd_sc_hd__inv_2 _6378_ (.A(_1680_),
    .Y(_1681_));
 sky130_fd_sc_hd__mux2_1 _6379_ (.A0(net88),
    .A1(net157),
    .S(net100),
    .X(_1683_));
 sky130_fd_sc_hd__mux2_1 _6380_ (.A0(_1669_),
    .A1(_1683_),
    .S(net62),
    .X(_1684_));
 sky130_fd_sc_hd__or2_1 _6381_ (.A(_1661_),
    .B(_1684_),
    .X(_1685_));
 sky130_fd_sc_hd__o21ai_2 _6382_ (.A1(_1659_),
    .A2(_1663_),
    .B1(_1685_),
    .Y(_1686_));
 sky130_fd_sc_hd__nor2_2 _6383_ (.A(net63),
    .B(_1686_),
    .Y(_1687_));
 sky130_fd_sc_hd__nand2_4 _6384_ (.A(_1619_),
    .B(_1687_),
    .Y(_1688_));
 sky130_fd_sc_hd__mux2_8 _6385_ (.A0(net157),
    .A1(net87),
    .S(net100),
    .X(_1689_));
 sky130_fd_sc_hd__and3_1 _6386_ (.A(_1619_),
    .B(_1687_),
    .C(_1689_),
    .X(_1690_));
 sky130_fd_sc_hd__xnor2_4 _6387_ (.A(_1688_),
    .B(_1689_),
    .Y(_1691_));
 sky130_fd_sc_hd__mux2_1 _6388_ (.A0(_0364_),
    .A1(net154),
    .S(net99),
    .X(_1692_));
 sky130_fd_sc_hd__mux2_1 _6389_ (.A0(_1683_),
    .A1(_1692_),
    .S(net62),
    .X(_1694_));
 sky130_fd_sc_hd__nor2_1 _6390_ (.A(_1661_),
    .B(_1694_),
    .Y(_1695_));
 sky130_fd_sc_hd__a21oi_1 _6391_ (.A1(_1661_),
    .A2(_1672_),
    .B1(_1695_),
    .Y(_1696_));
 sky130_fd_sc_hd__mux2_4 _6392_ (.A0(_1655_),
    .A1(_1696_),
    .S(_1646_),
    .X(_1697_));
 sky130_fd_sc_hd__and2_1 _6393_ (.A(net61),
    .B(_1697_),
    .X(_1698_));
 sky130_fd_sc_hd__nand2_1 _6394_ (.A(net61),
    .B(_1697_),
    .Y(_1699_));
 sky130_fd_sc_hd__mux2_2 _6395_ (.A0(net154),
    .A1(_0364_),
    .S(net99),
    .X(_1700_));
 sky130_fd_sc_hd__or2_2 _6396_ (.A(_1699_),
    .B(_1700_),
    .X(_1701_));
 sky130_fd_sc_hd__and2_1 _6397_ (.A(_1699_),
    .B(_1700_),
    .X(_1702_));
 sky130_fd_sc_hd__inv_2 _6398_ (.A(_1702_),
    .Y(_1703_));
 sky130_fd_sc_hd__nand2_4 _6399_ (.A(_1701_),
    .B(_1703_),
    .Y(_1705_));
 sky130_fd_sc_hd__mux2_1 _6400_ (.A0(net83),
    .A1(net146),
    .S(net100),
    .X(_1706_));
 sky130_fd_sc_hd__mux2_1 _6401_ (.A0(_1692_),
    .A1(_1706_),
    .S(net62),
    .X(_1707_));
 sky130_fd_sc_hd__mux2_1 _6402_ (.A0(_1684_),
    .A1(_1707_),
    .S(_1659_),
    .X(_1708_));
 sky130_fd_sc_hd__a2bb2o_2 _6403_ (.A1_N(_1620_),
    .A2_N(_1664_),
    .B1(_1708_),
    .B2(_1646_),
    .X(_1709_));
 sky130_fd_sc_hd__nand2_1 _6404_ (.A(net61),
    .B(_1709_),
    .Y(_1710_));
 sky130_fd_sc_hd__mux2_2 _6405_ (.A0(net144),
    .A1(net82),
    .S(net100),
    .X(_1711_));
 sky130_fd_sc_hd__and2_1 _6406_ (.A(_1710_),
    .B(_1711_),
    .X(_1712_));
 sky130_fd_sc_hd__or2_2 _6407_ (.A(_1710_),
    .B(_1711_),
    .X(_1713_));
 sky130_fd_sc_hd__mux2_1 _6408_ (.A0(_0430_),
    .A1(_3498_),
    .S(net99),
    .X(_1714_));
 sky130_fd_sc_hd__mux2_1 _6409_ (.A0(_1706_),
    .A1(_1714_),
    .S(net62),
    .X(_1716_));
 sky130_fd_sc_hd__or2_1 _6410_ (.A(_1661_),
    .B(_1716_),
    .X(_1717_));
 sky130_fd_sc_hd__o21ai_1 _6411_ (.A1(_1659_),
    .A2(_1694_),
    .B1(_1717_),
    .Y(_1718_));
 sky130_fd_sc_hd__mux2_1 _6412_ (.A0(_1673_),
    .A1(_1718_),
    .S(_1646_),
    .X(_1719_));
 sky130_fd_sc_hd__or2_2 _6413_ (.A(_1658_),
    .B(_1719_),
    .X(_1720_));
 sky130_fd_sc_hd__mux2_1 _6414_ (.A0(_3498_),
    .A1(net80),
    .S(net100),
    .X(_1721_));
 sky130_fd_sc_hd__and2b_1 _6415_ (.A_N(_1720_),
    .B(_1721_),
    .X(_1722_));
 sky130_fd_sc_hd__or2_2 _6416_ (.A(_1720_),
    .B(_1721_),
    .X(_1723_));
 sky130_fd_sc_hd__and2_1 _6417_ (.A(_1720_),
    .B(_1721_),
    .X(_1724_));
 sky130_fd_sc_hd__nand2_1 _6418_ (.A(_1720_),
    .B(_1721_),
    .Y(_1725_));
 sky130_fd_sc_hd__nand2_4 _6419_ (.A(_1723_),
    .B(_1725_),
    .Y(_1727_));
 sky130_fd_sc_hd__mux2_1 _6420_ (.A0(net77),
    .A1(_3496_),
    .S(net99),
    .X(_1728_));
 sky130_fd_sc_hd__mux2_1 _6421_ (.A0(_1714_),
    .A1(_1728_),
    .S(_1653_),
    .X(_1729_));
 sky130_fd_sc_hd__or2_1 _6422_ (.A(_1661_),
    .B(_1729_),
    .X(_1730_));
 sky130_fd_sc_hd__o21ai_1 _6423_ (.A1(_1659_),
    .A2(_1707_),
    .B1(_1730_),
    .Y(_1731_));
 sky130_fd_sc_hd__mux2_1 _6424_ (.A0(_1686_),
    .A1(_1731_),
    .S(_1646_),
    .X(_1732_));
 sky130_fd_sc_hd__nor2_1 _6425_ (.A(_1658_),
    .B(_1732_),
    .Y(_1733_));
 sky130_fd_sc_hd__mux2_4 _6426_ (.A0(net179),
    .A1(net75),
    .S(net100),
    .X(_1734_));
 sky130_fd_sc_hd__inv_2 _6427_ (.A(_1734_),
    .Y(_1735_));
 sky130_fd_sc_hd__nand2_2 _6428_ (.A(_1733_),
    .B(_1735_),
    .Y(_1736_));
 sky130_fd_sc_hd__or2_2 _6429_ (.A(_1733_),
    .B(_1735_),
    .X(_1738_));
 sky130_fd_sc_hd__mux2_1 _6430_ (.A0(net113),
    .A1(net137),
    .S(net99),
    .X(_1739_));
 sky130_fd_sc_hd__mux2_1 _6431_ (.A0(_1728_),
    .A1(_1739_),
    .S(net62),
    .X(_1740_));
 sky130_fd_sc_hd__mux2_1 _6432_ (.A0(_1716_),
    .A1(_1740_),
    .S(_1659_),
    .X(_1741_));
 sky130_fd_sc_hd__o221a_1 _6433_ (.A1(_1620_),
    .A2(_1696_),
    .B1(_1741_),
    .B2(net63),
    .C1(net61),
    .X(_1742_));
 sky130_fd_sc_hd__a31o_1 _6434_ (.A1(_1618_),
    .A2(_1646_),
    .A3(_1655_),
    .B1(_1742_),
    .X(_1743_));
 sky130_fd_sc_hd__mux2_2 _6435_ (.A0(net137),
    .A1(net113),
    .S(net100),
    .X(_1744_));
 sky130_fd_sc_hd__and2_1 _6436_ (.A(_1743_),
    .B(_1744_),
    .X(_1745_));
 sky130_fd_sc_hd__nor2_1 _6437_ (.A(_1743_),
    .B(_1744_),
    .Y(_1746_));
 sky130_fd_sc_hd__mux2_2 _6438_ (.A0(_0548_),
    .A1(net124),
    .S(net99),
    .X(_1747_));
 sky130_fd_sc_hd__mux2_1 _6439_ (.A0(_1739_),
    .A1(_1747_),
    .S(net62),
    .X(_1749_));
 sky130_fd_sc_hd__mux2_1 _6440_ (.A0(_1729_),
    .A1(_1749_),
    .S(_1659_),
    .X(_1750_));
 sky130_fd_sc_hd__mux2_1 _6441_ (.A0(_1708_),
    .A1(_1750_),
    .S(_1646_),
    .X(_1751_));
 sky130_fd_sc_hd__or2_1 _6442_ (.A(_1658_),
    .B(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__or2_1 _6443_ (.A(net61),
    .B(_1665_),
    .X(_1753_));
 sky130_fd_sc_hd__nand2_1 _6444_ (.A(_1752_),
    .B(_1753_),
    .Y(_1754_));
 sky130_fd_sc_hd__mux2_4 _6445_ (.A0(net123),
    .A1(net106),
    .S(net100),
    .X(_1755_));
 sky130_fd_sc_hd__nor2_1 _6446_ (.A(_1754_),
    .B(_1755_),
    .Y(_1756_));
 sky130_fd_sc_hd__nand2_1 _6447_ (.A(_1754_),
    .B(_1755_),
    .Y(_1757_));
 sky130_fd_sc_hd__mux2_1 _6448_ (.A0(net105),
    .A1(net176),
    .S(net99),
    .X(_1758_));
 sky130_fd_sc_hd__nand2_1 _6449_ (.A(_1653_),
    .B(_1758_),
    .Y(_1760_));
 sky130_fd_sc_hd__o21ai_2 _6450_ (.A1(_1653_),
    .A2(_1747_),
    .B1(_1760_),
    .Y(_1761_));
 sky130_fd_sc_hd__nand2_1 _6451_ (.A(_1661_),
    .B(_1740_),
    .Y(_1762_));
 sky130_fd_sc_hd__o21ai_2 _6452_ (.A1(_1661_),
    .A2(_1761_),
    .B1(_1762_),
    .Y(_1763_));
 sky130_fd_sc_hd__nand2_1 _6453_ (.A(net63),
    .B(_1718_),
    .Y(_1764_));
 sky130_fd_sc_hd__o211a_1 _6454_ (.A1(net63),
    .A2(_1763_),
    .B1(_1764_),
    .C1(_1657_),
    .X(_1765_));
 sky130_fd_sc_hd__o21bai_4 _6455_ (.A1(_1619_),
    .A2(_1674_),
    .B1_N(_1765_),
    .Y(_1766_));
 sky130_fd_sc_hd__mux2_2 _6456_ (.A0(net176),
    .A1(net105),
    .S(net99),
    .X(_1767_));
 sky130_fd_sc_hd__and2b_1 _6457_ (.A_N(_1767_),
    .B(_1766_),
    .X(_1768_));
 sky130_fd_sc_hd__o21a_1 _6458_ (.A1(_1756_),
    .A2(_1768_),
    .B1(_1757_),
    .X(_1769_));
 sky130_fd_sc_hd__o21bai_2 _6459_ (.A1(_1745_),
    .A2(_1769_),
    .B1_N(_1746_),
    .Y(_1771_));
 sky130_fd_sc_hd__inv_2 _6460_ (.A(_1771_),
    .Y(_1772_));
 sky130_fd_sc_hd__a21boi_1 _6461_ (.A1(_1736_),
    .A2(_1771_),
    .B1_N(_1738_),
    .Y(_1773_));
 sky130_fd_sc_hd__a21oi_1 _6462_ (.A1(_1727_),
    .A2(_1773_),
    .B1(_1722_),
    .Y(_1774_));
 sky130_fd_sc_hd__o21a_1 _6463_ (.A1(_1712_),
    .A2(_1774_),
    .B1(_1713_),
    .X(_1775_));
 sky130_fd_sc_hd__nand2b_1 _6464_ (.A_N(_1775_),
    .B(_1705_),
    .Y(_1776_));
 sky130_fd_sc_hd__a21bo_2 _6465_ (.A1(_1698_),
    .A2(_1700_),
    .B1_N(_1776_),
    .X(_1777_));
 sky130_fd_sc_hd__a21oi_4 _6466_ (.A1(_1691_),
    .A2(_1777_),
    .B1(_1690_),
    .Y(_1778_));
 sky130_fd_sc_hd__o21ai_4 _6467_ (.A1(_1681_),
    .A2(_1778_),
    .B1(_1676_),
    .Y(_1779_));
 sky130_fd_sc_hd__nand2_2 _6468_ (.A(_1666_),
    .B(_1667_),
    .Y(_1780_));
 sky130_fd_sc_hd__a21oi_4 _6469_ (.A1(_1779_),
    .A2(_1780_),
    .B1(_1668_),
    .Y(_1782_));
 sky130_fd_sc_hd__a21bo_2 _6470_ (.A1(net213),
    .A2(net201),
    .B1_N(_1656_),
    .X(_1783_));
 sky130_fd_sc_hd__a21oi_4 _6471_ (.A1(_1656_),
    .A2(_1782_),
    .B1(net224),
    .Y(_1784_));
 sky130_fd_sc_hd__and2b_4 _6472_ (.A_N(_1668_),
    .B(_1780_),
    .X(_1785_));
 sky130_fd_sc_hd__a21oi_1 _6473_ (.A1(net61),
    .A2(_1709_),
    .B1(_1711_),
    .Y(_1786_));
 sky130_fd_sc_hd__nand2b_4 _6474_ (.A_N(_1712_),
    .B(_1713_),
    .Y(_1787_));
 sky130_fd_sc_hd__or2_2 _6475_ (.A(_1733_),
    .B(_1734_),
    .X(_1788_));
 sky130_fd_sc_hd__nand2_4 _6476_ (.A(_1736_),
    .B(_1738_),
    .Y(_1789_));
 sky130_fd_sc_hd__inv_2 _6477_ (.A(_1789_),
    .Y(_1790_));
 sky130_fd_sc_hd__and2b_1 _6478_ (.A_N(_1743_),
    .B(_1744_),
    .X(_1791_));
 sky130_fd_sc_hd__or2_4 _6479_ (.A(_1745_),
    .B(_1746_),
    .X(_1793_));
 sky130_fd_sc_hd__and2b_4 _6480_ (.A_N(_1756_),
    .B(_1757_),
    .X(_1794_));
 sky130_fd_sc_hd__nor2_2 _6481_ (.A(_1766_),
    .B(_1767_),
    .Y(_1795_));
 sky130_fd_sc_hd__and2_1 _6482_ (.A(_1766_),
    .B(_1767_),
    .X(_1796_));
 sky130_fd_sc_hd__nor2_1 _6483_ (.A(_1653_),
    .B(_1758_),
    .Y(_1797_));
 sky130_fd_sc_hd__mux2_1 _6484_ (.A0(_1749_),
    .A1(_1797_),
    .S(_1659_),
    .X(_1798_));
 sky130_fd_sc_hd__nor2_1 _6485_ (.A(net63),
    .B(_1798_),
    .Y(_1799_));
 sky130_fd_sc_hd__a21oi_1 _6486_ (.A1(net63),
    .A2(_1731_),
    .B1(_1799_),
    .Y(_1800_));
 sky130_fd_sc_hd__a22o_4 _6487_ (.A1(_1618_),
    .A2(_1687_),
    .B1(_1800_),
    .B2(net61),
    .X(_1801_));
 sky130_fd_sc_hd__nor2_1 _6488_ (.A(_1620_),
    .B(_1658_),
    .Y(_1802_));
 sky130_fd_sc_hd__o2bb2a_2 _6489_ (.A1_N(_1763_),
    .A2_N(_1802_),
    .B1(_1657_),
    .B2(_1719_),
    .X(_1804_));
 sky130_fd_sc_hd__o2bb2a_2 _6490_ (.A1_N(_1798_),
    .A2_N(_1802_),
    .B1(net61),
    .B2(_1732_),
    .X(_1805_));
 sky130_fd_sc_hd__nand2_2 _6491_ (.A(_1804_),
    .B(_1805_),
    .Y(_1806_));
 sky130_fd_sc_hd__nor2_1 _6492_ (.A(net63),
    .B(_1648_),
    .Y(_1807_));
 sky130_fd_sc_hd__a221o_2 _6493_ (.A1(net63),
    .A2(_1750_),
    .B1(_1797_),
    .B2(_1807_),
    .C1(_1658_),
    .X(_1808_));
 sky130_fd_sc_hd__o21ai_4 _6494_ (.A1(net61),
    .A2(_1709_),
    .B1(_1808_),
    .Y(_1809_));
 sky130_fd_sc_hd__and2b_1 _6495_ (.A_N(_1761_),
    .B(_1807_),
    .X(_1810_));
 sky130_fd_sc_hd__a211o_1 _6496_ (.A1(_1647_),
    .A2(_1741_),
    .B1(_1810_),
    .C1(_1658_),
    .X(_1811_));
 sky130_fd_sc_hd__o21ai_4 _6497_ (.A1(net61),
    .A2(_1697_),
    .B1(_1811_),
    .Y(_1812_));
 sky130_fd_sc_hd__nand3b_4 _6498_ (.A_N(_1806_),
    .B(_1809_),
    .C(_1812_),
    .Y(_1813_));
 sky130_fd_sc_hd__nor2_2 _6499_ (.A(_1801_),
    .B(_1813_),
    .Y(_1815_));
 sky130_fd_sc_hd__o21bai_4 _6500_ (.A1(_1795_),
    .A2(_1815_),
    .B1_N(_1796_),
    .Y(_1816_));
 sky130_fd_sc_hd__a21o_1 _6501_ (.A1(_1752_),
    .A2(_1753_),
    .B1(_1755_),
    .X(_1817_));
 sky130_fd_sc_hd__o21ai_4 _6502_ (.A1(_1794_),
    .A2(_1816_),
    .B1(_1817_),
    .Y(_1818_));
 sky130_fd_sc_hd__a21oi_4 _6503_ (.A1(_1793_),
    .A2(_1818_),
    .B1(_1791_),
    .Y(_1819_));
 sky130_fd_sc_hd__o21ai_4 _6504_ (.A1(_1790_),
    .A2(_1819_),
    .B1(_1788_),
    .Y(_1820_));
 sky130_fd_sc_hd__a21o_1 _6505_ (.A1(_1723_),
    .A2(_1820_),
    .B1(_1724_),
    .X(_1821_));
 sky130_fd_sc_hd__a21o_1 _6506_ (.A1(_1787_),
    .A2(_1821_),
    .B1(_1786_),
    .X(_1822_));
 sky130_fd_sc_hd__a21oi_1 _6507_ (.A1(_1701_),
    .A2(_1822_),
    .B1(_1702_),
    .Y(_1823_));
 sky130_fd_sc_hd__a221o_1 _6508_ (.A1(_1688_),
    .A2(_1689_),
    .B1(_1701_),
    .B2(_1822_),
    .C1(_1702_),
    .X(_1824_));
 sky130_fd_sc_hd__o21a_1 _6509_ (.A1(_1688_),
    .A2(_1689_),
    .B1(_1824_),
    .X(_1826_));
 sky130_fd_sc_hd__a21oi_1 _6510_ (.A1(_1677_),
    .A2(_1826_),
    .B1(_1678_),
    .Y(_1827_));
 sky130_fd_sc_hd__a21o_1 _6511_ (.A1(_1657_),
    .A2(_1665_),
    .B1(_1667_),
    .X(_1828_));
 sky130_fd_sc_hd__o211a_1 _6512_ (.A1(_1785_),
    .A2(_1827_),
    .B1(_1828_),
    .C1(net224),
    .X(_1829_));
 sky130_fd_sc_hd__o21bai_4 _6513_ (.A1(net224),
    .A2(_1782_),
    .B1_N(_1829_),
    .Y(_1830_));
 sky130_fd_sc_hd__xor2_4 _6514_ (.A(_1783_),
    .B(_1830_),
    .X(_1831_));
 sky130_fd_sc_hd__nand2b_2 _6515_ (.A_N(net44),
    .B(_1831_),
    .Y(_1832_));
 sky130_fd_sc_hd__mux2_4 _6516_ (.A0(_1779_),
    .A1(_1827_),
    .S(net224),
    .X(_1833_));
 sky130_fd_sc_hd__xnor2_4 _6517_ (.A(_1785_),
    .B(_1833_),
    .Y(_1834_));
 sky130_fd_sc_hd__nand2b_2 _6518_ (.A_N(_1832_),
    .B(_1834_),
    .Y(_1835_));
 sky130_fd_sc_hd__mux2_1 _6519_ (.A0(_1777_),
    .A1(_1823_),
    .S(net226),
    .X(_1837_));
 sky130_fd_sc_hd__xnor2_2 _6520_ (.A(_1691_),
    .B(_1837_),
    .Y(_1838_));
 sky130_fd_sc_hd__inv_2 _6521_ (.A(_1838_),
    .Y(_1839_));
 sky130_fd_sc_hd__mux2_4 _6522_ (.A0(_1778_),
    .A1(_1826_),
    .S(net224),
    .X(_1840_));
 sky130_fd_sc_hd__xnor2_4 _6523_ (.A(_1680_),
    .B(_1840_),
    .Y(_1841_));
 sky130_fd_sc_hd__or2_1 _6524_ (.A(_1839_),
    .B(_1841_),
    .X(_1842_));
 sky130_fd_sc_hd__or2_2 _6525_ (.A(_1835_),
    .B(_1842_),
    .X(_1843_));
 sky130_fd_sc_hd__mux2_4 _6526_ (.A0(_1775_),
    .A1(_1822_),
    .S(net226),
    .X(_1844_));
 sky130_fd_sc_hd__xnor2_4 _6527_ (.A(_1705_),
    .B(_1844_),
    .Y(_1845_));
 sky130_fd_sc_hd__mux2_4 _6528_ (.A0(_1774_),
    .A1(_1821_),
    .S(net226),
    .X(_1846_));
 sky130_fd_sc_hd__xor2_4 _6529_ (.A(_1787_),
    .B(_1846_),
    .X(_1848_));
 sky130_fd_sc_hd__nor2_1 _6530_ (.A(_1845_),
    .B(_1848_),
    .Y(_1849_));
 sky130_fd_sc_hd__nor2_1 _6531_ (.A(net226),
    .B(_1773_),
    .Y(_1850_));
 sky130_fd_sc_hd__a21oi_4 _6532_ (.A1(net226),
    .A2(_1820_),
    .B1(_1850_),
    .Y(_1851_));
 sky130_fd_sc_hd__xor2_4 _6533_ (.A(_1727_),
    .B(_1851_),
    .X(_1852_));
 sky130_fd_sc_hd__inv_2 _6534_ (.A(_1852_),
    .Y(_1853_));
 sky130_fd_sc_hd__mux2_4 _6535_ (.A0(_1772_),
    .A1(_1819_),
    .S(net226),
    .X(_1854_));
 sky130_fd_sc_hd__xnor2_4 _6536_ (.A(_1789_),
    .B(_1854_),
    .Y(_1855_));
 sky130_fd_sc_hd__inv_2 _6537_ (.A(_1855_),
    .Y(_1856_));
 sky130_fd_sc_hd__or2_1 _6538_ (.A(_1852_),
    .B(_1855_),
    .X(_1857_));
 sky130_fd_sc_hd__or3_1 _6539_ (.A(_1845_),
    .B(_1848_),
    .C(_1857_),
    .X(_1859_));
 sky130_fd_sc_hd__or2_4 _6540_ (.A(_1843_),
    .B(_1859_),
    .X(_1860_));
 sky130_fd_sc_hd__nor2_1 _6541_ (.A(net226),
    .B(_1769_),
    .Y(_1861_));
 sky130_fd_sc_hd__a21oi_4 _6542_ (.A1(net226),
    .A2(_1818_),
    .B1(_1861_),
    .Y(_1862_));
 sky130_fd_sc_hd__xor2_4 _6543_ (.A(_1793_),
    .B(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__mux2_4 _6544_ (.A0(_1768_),
    .A1(_1816_),
    .S(net226),
    .X(_1864_));
 sky130_fd_sc_hd__xor2_4 _6545_ (.A(_1794_),
    .B(_1864_),
    .X(_1865_));
 sky130_fd_sc_hd__inv_2 _6546_ (.A(_1865_),
    .Y(_1866_));
 sky130_fd_sc_hd__nand2_4 _6547_ (.A(_1863_),
    .B(_1866_),
    .Y(_1867_));
 sky130_fd_sc_hd__and2_2 _6548_ (.A(net225),
    .B(_1813_),
    .X(_1868_));
 sky130_fd_sc_hd__xnor2_4 _6549_ (.A(_1801_),
    .B(_1868_),
    .Y(_1870_));
 sky130_fd_sc_hd__or4_1 _6550_ (.A(net221),
    .B(_1795_),
    .C(_1796_),
    .D(_1815_),
    .X(_1871_));
 sky130_fd_sc_hd__o22ai_2 _6551_ (.A1(_1795_),
    .A2(_1796_),
    .B1(_1815_),
    .B2(net221),
    .Y(_1872_));
 sky130_fd_sc_hd__nand2_2 _6552_ (.A(_1871_),
    .B(_1872_),
    .Y(_1873_));
 sky130_fd_sc_hd__inv_2 _6553_ (.A(_1873_),
    .Y(_1874_));
 sky130_fd_sc_hd__nand2_4 _6554_ (.A(_1870_),
    .B(_1874_),
    .Y(_1875_));
 sky130_fd_sc_hd__nor2_4 _6555_ (.A(_1867_),
    .B(_1875_),
    .Y(_1876_));
 sky130_fd_sc_hd__nor2_8 _6556_ (.A(_1860_),
    .B(_1876_),
    .Y(_1877_));
 sky130_fd_sc_hd__or2_1 _6557_ (.A(_1589_),
    .B(_1877_),
    .X(_1878_));
 sky130_fd_sc_hd__nor2_1 _6558_ (.A(_1602_),
    .B(_1878_),
    .Y(_1879_));
 sky130_fd_sc_hd__and2_1 _6559_ (.A(_1602_),
    .B(_1878_),
    .X(_1881_));
 sky130_fd_sc_hd__nor2_1 _6560_ (.A(_1879_),
    .B(_1881_),
    .Y(_1882_));
 sky130_fd_sc_hd__a21oi_1 _6561_ (.A1(_1813_),
    .A2(_1876_),
    .B1(_1859_),
    .Y(_1883_));
 sky130_fd_sc_hd__nor2_1 _6562_ (.A(_1843_),
    .B(_1883_),
    .Y(_1884_));
 sky130_fd_sc_hd__or2_2 _6563_ (.A(_1615_),
    .B(net39),
    .X(_1885_));
 sky130_fd_sc_hd__nand2_1 _6564_ (.A(_1589_),
    .B(_1877_),
    .Y(_1886_));
 sky130_fd_sc_hd__and2_1 _6565_ (.A(_1878_),
    .B(_1886_),
    .X(_1887_));
 sky130_fd_sc_hd__and2b_1 _6566_ (.A_N(_1885_),
    .B(_1887_),
    .X(_1888_));
 sky130_fd_sc_hd__xnor2_1 _6567_ (.A(_1885_),
    .B(_1887_),
    .Y(_1889_));
 sky130_fd_sc_hd__a21oi_2 _6568_ (.A1(_1849_),
    .A2(_1857_),
    .B1(_1842_),
    .Y(_1890_));
 sky130_fd_sc_hd__a31o_2 _6569_ (.A1(_1804_),
    .A2(_1805_),
    .A3(_1809_),
    .B1(_1472_),
    .X(_1892_));
 sky130_fd_sc_hd__xnor2_4 _6570_ (.A(_1812_),
    .B(_1892_),
    .Y(_1893_));
 sky130_fd_sc_hd__nand2_2 _6571_ (.A(net224),
    .B(_1806_),
    .Y(_1894_));
 sky130_fd_sc_hd__xnor2_4 _6572_ (.A(_1809_),
    .B(_1894_),
    .Y(_1895_));
 sky130_fd_sc_hd__a31oi_4 _6573_ (.A1(_1806_),
    .A2(_1893_),
    .A3(_1895_),
    .B1(_1875_),
    .Y(_1896_));
 sky130_fd_sc_hd__o32ai_4 _6574_ (.A1(_1860_),
    .A2(_1867_),
    .A3(_1896_),
    .B1(_1890_),
    .B2(_1835_),
    .Y(_1897_));
 sky130_fd_sc_hd__mux2_8 _6575_ (.A0(_3435_),
    .A1(_1249_),
    .S(net97),
    .X(_1898_));
 sky130_fd_sc_hd__nand2b_1 _6576_ (.A_N(_1897_),
    .B(_1898_),
    .Y(_1899_));
 sky130_fd_sc_hd__nand2_1 _6577_ (.A(_1615_),
    .B(net39),
    .Y(_1900_));
 sky130_fd_sc_hd__nand2_1 _6578_ (.A(_1885_),
    .B(_1900_),
    .Y(_1901_));
 sky130_fd_sc_hd__nor2_1 _6579_ (.A(_1899_),
    .B(_1901_),
    .Y(_1903_));
 sky130_fd_sc_hd__xor2_4 _6580_ (.A(_1897_),
    .B(_1898_),
    .X(_1904_));
 sky130_fd_sc_hd__nor2_1 _6581_ (.A(_1870_),
    .B(_1873_),
    .Y(_1905_));
 sky130_fd_sc_hd__o21a_1 _6582_ (.A1(_1865_),
    .A2(_1905_),
    .B1(_1863_),
    .X(_1906_));
 sky130_fd_sc_hd__nor2_1 _6583_ (.A(_1472_),
    .B(_1805_),
    .Y(_1907_));
 sky130_fd_sc_hd__xnor2_1 _6584_ (.A(_1804_),
    .B(_1907_),
    .Y(_1908_));
 sky130_fd_sc_hd__o21a_1 _6585_ (.A1(_1838_),
    .A2(_1841_),
    .B1(_1834_),
    .X(_1909_));
 sky130_fd_sc_hd__a21oi_2 _6586_ (.A1(_1853_),
    .A2(_1855_),
    .B1(_1848_),
    .Y(_1910_));
 sky130_fd_sc_hd__o32ai_4 _6587_ (.A1(_1843_),
    .A2(_1845_),
    .A3(_1910_),
    .B1(_1909_),
    .B2(_1832_),
    .Y(_1911_));
 sky130_fd_sc_hd__mux2_8 _6588_ (.A0(_1906_),
    .A1(_1911_),
    .S(_1860_),
    .X(_1912_));
 sky130_fd_sc_hd__and2b_2 _6589_ (.A_N(_1609_),
    .B(_1912_),
    .X(_1914_));
 sky130_fd_sc_hd__xor2_2 _6590_ (.A(_1609_),
    .B(_1912_),
    .X(_1915_));
 sky130_fd_sc_hd__nand2_2 _6591_ (.A(_1784_),
    .B(_1915_),
    .Y(_1916_));
 sky130_fd_sc_hd__xnor2_4 _6592_ (.A(_1904_),
    .B(_1914_),
    .Y(_1917_));
 sky130_fd_sc_hd__o22a_1 _6593_ (.A1(_1904_),
    .A2(_1914_),
    .B1(_1916_),
    .B2(_1917_),
    .X(_1918_));
 sky130_fd_sc_hd__and2_1 _6594_ (.A(_1899_),
    .B(_1901_),
    .X(_1919_));
 sky130_fd_sc_hd__or2_1 _6595_ (.A(_1903_),
    .B(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__nor2_1 _6596_ (.A(_1918_),
    .B(_1920_),
    .Y(_1921_));
 sky130_fd_sc_hd__o21a_1 _6597_ (.A1(_1903_),
    .A2(_1921_),
    .B1(_1889_),
    .X(_1922_));
 sky130_fd_sc_hd__o21a_1 _6598_ (.A1(_1888_),
    .A2(_1922_),
    .B1(_1882_),
    .X(_1923_));
 sky130_fd_sc_hd__o21ai_2 _6599_ (.A1(_1879_),
    .A2(_1923_),
    .B1(_1604_),
    .Y(_1925_));
 sky130_fd_sc_hd__a21oi_2 _6600_ (.A1(_1603_),
    .A2(_1925_),
    .B1(_1599_),
    .Y(_1926_));
 sky130_fd_sc_hd__and3_1 _6601_ (.A(_1599_),
    .B(_1603_),
    .C(_1925_),
    .X(_1927_));
 sky130_fd_sc_hd__or2_2 _6602_ (.A(_1926_),
    .B(_1927_),
    .X(_1928_));
 sky130_fd_sc_hd__o22ai_4 _6603_ (.A1(_1332_),
    .A2(_1597_),
    .B1(_1598_),
    .B2(_1595_),
    .Y(_1929_));
 sky130_fd_sc_hd__o22ai_4 _6604_ (.A1(_1596_),
    .A2(_1597_),
    .B1(_1926_),
    .B2(_1929_),
    .Y(_1930_));
 sky130_fd_sc_hd__nor3_1 _6605_ (.A(_1889_),
    .B(_1903_),
    .C(_1921_),
    .Y(_1931_));
 sky130_fd_sc_hd__nor2_2 _6606_ (.A(_1922_),
    .B(_1931_),
    .Y(_1932_));
 sky130_fd_sc_hd__or2_1 _6607_ (.A(_1930_),
    .B(_1932_),
    .X(_1933_));
 sky130_fd_sc_hd__and2_1 _6608_ (.A(_1930_),
    .B(_1932_),
    .X(_1934_));
 sky130_fd_sc_hd__nand2_1 _6609_ (.A(_1930_),
    .B(_1932_),
    .Y(_1936_));
 sky130_fd_sc_hd__nand2_1 _6610_ (.A(_1933_),
    .B(_1936_),
    .Y(_1937_));
 sky130_fd_sc_hd__and2_1 _6611_ (.A(_1918_),
    .B(_1920_),
    .X(_1938_));
 sky130_fd_sc_hd__nor2_1 _6612_ (.A(_1921_),
    .B(_1938_),
    .Y(_1939_));
 sky130_fd_sc_hd__xor2_2 _6613_ (.A(_1916_),
    .B(_1917_),
    .X(_1940_));
 sky130_fd_sc_hd__or2_1 _6614_ (.A(_1784_),
    .B(_1915_),
    .X(_1941_));
 sky130_fd_sc_hd__and2_2 _6615_ (.A(_1916_),
    .B(_1941_),
    .X(_1942_));
 sky130_fd_sc_hd__or4_1 _6616_ (.A(_1932_),
    .B(_1939_),
    .C(_1940_),
    .D(_1942_),
    .X(_1943_));
 sky130_fd_sc_hd__nor3_1 _6617_ (.A(_1882_),
    .B(_1888_),
    .C(_1922_),
    .Y(_1944_));
 sky130_fd_sc_hd__or2_2 _6618_ (.A(_1923_),
    .B(_1944_),
    .X(_1945_));
 sky130_fd_sc_hd__inv_2 _6619_ (.A(_1945_),
    .Y(_1947_));
 sky130_fd_sc_hd__nand2_1 _6620_ (.A(_1932_),
    .B(_1945_),
    .Y(_1948_));
 sky130_fd_sc_hd__nor2_1 _6621_ (.A(_1932_),
    .B(_1945_),
    .Y(_1949_));
 sky130_fd_sc_hd__inv_2 _6622_ (.A(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__nand2_1 _6623_ (.A(_1948_),
    .B(_1950_),
    .Y(_1951_));
 sky130_fd_sc_hd__or3b_1 _6624_ (.A(net22),
    .B(net24),
    .C_N(_1943_),
    .X(_1952_));
 sky130_fd_sc_hd__o21ai_1 _6625_ (.A1(_1943_),
    .A2(_1947_),
    .B1(_1930_),
    .Y(_1953_));
 sky130_fd_sc_hd__or3_1 _6626_ (.A(_1604_),
    .B(_1879_),
    .C(_1923_),
    .X(_1954_));
 sky130_fd_sc_hd__and2_1 _6627_ (.A(_1925_),
    .B(_1954_),
    .X(_1955_));
 sky130_fd_sc_hd__xnor2_1 _6628_ (.A(_1953_),
    .B(_1955_),
    .Y(_1956_));
 sky130_fd_sc_hd__xnor2_1 _6629_ (.A(_1952_),
    .B(_1956_),
    .Y(_1958_));
 sky130_fd_sc_hd__clkinv_4 _6630_ (.A(net18),
    .Y(_1959_));
 sky130_fd_sc_hd__and2_1 _6631_ (.A(_1930_),
    .B(net19),
    .X(_1960_));
 sky130_fd_sc_hd__a21o_1 _6632_ (.A1(_1933_),
    .A2(_1947_),
    .B1(_1934_),
    .X(_1961_));
 sky130_fd_sc_hd__a21o_1 _6633_ (.A1(_1959_),
    .A2(_1961_),
    .B1(_1960_),
    .X(_1962_));
 sky130_fd_sc_hd__nand2_1 _6634_ (.A(_1928_),
    .B(_1962_),
    .Y(_1963_));
 sky130_fd_sc_hd__xnor2_2 _6635_ (.A(_1928_),
    .B(_1962_),
    .Y(_1964_));
 sky130_fd_sc_hd__clkinv_2 _6636_ (.A(net16),
    .Y(_1965_));
 sky130_fd_sc_hd__or2_2 _6637_ (.A(net23),
    .B(net18),
    .X(_1966_));
 sky130_fd_sc_hd__inv_2 _6638_ (.A(_1966_),
    .Y(_1967_));
 sky130_fd_sc_hd__o211a_1 _6639_ (.A1(net21),
    .A2(net18),
    .B1(net17),
    .C1(_1966_),
    .X(_1969_));
 sky130_fd_sc_hd__inv_2 _6640_ (.A(_1969_),
    .Y(_1970_));
 sky130_fd_sc_hd__or2_1 _6641_ (.A(_1877_),
    .B(net39),
    .X(_1971_));
 sky130_fd_sc_hd__mux2_1 _6642_ (.A0(_1863_),
    .A1(_1866_),
    .S(net34),
    .X(_1972_));
 sky130_fd_sc_hd__mux2_1 _6643_ (.A0(_1874_),
    .A1(_1870_),
    .S(net34),
    .X(_1973_));
 sky130_fd_sc_hd__mux2_1 _6644_ (.A0(_1972_),
    .A1(_1973_),
    .S(net37),
    .X(_1974_));
 sky130_fd_sc_hd__nor2_1 _6645_ (.A(_1971_),
    .B(_1974_),
    .Y(_1975_));
 sky130_fd_sc_hd__mux2_1 _6646_ (.A0(_1865_),
    .A1(_1873_),
    .S(net34),
    .X(_1976_));
 sky130_fd_sc_hd__inv_2 _6647_ (.A(_1976_),
    .Y(_1977_));
 sky130_fd_sc_hd__mux2_1 _6648_ (.A0(_1870_),
    .A1(_1893_),
    .S(net34),
    .X(_1978_));
 sky130_fd_sc_hd__mux2_1 _6649_ (.A0(_1977_),
    .A1(_1978_),
    .S(net36),
    .X(_1980_));
 sky130_fd_sc_hd__or2_1 _6650_ (.A(net38),
    .B(_1980_),
    .X(_1981_));
 sky130_fd_sc_hd__inv_2 _6651_ (.A(_1981_),
    .Y(_1982_));
 sky130_fd_sc_hd__nor2_1 _6652_ (.A(net44),
    .B(_1877_),
    .Y(_1983_));
 sky130_fd_sc_hd__a22o_1 _6653_ (.A1(net44),
    .A2(_1975_),
    .B1(_1982_),
    .B2(_1983_),
    .X(_1984_));
 sky130_fd_sc_hd__or2_1 _6654_ (.A(net36),
    .B(_1973_),
    .X(_1985_));
 sky130_fd_sc_hd__nor2_2 _6655_ (.A(net38),
    .B(_1985_),
    .Y(_1986_));
 sky130_fd_sc_hd__a22o_1 _6656_ (.A1(net44),
    .A2(_1982_),
    .B1(_1983_),
    .B2(_1986_),
    .X(_1987_));
 sky130_fd_sc_hd__mux2_1 _6657_ (.A0(_1987_),
    .A1(_1984_),
    .S(net20),
    .X(_1988_));
 sky130_fd_sc_hd__mux2_1 _6658_ (.A0(_1853_),
    .A1(_1856_),
    .S(net34),
    .X(_1989_));
 sky130_fd_sc_hd__and2b_1 _6659_ (.A_N(net36),
    .B(_1989_),
    .X(_1991_));
 sky130_fd_sc_hd__a21oi_2 _6660_ (.A1(net36),
    .A2(_1972_),
    .B1(_1991_),
    .Y(_1992_));
 sky130_fd_sc_hd__inv_2 _6661_ (.A(_1992_),
    .Y(_1993_));
 sky130_fd_sc_hd__mux2_1 _6662_ (.A0(_1993_),
    .A1(_1985_),
    .S(net38),
    .X(_1994_));
 sky130_fd_sc_hd__or2_2 _6663_ (.A(net36),
    .B(_1978_),
    .X(_1995_));
 sky130_fd_sc_hd__inv_2 _6664_ (.A(_1995_),
    .Y(_1996_));
 sky130_fd_sc_hd__mux2_1 _6665_ (.A0(_1856_),
    .A1(_1863_),
    .S(net35),
    .X(_1997_));
 sky130_fd_sc_hd__inv_2 _6666_ (.A(_1997_),
    .Y(_1998_));
 sky130_fd_sc_hd__mux2_1 _6667_ (.A0(_1998_),
    .A1(_1976_),
    .S(net36),
    .X(_1999_));
 sky130_fd_sc_hd__mux2_1 _6668_ (.A0(_1999_),
    .A1(_1996_),
    .S(net38),
    .X(_2000_));
 sky130_fd_sc_hd__inv_2 _6669_ (.A(_2000_),
    .Y(_2002_));
 sky130_fd_sc_hd__mux2_1 _6670_ (.A0(_2002_),
    .A1(_1994_),
    .S(net45),
    .X(_2003_));
 sky130_fd_sc_hd__mux2_1 _6671_ (.A0(_1975_),
    .A1(_2000_),
    .S(net44),
    .X(_2004_));
 sky130_fd_sc_hd__inv_2 _6672_ (.A(_2004_),
    .Y(_2005_));
 sky130_fd_sc_hd__mux2_1 _6673_ (.A0(_2005_),
    .A1(_2003_),
    .S(net20),
    .X(_2006_));
 sky130_fd_sc_hd__inv_2 _6674_ (.A(_2006_),
    .Y(_2007_));
 sky130_fd_sc_hd__and2_1 _6675_ (.A(net23),
    .B(_2007_),
    .X(_2008_));
 sky130_fd_sc_hd__mux2_1 _6676_ (.A0(_1848_),
    .A1(_1852_),
    .S(net34),
    .X(_2009_));
 sky130_fd_sc_hd__inv_2 _6677_ (.A(_2009_),
    .Y(_2010_));
 sky130_fd_sc_hd__mux2_1 _6678_ (.A0(_2010_),
    .A1(_1997_),
    .S(net37),
    .X(_2011_));
 sky130_fd_sc_hd__and2b_1 _6679_ (.A_N(net38),
    .B(_2011_),
    .X(_2013_));
 sky130_fd_sc_hd__a21oi_1 _6680_ (.A1(net39),
    .A2(_1980_),
    .B1(_2013_),
    .Y(_2014_));
 sky130_fd_sc_hd__nand2_1 _6681_ (.A(net45),
    .B(_2014_),
    .Y(_2015_));
 sky130_fd_sc_hd__o21ai_1 _6682_ (.A1(net44),
    .A2(_1994_),
    .B1(_2015_),
    .Y(_2016_));
 sky130_fd_sc_hd__mux2_1 _6683_ (.A0(_1845_),
    .A1(_1848_),
    .S(net34),
    .X(_2017_));
 sky130_fd_sc_hd__a2bb2o_1 _6684_ (.A1_N(net37),
    .A2_N(_2017_),
    .B1(_1974_),
    .B2(net38),
    .X(_2018_));
 sky130_fd_sc_hd__a21oi_1 _6685_ (.A1(net37),
    .A2(_1989_),
    .B1(_2018_),
    .Y(_2019_));
 sky130_fd_sc_hd__mux2_1 _6686_ (.A0(_2014_),
    .A1(_2019_),
    .S(net45),
    .X(_2020_));
 sky130_fd_sc_hd__mux2_1 _6687_ (.A0(_2016_),
    .A1(_2020_),
    .S(net21),
    .X(_2021_));
 sky130_fd_sc_hd__mux2_1 _6688_ (.A0(_1839_),
    .A1(_1845_),
    .S(net34),
    .X(_2022_));
 sky130_fd_sc_hd__mux2_1 _6689_ (.A0(_2022_),
    .A1(_2009_),
    .S(net36),
    .X(_2024_));
 sky130_fd_sc_hd__mux2_1 _6690_ (.A0(_2024_),
    .A1(_1999_),
    .S(net38),
    .X(_2025_));
 sky130_fd_sc_hd__nor2_2 _6691_ (.A(net39),
    .B(_1995_),
    .Y(_2026_));
 sky130_fd_sc_hd__a21o_1 _6692_ (.A1(_1877_),
    .A2(_2026_),
    .B1(_2025_),
    .X(_2027_));
 sky130_fd_sc_hd__mux2_1 _6693_ (.A0(_2019_),
    .A1(_2027_),
    .S(net45),
    .X(_2028_));
 sky130_fd_sc_hd__mux2_1 _6694_ (.A0(_1841_),
    .A1(_1839_),
    .S(net35),
    .X(_2029_));
 sky130_fd_sc_hd__mux2_1 _6695_ (.A0(_2029_),
    .A1(_2017_),
    .S(net36),
    .X(_2030_));
 sky130_fd_sc_hd__a21o_1 _6696_ (.A1(net38),
    .A2(_1992_),
    .B1(_2030_),
    .X(_2031_));
 sky130_fd_sc_hd__mux2_1 _6697_ (.A0(_2031_),
    .A1(_1986_),
    .S(_1877_),
    .X(_2032_));
 sky130_fd_sc_hd__mux2_1 _6698_ (.A0(_2027_),
    .A1(_2032_),
    .S(net44),
    .X(_2033_));
 sky130_fd_sc_hd__mux2_1 _6699_ (.A0(_2028_),
    .A1(_2033_),
    .S(net20),
    .X(_2035_));
 sky130_fd_sc_hd__mux2_1 _6700_ (.A0(_2021_),
    .A1(_2035_),
    .S(net23),
    .X(_2036_));
 sky130_fd_sc_hd__and2_1 _6701_ (.A(net18),
    .B(_2036_),
    .X(_2037_));
 sky130_fd_sc_hd__a221o_1 _6702_ (.A1(_1967_),
    .A2(_1988_),
    .B1(_2008_),
    .B2(_1959_),
    .C1(_2037_),
    .X(_2038_));
 sky130_fd_sc_hd__mux2_1 _6703_ (.A0(_1984_),
    .A1(_2004_),
    .S(net20),
    .X(_2039_));
 sky130_fd_sc_hd__nand2_1 _6704_ (.A(net20),
    .B(_2016_),
    .Y(_2040_));
 sky130_fd_sc_hd__o21a_1 _6705_ (.A1(net21),
    .A2(_2003_),
    .B1(_2040_),
    .X(_2041_));
 sky130_fd_sc_hd__inv_2 _6706_ (.A(_2041_),
    .Y(_2042_));
 sky130_fd_sc_hd__and2_1 _6707_ (.A(net23),
    .B(_2042_),
    .X(_2043_));
 sky130_fd_sc_hd__mux2_1 _6708_ (.A0(_2020_),
    .A1(_2028_),
    .S(net21),
    .X(_2044_));
 sky130_fd_sc_hd__nor2_1 _6709_ (.A(_1834_),
    .B(net34),
    .Y(_2046_));
 sky130_fd_sc_hd__a221o_1 _6710_ (.A1(_1841_),
    .A2(net34),
    .B1(_2022_),
    .B2(net36),
    .C1(net38),
    .X(_2047_));
 sky130_fd_sc_hd__a2bb2o_1 _6711_ (.A1_N(_2046_),
    .A2_N(_2047_),
    .B1(net38),
    .B2(_2011_),
    .X(_2048_));
 sky130_fd_sc_hd__a21bo_1 _6712_ (.A1(_1877_),
    .A2(_1982_),
    .B1_N(_2048_),
    .X(_2049_));
 sky130_fd_sc_hd__mux2_1 _6713_ (.A0(_2032_),
    .A1(_2049_),
    .S(net44),
    .X(_2050_));
 sky130_fd_sc_hd__mux2_1 _6714_ (.A0(_2033_),
    .A1(_2050_),
    .S(net20),
    .X(_2051_));
 sky130_fd_sc_hd__mux2_1 _6715_ (.A0(_2044_),
    .A1(_2051_),
    .S(net23),
    .X(_2052_));
 sky130_fd_sc_hd__and2_1 _6716_ (.A(net18),
    .B(_2052_),
    .X(_2053_));
 sky130_fd_sc_hd__a221o_1 _6717_ (.A1(_1967_),
    .A2(_2039_),
    .B1(_2043_),
    .B2(_1959_),
    .C1(_2053_),
    .X(_2054_));
 sky130_fd_sc_hd__mux2_1 _6718_ (.A0(_1831_),
    .A1(_1834_),
    .S(net35),
    .X(_2055_));
 sky130_fd_sc_hd__inv_2 _6719_ (.A(_2055_),
    .Y(_2057_));
 sky130_fd_sc_hd__a211o_4 _6720_ (.A1(net36),
    .A2(_2029_),
    .B1(_2057_),
    .C1(_1971_),
    .X(_2058_));
 sky130_fd_sc_hd__mux2_1 _6721_ (.A0(_2049_),
    .A1(_2058_),
    .S(net44),
    .X(_2059_));
 sky130_fd_sc_hd__mux2_1 _6722_ (.A0(_2059_),
    .A1(_1942_),
    .S(net22),
    .X(_2060_));
 sky130_fd_sc_hd__mux2_1 _6723_ (.A0(_1940_),
    .A1(_1939_),
    .S(net22),
    .X(_2061_));
 sky130_fd_sc_hd__mux2_1 _6724_ (.A0(_2060_),
    .A1(_2061_),
    .S(net24),
    .X(_2062_));
 sky130_fd_sc_hd__inv_2 _6725_ (.A(_2062_),
    .Y(_2063_));
 sky130_fd_sc_hd__mux2_1 _6726_ (.A0(_2052_),
    .A1(_2062_),
    .S(net18),
    .X(_2064_));
 sky130_fd_sc_hd__mux2_1 _6727_ (.A0(_2007_),
    .A1(_2021_),
    .S(net23),
    .X(_2065_));
 sky130_fd_sc_hd__mux2_2 _6728_ (.A0(_2050_),
    .A1(_2059_),
    .S(net20),
    .X(_2066_));
 sky130_fd_sc_hd__mux2_1 _6729_ (.A0(_2035_),
    .A1(_2066_),
    .S(net23),
    .X(_2068_));
 sky130_fd_sc_hd__inv_2 _6730_ (.A(_2068_),
    .Y(_2069_));
 sky130_fd_sc_hd__mux2_1 _6731_ (.A0(_2065_),
    .A1(_2068_),
    .S(net18),
    .X(_2070_));
 sky130_fd_sc_hd__or4_1 _6732_ (.A(_2038_),
    .B(_2054_),
    .C(_2064_),
    .D(_2070_),
    .X(_2071_));
 sky130_fd_sc_hd__mux2_1 _6733_ (.A0(_1942_),
    .A1(_1940_),
    .S(net22),
    .X(_2072_));
 sky130_fd_sc_hd__inv_2 _6734_ (.A(_2072_),
    .Y(_2073_));
 sky130_fd_sc_hd__mux2_1 _6735_ (.A0(_2066_),
    .A1(_2072_),
    .S(net24),
    .X(_2074_));
 sky130_fd_sc_hd__mux2_1 _6736_ (.A0(_2036_),
    .A1(_2074_),
    .S(net19),
    .X(_2075_));
 sky130_fd_sc_hd__nand2b_1 _6737_ (.A_N(_1895_),
    .B(net35),
    .Y(_2076_));
 sky130_fd_sc_hd__o21ai_1 _6738_ (.A1(_1893_),
    .A2(net35),
    .B1(_2076_),
    .Y(_2077_));
 sky130_fd_sc_hd__mux2_1 _6739_ (.A0(_2077_),
    .A1(_2026_),
    .S(net45),
    .X(_2079_));
 sky130_fd_sc_hd__a22o_1 _6740_ (.A1(net44),
    .A2(_1986_),
    .B1(_2026_),
    .B2(_1983_),
    .X(_2080_));
 sky130_fd_sc_hd__mux2_1 _6741_ (.A0(_2079_),
    .A1(_2080_),
    .S(net20),
    .X(_2081_));
 sky130_fd_sc_hd__mux2_1 _6742_ (.A0(_2081_),
    .A1(_1988_),
    .S(net23),
    .X(_2082_));
 sky130_fd_sc_hd__mux2_1 _6743_ (.A0(_2065_),
    .A1(_2082_),
    .S(_1959_),
    .X(_2083_));
 sky130_fd_sc_hd__inv_2 _6744_ (.A(_2083_),
    .Y(_2084_));
 sky130_fd_sc_hd__mux2_1 _6745_ (.A0(_2042_),
    .A1(_2044_),
    .S(net24),
    .X(_2085_));
 sky130_fd_sc_hd__mux2_1 _6746_ (.A0(_2051_),
    .A1(_2060_),
    .S(net23),
    .X(_2086_));
 sky130_fd_sc_hd__mux2_1 _6747_ (.A0(_2085_),
    .A1(_2086_),
    .S(net18),
    .X(_2087_));
 sky130_fd_sc_hd__a21o_1 _6748_ (.A1(_1948_),
    .A2(_2061_),
    .B1(_1949_),
    .X(_2088_));
 sky130_fd_sc_hd__mux2_1 _6749_ (.A0(_2086_),
    .A1(_2088_),
    .S(net18),
    .X(_2090_));
 sky130_fd_sc_hd__o41a_1 _6750_ (.A1(_1988_),
    .A2(_2008_),
    .A3(_2039_),
    .A4(_2043_),
    .B1(net18),
    .X(_2091_));
 sky130_fd_sc_hd__mux2_1 _6751_ (.A0(_2080_),
    .A1(_1987_),
    .S(net20),
    .X(_2092_));
 sky130_fd_sc_hd__o31a_1 _6752_ (.A1(_2081_),
    .A2(_2091_),
    .A3(_2092_),
    .B1(_1966_),
    .X(_2093_));
 sky130_fd_sc_hd__mux2_1 _6753_ (.A0(_2092_),
    .A1(_2039_),
    .S(net23),
    .X(_2094_));
 sky130_fd_sc_hd__mux2_1 _6754_ (.A0(_2085_),
    .A1(_2094_),
    .S(_1959_),
    .X(_2095_));
 sky130_fd_sc_hd__a221o_1 _6755_ (.A1(net45),
    .A2(_2077_),
    .B1(_2079_),
    .B2(net20),
    .C1(_1908_),
    .X(_2096_));
 sky130_fd_sc_hd__o21ba_1 _6756_ (.A1(_1895_),
    .A2(net35),
    .B1_N(_2096_),
    .X(_2097_));
 sky130_fd_sc_hd__or4_1 _6757_ (.A(_2075_),
    .B(_2083_),
    .C(_2087_),
    .D(_2095_),
    .X(_2098_));
 sky130_fd_sc_hd__o21a_1 _6758_ (.A1(_2071_),
    .A2(_2098_),
    .B1(net17),
    .X(_2099_));
 sky130_fd_sc_hd__mux2_2 _6759_ (.A0(_2095_),
    .A1(_2090_),
    .S(net17),
    .X(_2101_));
 sky130_fd_sc_hd__or4b_1 _6760_ (.A(_2093_),
    .B(_2099_),
    .C(_2101_),
    .D_N(_2097_),
    .X(_2102_));
 sky130_fd_sc_hd__o21ai_1 _6761_ (.A1(_1934_),
    .A2(_1939_),
    .B1(_1933_),
    .Y(_2103_));
 sky130_fd_sc_hd__mux2_1 _6762_ (.A0(_2073_),
    .A1(_2103_),
    .S(net24),
    .X(_2104_));
 sky130_fd_sc_hd__mux2_1 _6763_ (.A0(_2069_),
    .A1(_2104_),
    .S(net19),
    .X(_2105_));
 sky130_fd_sc_hd__mux2_2 _6764_ (.A0(_2084_),
    .A1(_2105_),
    .S(net17),
    .X(_2106_));
 sky130_fd_sc_hd__a21o_1 _6765_ (.A1(_1970_),
    .A2(_2102_),
    .B1(_2106_),
    .X(_2107_));
 sky130_fd_sc_hd__mux2_2 _6766_ (.A0(_0668_),
    .A1(_0646_),
    .S(net97),
    .X(_2108_));
 sky130_fd_sc_hd__mux2_8 _6767_ (.A0(net231),
    .A1(net234),
    .S(net98),
    .X(_2109_));
 sky130_fd_sc_hd__xor2_1 _6768_ (.A(_2101_),
    .B(_2106_),
    .X(_2110_));
 sky130_fd_sc_hd__o21ai_1 _6769_ (.A1(_2107_),
    .A2(_2109_),
    .B1(_2110_),
    .Y(_2112_));
 sky130_fd_sc_hd__nand2_1 _6770_ (.A(net231),
    .B(net212),
    .Y(_2113_));
 sky130_fd_sc_hd__o21a_2 _6771_ (.A1(_0646_),
    .A2(_0333_),
    .B1(_2113_),
    .X(_2114_));
 sky130_fd_sc_hd__o21ai_4 _6772_ (.A1(_1784_),
    .A2(_2058_),
    .B1(_2114_),
    .Y(_2115_));
 sky130_fd_sc_hd__nor3_4 _6773_ (.A(\cmd[7] ),
    .B(\cmd[6] ),
    .C(_2115_),
    .Y(_2116_));
 sky130_fd_sc_hd__or3_4 _6774_ (.A(\cmd[7] ),
    .B(\cmd[6] ),
    .C(_2115_),
    .X(_2117_));
 sky130_fd_sc_hd__o31a_1 _6775_ (.A1(_2101_),
    .A2(_2107_),
    .A3(_2109_),
    .B1(_2116_),
    .X(_2118_));
 sky130_fd_sc_hd__nand2_1 _6776_ (.A(_2112_),
    .B(_2118_),
    .Y(_2119_));
 sky130_fd_sc_hd__nand2_4 _6777_ (.A(net163),
    .B(net64),
    .Y(_2120_));
 sky130_fd_sc_hd__or2_4 _6778_ (.A(_3476_),
    .B(net86),
    .X(_2121_));
 sky130_fd_sc_hd__nand2_2 _6779_ (.A(net128),
    .B(net87),
    .Y(_2123_));
 sky130_fd_sc_hd__nand2_1 _6780_ (.A(_0367_),
    .B(_2123_),
    .Y(_2124_));
 sky130_fd_sc_hd__o21ai_4 _6781_ (.A1(_0355_),
    .A2(_2121_),
    .B1(_2124_),
    .Y(_2125_));
 sky130_fd_sc_hd__xor2_4 _6782_ (.A(_2120_),
    .B(_2125_),
    .X(_2126_));
 sky130_fd_sc_hd__xnor2_2 _6783_ (.A(_0375_),
    .B(_2121_),
    .Y(_2127_));
 sky130_fd_sc_hd__and3_2 _6784_ (.A(net163),
    .B(net87),
    .C(_2127_),
    .X(_2128_));
 sky130_fd_sc_hd__o21ba_2 _6785_ (.A1(_0376_),
    .A2(_2121_),
    .B1_N(_2128_),
    .X(_2129_));
 sky130_fd_sc_hd__and2b_1 _6786_ (.A_N(_2129_),
    .B(_2126_),
    .X(_2130_));
 sky130_fd_sc_hd__nor2_1 _6787_ (.A(net69),
    .B(net161),
    .Y(_2131_));
 sky130_fd_sc_hd__xnor2_2 _6788_ (.A(_2126_),
    .B(_2129_),
    .Y(_2132_));
 sky130_fd_sc_hd__and2_1 _6789_ (.A(_2131_),
    .B(_2132_),
    .X(_2134_));
 sky130_fd_sc_hd__nor2_1 _6790_ (.A(net69),
    .B(net166),
    .Y(_2135_));
 sky130_fd_sc_hd__nor2_2 _6791_ (.A(net67),
    .B(_2123_),
    .Y(_2136_));
 sky130_fd_sc_hd__a21oi_1 _6792_ (.A1(net128),
    .A2(net65),
    .B1(_0354_),
    .Y(_2137_));
 sky130_fd_sc_hd__nor2_1 _6793_ (.A(_2136_),
    .B(_2137_),
    .Y(_2138_));
 sky130_fd_sc_hd__and2_1 _6794_ (.A(_2135_),
    .B(_2138_),
    .X(_2139_));
 sky130_fd_sc_hd__xnor2_1 _6795_ (.A(_2135_),
    .B(_2138_),
    .Y(_2140_));
 sky130_fd_sc_hd__o22a_1 _6796_ (.A1(_0367_),
    .A2(_2123_),
    .B1(_2125_),
    .B2(_2120_),
    .X(_2141_));
 sky130_fd_sc_hd__or2_1 _6797_ (.A(_2140_),
    .B(_2141_),
    .X(_2142_));
 sky130_fd_sc_hd__nand2_1 _6798_ (.A(_2140_),
    .B(_2141_),
    .Y(_2143_));
 sky130_fd_sc_hd__nand2_1 _6799_ (.A(_2142_),
    .B(_2143_),
    .Y(_2145_));
 sky130_fd_sc_hd__or3_2 _6800_ (.A(net161),
    .B(net202),
    .C(_2145_),
    .X(_2146_));
 sky130_fd_sc_hd__o21ai_1 _6801_ (.A1(net161),
    .A2(net201),
    .B1(_2145_),
    .Y(_2147_));
 sky130_fd_sc_hd__and2_1 _6802_ (.A(_2146_),
    .B(_2147_),
    .X(_2148_));
 sky130_fd_sc_hd__o21a_1 _6803_ (.A1(_2130_),
    .A2(_2134_),
    .B1(_2148_),
    .X(_2149_));
 sky130_fd_sc_hd__nand2_1 _6804_ (.A(_2142_),
    .B(_2146_),
    .Y(_2150_));
 sky130_fd_sc_hd__nor2_1 _6805_ (.A(net166),
    .B(net201),
    .Y(_2151_));
 sky130_fd_sc_hd__nor2_2 _6806_ (.A(net69),
    .B(net127),
    .Y(_2152_));
 sky130_fd_sc_hd__xnor2_1 _6807_ (.A(_0353_),
    .B(_2152_),
    .Y(_2153_));
 sky130_fd_sc_hd__nand2_2 _6808_ (.A(_2151_),
    .B(_2153_),
    .Y(_2154_));
 sky130_fd_sc_hd__or2_1 _6809_ (.A(_2151_),
    .B(_2153_),
    .X(_2156_));
 sky130_fd_sc_hd__and2_2 _6810_ (.A(_2154_),
    .B(_2156_),
    .X(_2157_));
 sky130_fd_sc_hd__o21ai_4 _6811_ (.A1(_2136_),
    .A2(_2139_),
    .B1(_2157_),
    .Y(_2158_));
 sky130_fd_sc_hd__or3_1 _6812_ (.A(_2136_),
    .B(_2139_),
    .C(_2157_),
    .X(_2159_));
 sky130_fd_sc_hd__nand2_2 _6813_ (.A(_2158_),
    .B(_2159_),
    .Y(_2160_));
 sky130_fd_sc_hd__a21o_1 _6814_ (.A1(_2142_),
    .A2(_2146_),
    .B1(_2160_),
    .X(_2161_));
 sky130_fd_sc_hd__xnor2_2 _6815_ (.A(_2150_),
    .B(_2160_),
    .Y(_2162_));
 sky130_fd_sc_hd__nand2_2 _6816_ (.A(_2149_),
    .B(_2162_),
    .Y(_2163_));
 sky130_fd_sc_hd__o31a_4 _6817_ (.A1(net69),
    .A2(net127),
    .A3(_0353_),
    .B1(_2154_),
    .X(_2164_));
 sky130_fd_sc_hd__o21a_1 _6818_ (.A1(net127),
    .A2(net201),
    .B1(_0390_),
    .X(_2165_));
 sky130_fd_sc_hd__or2_4 _6819_ (.A(_2152_),
    .B(_2165_),
    .X(_2167_));
 sky130_fd_sc_hd__xnor2_4 _6820_ (.A(_2164_),
    .B(_2167_),
    .Y(_2168_));
 sky130_fd_sc_hd__nand2_2 _6821_ (.A(_2158_),
    .B(_2161_),
    .Y(_2169_));
 sky130_fd_sc_hd__xor2_4 _6822_ (.A(_2168_),
    .B(_2169_),
    .X(_2170_));
 sky130_fd_sc_hd__nor2_1 _6823_ (.A(_2163_),
    .B(_2170_),
    .Y(_2171_));
 sky130_fd_sc_hd__or2_1 _6824_ (.A(_2161_),
    .B(_2168_),
    .X(_2172_));
 sky130_fd_sc_hd__o21bai_2 _6825_ (.A1(_2154_),
    .A2(_2165_),
    .B1_N(_2152_),
    .Y(_2173_));
 sky130_fd_sc_hd__o21a_1 _6826_ (.A1(_1216_),
    .A2(_2173_),
    .B1(_2158_),
    .X(_2174_));
 sky130_fd_sc_hd__nor3_1 _6827_ (.A(_1216_),
    .B(_2158_),
    .C(_2173_),
    .Y(_2175_));
 sky130_fd_sc_hd__nor2_1 _6828_ (.A(_2172_),
    .B(_2174_),
    .Y(_2176_));
 sky130_fd_sc_hd__o21a_1 _6829_ (.A1(_2174_),
    .A2(_2175_),
    .B1(_2172_),
    .X(_2178_));
 sky130_fd_sc_hd__nor2_1 _6830_ (.A(_2176_),
    .B(_2178_),
    .Y(_2179_));
 sky130_fd_sc_hd__xor2_1 _6831_ (.A(_2171_),
    .B(_2179_),
    .X(_2180_));
 sky130_fd_sc_hd__or2_1 _6832_ (.A(_2149_),
    .B(_2162_),
    .X(_2181_));
 sky130_fd_sc_hd__and2_2 _6833_ (.A(_2163_),
    .B(_2181_),
    .X(_2182_));
 sky130_fd_sc_hd__nor3_1 _6834_ (.A(_2130_),
    .B(_2134_),
    .C(_2148_),
    .Y(_2183_));
 sky130_fd_sc_hd__or2_1 _6835_ (.A(_2149_),
    .B(_2183_),
    .X(_2184_));
 sky130_fd_sc_hd__xnor2_1 _6836_ (.A(_2131_),
    .B(_2132_),
    .Y(_2185_));
 sky130_fd_sc_hd__a21oi_2 _6837_ (.A1(net163),
    .A2(net87),
    .B1(_2127_),
    .Y(_2186_));
 sky130_fd_sc_hd__nor2_4 _6838_ (.A(_2128_),
    .B(_2186_),
    .Y(_2187_));
 sky130_fd_sc_hd__or3_2 _6839_ (.A(net127),
    .B(net81),
    .C(_0433_),
    .X(_2189_));
 sky130_fd_sc_hd__o21ai_1 _6840_ (.A1(net127),
    .A2(net81),
    .B1(_0433_),
    .Y(_2190_));
 sky130_fd_sc_hd__nand2_1 _6841_ (.A(_2189_),
    .B(_2190_),
    .Y(_2191_));
 sky130_fd_sc_hd__or3_2 _6842_ (.A(net166),
    .B(net85),
    .C(_2191_),
    .X(_2192_));
 sky130_fd_sc_hd__nand2_2 _6843_ (.A(_2189_),
    .B(_2192_),
    .Y(_2193_));
 sky130_fd_sc_hd__nand2_4 _6844_ (.A(net157),
    .B(net64),
    .Y(_2194_));
 sky130_fd_sc_hd__xor2_4 _6845_ (.A(_2187_),
    .B(_2193_),
    .X(_2195_));
 sky130_fd_sc_hd__inv_2 _6846_ (.A(_2195_),
    .Y(_2196_));
 sky130_fd_sc_hd__o2bb2a_1 _6847_ (.A1_N(_2187_),
    .A2_N(_2193_),
    .B1(_2194_),
    .B2(_2196_),
    .X(_2197_));
 sky130_fd_sc_hd__nor2_2 _6848_ (.A(_2185_),
    .B(_2197_),
    .Y(_2198_));
 sky130_fd_sc_hd__and2_1 _6849_ (.A(_2185_),
    .B(_2197_),
    .X(_2200_));
 sky130_fd_sc_hd__or2_4 _6850_ (.A(_2198_),
    .B(_2200_),
    .X(_2201_));
 sky130_fd_sc_hd__or2_4 _6851_ (.A(net71),
    .B(net144),
    .X(_2202_));
 sky130_fd_sc_hd__and3_2 _6852_ (.A(net154),
    .B(net199),
    .C(_2202_),
    .X(_2203_));
 sky130_fd_sc_hd__nand2b_1 _6853_ (.A_N(_2201_),
    .B(_2203_),
    .Y(_2204_));
 sky130_fd_sc_hd__or2_4 _6854_ (.A(net71),
    .B(net149),
    .X(_2205_));
 sky130_fd_sc_hd__or3_2 _6855_ (.A(net144),
    .B(net200),
    .C(_2205_),
    .X(_2206_));
 sky130_fd_sc_hd__a21oi_2 _6856_ (.A1(_2204_),
    .A2(_2206_),
    .B1(_2184_),
    .Y(_2207_));
 sky130_fd_sc_hd__and3_1 _6857_ (.A(_2184_),
    .B(_2204_),
    .C(_2206_),
    .X(_2208_));
 sky130_fd_sc_hd__nor2_2 _6858_ (.A(_2207_),
    .B(_2208_),
    .Y(_2209_));
 sky130_fd_sc_hd__a21o_2 _6859_ (.A1(_2198_),
    .A2(_2209_),
    .B1(_2207_),
    .X(_2211_));
 sky130_fd_sc_hd__nand2_2 _6860_ (.A(_2182_),
    .B(_2211_),
    .Y(_2212_));
 sky130_fd_sc_hd__xnor2_2 _6861_ (.A(_2182_),
    .B(_2211_),
    .Y(_2213_));
 sky130_fd_sc_hd__xnor2_2 _6862_ (.A(_2198_),
    .B(_2209_),
    .Y(_2214_));
 sky130_fd_sc_hd__xor2_4 _6863_ (.A(_2201_),
    .B(_2203_),
    .X(_2215_));
 sky130_fd_sc_hd__and4_4 _6864_ (.A(net154),
    .B(_3496_),
    .C(net88),
    .D(net199),
    .X(_2216_));
 sky130_fd_sc_hd__nand2_4 _6865_ (.A(net64),
    .B(_2216_),
    .Y(_2217_));
 sky130_fd_sc_hd__xnor2_4 _6866_ (.A(_2194_),
    .B(_2195_),
    .Y(_2218_));
 sky130_fd_sc_hd__nand2b_1 _6867_ (.A_N(_2217_),
    .B(_2218_),
    .Y(_2219_));
 sky130_fd_sc_hd__xnor2_4 _6868_ (.A(_2217_),
    .B(_2218_),
    .Y(_2220_));
 sky130_fd_sc_hd__o21ai_1 _6869_ (.A1(net166),
    .A2(net85),
    .B1(_2191_),
    .Y(_2222_));
 sky130_fd_sc_hd__nand2_1 _6870_ (.A(_2192_),
    .B(_2222_),
    .Y(_2223_));
 sky130_fd_sc_hd__or3_2 _6871_ (.A(net127),
    .B(_0433_),
    .C(_0498_),
    .X(_2224_));
 sky130_fd_sc_hd__inv_2 _6872_ (.A(_2224_),
    .Y(_2225_));
 sky130_fd_sc_hd__nand2_4 _6873_ (.A(net163),
    .B(_0372_),
    .Y(_2226_));
 sky130_fd_sc_hd__a21oi_2 _6874_ (.A1(net128),
    .A2(net80),
    .B1(_0500_),
    .Y(_2227_));
 sky130_fd_sc_hd__nor2_2 _6875_ (.A(_2225_),
    .B(_2227_),
    .Y(_2228_));
 sky130_fd_sc_hd__o21a_1 _6876_ (.A1(_2226_),
    .A2(_2227_),
    .B1(_2224_),
    .X(_2229_));
 sky130_fd_sc_hd__xnor2_1 _6877_ (.A(_2223_),
    .B(_2229_),
    .Y(_2230_));
 sky130_fd_sc_hd__and3b_1 _6878_ (.A_N(_2230_),
    .B(net87),
    .C(net157),
    .X(_2231_));
 sky130_fd_sc_hd__o21ba_1 _6879_ (.A1(_2223_),
    .A2(_2229_),
    .B1_N(_2231_),
    .X(_2233_));
 sky130_fd_sc_hd__nand2b_1 _6880_ (.A_N(_2233_),
    .B(_2220_),
    .Y(_2234_));
 sky130_fd_sc_hd__xnor2_2 _6881_ (.A(_2220_),
    .B(_2233_),
    .Y(_2235_));
 sky130_fd_sc_hd__o21ai_1 _6882_ (.A1(net144),
    .A2(net200),
    .B1(_2205_),
    .Y(_2236_));
 sky130_fd_sc_hd__a21o_1 _6883_ (.A1(net154),
    .A2(net64),
    .B1(_2216_),
    .X(_2237_));
 sky130_fd_sc_hd__nand2_1 _6884_ (.A(_2217_),
    .B(_2237_),
    .Y(_2238_));
 sky130_fd_sc_hd__o2bb2a_1 _6885_ (.A1_N(_2206_),
    .A2_N(_2236_),
    .B1(_2238_),
    .B2(_2202_),
    .X(_2239_));
 sky130_fd_sc_hd__nand2b_2 _6886_ (.A_N(_2239_),
    .B(_2235_),
    .Y(_2240_));
 sky130_fd_sc_hd__and2_1 _6887_ (.A(_2219_),
    .B(_2234_),
    .X(_2241_));
 sky130_fd_sc_hd__xnor2_1 _6888_ (.A(_2215_),
    .B(_2240_),
    .Y(_2242_));
 sky130_fd_sc_hd__or2_1 _6889_ (.A(_2241_),
    .B(_2242_),
    .X(_2244_));
 sky130_fd_sc_hd__o21ai_2 _6890_ (.A1(_2215_),
    .A2(_2240_),
    .B1(_2244_),
    .Y(_2245_));
 sky130_fd_sc_hd__nand2b_2 _6891_ (.A_N(_2214_),
    .B(_2245_),
    .Y(_2246_));
 sky130_fd_sc_hd__xor2_1 _6892_ (.A(_2213_),
    .B(_2246_),
    .X(_2247_));
 sky130_fd_sc_hd__xor2_1 _6893_ (.A(_2214_),
    .B(_2245_),
    .X(_2248_));
 sky130_fd_sc_hd__nand2_1 _6894_ (.A(_2241_),
    .B(_2242_),
    .Y(_2249_));
 sky130_fd_sc_hd__and2_1 _6895_ (.A(_2244_),
    .B(_2249_),
    .X(_2250_));
 sky130_fd_sc_hd__xnor2_1 _6896_ (.A(_2235_),
    .B(_2239_),
    .Y(_2251_));
 sky130_fd_sc_hd__xor2_1 _6897_ (.A(_2202_),
    .B(_2238_),
    .X(_2252_));
 sky130_fd_sc_hd__nand2_1 _6898_ (.A(net146),
    .B(net88),
    .Y(_2253_));
 sky130_fd_sc_hd__nand2_1 _6899_ (.A(net137),
    .B(net199),
    .Y(_2255_));
 sky130_fd_sc_hd__or2_1 _6900_ (.A(_2253_),
    .B(_2255_),
    .X(_2256_));
 sky130_fd_sc_hd__o22a_1 _6901_ (.A1(net149),
    .A2(net91),
    .B1(net200),
    .B2(net179),
    .X(_2257_));
 sky130_fd_sc_hd__or2_4 _6902_ (.A(net179),
    .B(net84),
    .X(_2258_));
 sky130_fd_sc_hd__or4_4 _6903_ (.A(_2205_),
    .B(_2216_),
    .C(_2257_),
    .D(_2258_),
    .X(_2259_));
 sky130_fd_sc_hd__o22ai_2 _6904_ (.A1(_2216_),
    .A2(_2257_),
    .B1(_2258_),
    .B2(_2205_),
    .Y(_2260_));
 sky130_fd_sc_hd__nand2_2 _6905_ (.A(_2259_),
    .B(_2260_),
    .Y(_2261_));
 sky130_fd_sc_hd__o21a_1 _6906_ (.A1(net144),
    .A2(net67),
    .B1(_2256_),
    .X(_2262_));
 sky130_fd_sc_hd__o21ba_1 _6907_ (.A1(net67),
    .A2(_2256_),
    .B1_N(_2262_),
    .X(_2263_));
 sky130_fd_sc_hd__o22a_1 _6908_ (.A1(net67),
    .A2(_2256_),
    .B1(_2261_),
    .B2(_2262_),
    .X(_2264_));
 sky130_fd_sc_hd__and2b_1 _6909_ (.A_N(_2264_),
    .B(_2252_),
    .X(_2266_));
 sky130_fd_sc_hd__o21a_1 _6910_ (.A1(net161),
    .A2(net89),
    .B1(_2230_),
    .X(_2267_));
 sky130_fd_sc_hd__nor2_1 _6911_ (.A(_2231_),
    .B(_2267_),
    .Y(_2268_));
 sky130_fd_sc_hd__or3_1 _6912_ (.A(_2231_),
    .B(_2259_),
    .C(_2267_),
    .X(_2269_));
 sky130_fd_sc_hd__xnor2_2 _6913_ (.A(_2259_),
    .B(_2268_),
    .Y(_2270_));
 sky130_fd_sc_hd__xnor2_4 _6914_ (.A(_2226_),
    .B(_2228_),
    .Y(_2271_));
 sky130_fd_sc_hd__nor2_2 _6915_ (.A(net127),
    .B(net110),
    .Y(_2272_));
 sky130_fd_sc_hd__and3_2 _6916_ (.A(net128),
    .B(net76),
    .C(_0611_),
    .X(_2273_));
 sky130_fd_sc_hd__nor2_4 _6917_ (.A(net166),
    .B(net79),
    .Y(_2274_));
 sky130_fd_sc_hd__a21oi_2 _6918_ (.A1(_3475_),
    .A2(net76),
    .B1(_0611_),
    .Y(_2275_));
 sky130_fd_sc_hd__nor2_4 _6919_ (.A(_2273_),
    .B(_2275_),
    .Y(_2277_));
 sky130_fd_sc_hd__a21oi_2 _6920_ (.A1(_2274_),
    .A2(_2277_),
    .B1(_2273_),
    .Y(_2278_));
 sky130_fd_sc_hd__nand2b_1 _6921_ (.A_N(_2278_),
    .B(_2271_),
    .Y(_2279_));
 sky130_fd_sc_hd__nor2_2 _6922_ (.A(net161),
    .B(net84),
    .Y(_2280_));
 sky130_fd_sc_hd__xnor2_2 _6923_ (.A(_2271_),
    .B(_2278_),
    .Y(_2281_));
 sky130_fd_sc_hd__a21bo_1 _6924_ (.A1(_2280_),
    .A2(_2281_),
    .B1_N(_2279_),
    .X(_2282_));
 sky130_fd_sc_hd__xnor2_1 _6925_ (.A(_2270_),
    .B(_2282_),
    .Y(_2283_));
 sky130_fd_sc_hd__and2b_1 _6926_ (.A_N(_2252_),
    .B(_2264_),
    .X(_2284_));
 sky130_fd_sc_hd__or2_1 _6927_ (.A(_2266_),
    .B(_2284_),
    .X(_2285_));
 sky130_fd_sc_hd__nor2_1 _6928_ (.A(_2283_),
    .B(_2285_),
    .Y(_2286_));
 sky130_fd_sc_hd__o21a_1 _6929_ (.A1(_2266_),
    .A2(_2286_),
    .B1(_2251_),
    .X(_2288_));
 sky130_fd_sc_hd__a21bo_2 _6930_ (.A1(_2270_),
    .A2(_2282_),
    .B1_N(_2269_),
    .X(_2289_));
 sky130_fd_sc_hd__nor3_1 _6931_ (.A(_2251_),
    .B(_2266_),
    .C(_2286_),
    .Y(_2290_));
 sky130_fd_sc_hd__or2_2 _6932_ (.A(_2288_),
    .B(_2290_),
    .X(_2291_));
 sky130_fd_sc_hd__and2b_1 _6933_ (.A_N(_2291_),
    .B(_2289_),
    .X(_2292_));
 sky130_fd_sc_hd__o21ai_1 _6934_ (.A1(_2288_),
    .A2(_2292_),
    .B1(_2250_),
    .Y(_2293_));
 sky130_fd_sc_hd__nor2_1 _6935_ (.A(_2248_),
    .B(_2293_),
    .Y(_2294_));
 sky130_fd_sc_hd__and2_1 _6936_ (.A(_2248_),
    .B(_2293_),
    .X(_2295_));
 sky130_fd_sc_hd__or2_2 _6937_ (.A(_2294_),
    .B(_2295_),
    .X(_2296_));
 sky130_fd_sc_hd__inv_2 _6938_ (.A(_2296_),
    .Y(_2297_));
 sky130_fd_sc_hd__xnor2_2 _6939_ (.A(_2289_),
    .B(_2291_),
    .Y(_2299_));
 sky130_fd_sc_hd__nand2_1 _6940_ (.A(_2283_),
    .B(_2285_),
    .Y(_2300_));
 sky130_fd_sc_hd__nand2b_2 _6941_ (.A_N(_2286_),
    .B(_2300_),
    .Y(_2301_));
 sky130_fd_sc_hd__xor2_2 _6942_ (.A(_2261_),
    .B(_2263_),
    .X(_2302_));
 sky130_fd_sc_hd__xor2_1 _6943_ (.A(_2253_),
    .B(_2255_),
    .X(_2303_));
 sky130_fd_sc_hd__nor2_2 _6944_ (.A(net134),
    .B(net84),
    .Y(_2304_));
 sky130_fd_sc_hd__or2_2 _6945_ (.A(net71),
    .B(net134),
    .X(_2305_));
 sky130_fd_sc_hd__or3_1 _6946_ (.A(net134),
    .B(net84),
    .C(_2202_),
    .X(_2306_));
 sky130_fd_sc_hd__or4b_2 _6947_ (.A(net134),
    .B(_0363_),
    .C(_2202_),
    .D_N(_2303_),
    .X(_2307_));
 sky130_fd_sc_hd__o22a_1 _6948_ (.A1(net71),
    .A2(net179),
    .B1(net84),
    .B2(net149),
    .X(_2308_));
 sky130_fd_sc_hd__o21ba_1 _6949_ (.A1(_2205_),
    .A2(_2258_),
    .B1_N(_2308_),
    .X(_2310_));
 sky130_fd_sc_hd__nand2_2 _6950_ (.A(net124),
    .B(net64),
    .Y(_2311_));
 sky130_fd_sc_hd__and4_2 _6951_ (.A(_3496_),
    .B(net124),
    .C(net64),
    .D(net199),
    .X(_2312_));
 sky130_fd_sc_hd__nand2_2 _6952_ (.A(net154),
    .B(net83),
    .Y(_2313_));
 sky130_fd_sc_hd__o22a_1 _6953_ (.A1(net179),
    .A2(net66),
    .B1(net200),
    .B2(net123),
    .X(_2314_));
 sky130_fd_sc_hd__nor2_4 _6954_ (.A(_2312_),
    .B(_2314_),
    .Y(_2315_));
 sky130_fd_sc_hd__and3_1 _6955_ (.A(net154),
    .B(net83),
    .C(_2315_),
    .X(_2316_));
 sky130_fd_sc_hd__o21ai_2 _6956_ (.A1(_2312_),
    .A2(_2316_),
    .B1(_2310_),
    .Y(_2317_));
 sky130_fd_sc_hd__or3_1 _6957_ (.A(_2310_),
    .B(_2312_),
    .C(_2316_),
    .X(_2318_));
 sky130_fd_sc_hd__and2_1 _6958_ (.A(_2317_),
    .B(_2318_),
    .X(_2319_));
 sky130_fd_sc_hd__a31o_1 _6959_ (.A1(_3464_),
    .A2(net146),
    .A3(_2304_),
    .B1(_2303_),
    .X(_2321_));
 sky130_fd_sc_hd__nand2_1 _6960_ (.A(_2307_),
    .B(_2321_),
    .Y(_2322_));
 sky130_fd_sc_hd__inv_2 _6961_ (.A(_2322_),
    .Y(_2323_));
 sky130_fd_sc_hd__nand2_1 _6962_ (.A(_2319_),
    .B(_2323_),
    .Y(_2324_));
 sky130_fd_sc_hd__a21o_2 _6963_ (.A1(_2307_),
    .A2(_2324_),
    .B1(_2302_),
    .X(_2325_));
 sky130_fd_sc_hd__xnor2_2 _6964_ (.A(_2280_),
    .B(_2281_),
    .Y(_2326_));
 sky130_fd_sc_hd__nor2_2 _6965_ (.A(_2317_),
    .B(_2326_),
    .Y(_2327_));
 sky130_fd_sc_hd__and2_1 _6966_ (.A(_2317_),
    .B(_2326_),
    .X(_2328_));
 sky130_fd_sc_hd__nor2_4 _6967_ (.A(_2327_),
    .B(_2328_),
    .Y(_2329_));
 sky130_fd_sc_hd__xnor2_4 _6968_ (.A(_2274_),
    .B(_2277_),
    .Y(_2330_));
 sky130_fd_sc_hd__or2_4 _6969_ (.A(_3476_),
    .B(net107),
    .X(_2332_));
 sky130_fd_sc_hd__xor2_1 _6970_ (.A(_0596_),
    .B(_2272_),
    .X(_2333_));
 sky130_fd_sc_hd__or3b_1 _6971_ (.A(net166),
    .B(net74),
    .C_N(_2333_),
    .X(_2334_));
 sky130_fd_sc_hd__a21bo_4 _6972_ (.A1(_0596_),
    .A2(_2272_),
    .B1_N(_2334_),
    .X(_2335_));
 sky130_fd_sc_hd__nand2b_1 _6973_ (.A_N(_2330_),
    .B(_2335_),
    .Y(_2336_));
 sky130_fd_sc_hd__nor2_1 _6974_ (.A(net161),
    .B(net82),
    .Y(_2337_));
 sky130_fd_sc_hd__xor2_4 _6975_ (.A(_2330_),
    .B(_2335_),
    .X(_2338_));
 sky130_fd_sc_hd__o31ai_4 _6976_ (.A1(net161),
    .A2(net82),
    .A3(_2338_),
    .B1(_2336_),
    .Y(_2339_));
 sky130_fd_sc_hd__xor2_4 _6977_ (.A(_2329_),
    .B(_2339_),
    .X(_2340_));
 sky130_fd_sc_hd__nand3_1 _6978_ (.A(_2302_),
    .B(_2307_),
    .C(_2324_),
    .Y(_2341_));
 sky130_fd_sc_hd__and2_1 _6979_ (.A(_2325_),
    .B(_2341_),
    .X(_2343_));
 sky130_fd_sc_hd__nand2_4 _6980_ (.A(_2340_),
    .B(_2343_),
    .Y(_2344_));
 sky130_fd_sc_hd__a21oi_4 _6981_ (.A1(_2325_),
    .A2(_2344_),
    .B1(_2301_),
    .Y(_2345_));
 sky130_fd_sc_hd__a21o_2 _6982_ (.A1(_2329_),
    .A2(_2339_),
    .B1(_2327_),
    .X(_2346_));
 sky130_fd_sc_hd__and3_1 _6983_ (.A(_2301_),
    .B(_2325_),
    .C(_2344_),
    .X(_2347_));
 sky130_fd_sc_hd__or2_2 _6984_ (.A(_2345_),
    .B(_2347_),
    .X(_2348_));
 sky130_fd_sc_hd__and2b_1 _6985_ (.A_N(_2348_),
    .B(_2346_),
    .X(_2349_));
 sky130_fd_sc_hd__o21ai_4 _6986_ (.A1(_2345_),
    .A2(_2349_),
    .B1(_2299_),
    .Y(_2350_));
 sky130_fd_sc_hd__or3_1 _6987_ (.A(_2250_),
    .B(_2288_),
    .C(_2292_),
    .X(_2351_));
 sky130_fd_sc_hd__and2_2 _6988_ (.A(_2293_),
    .B(_2351_),
    .X(_2352_));
 sky130_fd_sc_hd__and2b_1 _6989_ (.A_N(_2350_),
    .B(_2352_),
    .X(_2354_));
 sky130_fd_sc_hd__xor2_4 _6990_ (.A(_2350_),
    .B(_2352_),
    .X(_2355_));
 sky130_fd_sc_hd__or3_1 _6991_ (.A(_2299_),
    .B(_2345_),
    .C(_2349_),
    .X(_2356_));
 sky130_fd_sc_hd__nand2_1 _6992_ (.A(_2350_),
    .B(_2356_),
    .Y(_2357_));
 sky130_fd_sc_hd__xnor2_2 _6993_ (.A(_2346_),
    .B(_2348_),
    .Y(_2358_));
 sky130_fd_sc_hd__or2_2 _6994_ (.A(_2340_),
    .B(_2343_),
    .X(_2359_));
 sky130_fd_sc_hd__nand2_4 _6995_ (.A(_2344_),
    .B(_2359_),
    .Y(_2360_));
 sky130_fd_sc_hd__xnor2_1 _6996_ (.A(_2319_),
    .B(_2323_),
    .Y(_2361_));
 sky130_fd_sc_hd__o21ai_1 _6997_ (.A1(net144),
    .A2(net84),
    .B1(_2305_),
    .Y(_2362_));
 sky130_fd_sc_hd__and2_1 _6998_ (.A(_2306_),
    .B(_2362_),
    .X(_2363_));
 sky130_fd_sc_hd__nand2_4 _6999_ (.A(net146),
    .B(net83),
    .Y(_2365_));
 sky130_fd_sc_hd__o22a_1 _7000_ (.A1(net134),
    .A2(net66),
    .B1(net200),
    .B2(net176),
    .X(_2366_));
 sky130_fd_sc_hd__nor2_4 _7001_ (.A(net176),
    .B(net66),
    .Y(_2367_));
 sky130_fd_sc_hd__nand2_2 _7002_ (.A(net137),
    .B(_2367_),
    .Y(_2368_));
 sky130_fd_sc_hd__a21o_2 _7003_ (.A1(net137),
    .A2(_2367_),
    .B1(_2366_),
    .X(_2369_));
 sky130_fd_sc_hd__nor2_1 _7004_ (.A(_2365_),
    .B(_2369_),
    .Y(_2370_));
 sky130_fd_sc_hd__nand2_2 _7005_ (.A(_2363_),
    .B(_2370_),
    .Y(_2371_));
 sky130_fd_sc_hd__xnor2_4 _7006_ (.A(_2313_),
    .B(_2315_),
    .Y(_2372_));
 sky130_fd_sc_hd__and3_1 _7007_ (.A(net137),
    .B(_2367_),
    .C(_2372_),
    .X(_2373_));
 sky130_fd_sc_hd__xnor2_4 _7008_ (.A(_2368_),
    .B(_2372_),
    .Y(_2374_));
 sky130_fd_sc_hd__nand2_2 _7009_ (.A(net181),
    .B(net88),
    .Y(_2376_));
 sky130_fd_sc_hd__or3_1 _7010_ (.A(net71),
    .B(net122),
    .C(_2376_),
    .X(_2377_));
 sky130_fd_sc_hd__o21ai_2 _7011_ (.A1(net71),
    .A2(net123),
    .B1(_2376_),
    .Y(_2378_));
 sky130_fd_sc_hd__nor2_1 _7012_ (.A(net149),
    .B(net79),
    .Y(_2379_));
 sky130_fd_sc_hd__and3_1 _7013_ (.A(_2377_),
    .B(_2378_),
    .C(_2379_),
    .X(_2380_));
 sky130_fd_sc_hd__a21bo_4 _7014_ (.A1(_2378_),
    .A2(_2379_),
    .B1_N(_2377_),
    .X(_2381_));
 sky130_fd_sc_hd__xnor2_4 _7015_ (.A(_2374_),
    .B(_2381_),
    .Y(_2382_));
 sky130_fd_sc_hd__or2_1 _7016_ (.A(_2363_),
    .B(_2370_),
    .X(_2383_));
 sky130_fd_sc_hd__nand2_2 _7017_ (.A(_2371_),
    .B(_2383_),
    .Y(_2384_));
 sky130_fd_sc_hd__or2_1 _7018_ (.A(_2382_),
    .B(_2384_),
    .X(_2385_));
 sky130_fd_sc_hd__a21o_1 _7019_ (.A1(_2371_),
    .A2(_2385_),
    .B1(_2361_),
    .X(_2387_));
 sky130_fd_sc_hd__a21o_1 _7020_ (.A1(_2374_),
    .A2(_2381_),
    .B1(_2373_),
    .X(_2388_));
 sky130_fd_sc_hd__xnor2_2 _7021_ (.A(_2337_),
    .B(_2338_),
    .Y(_2389_));
 sky130_fd_sc_hd__xnor2_1 _7022_ (.A(_2388_),
    .B(_2389_),
    .Y(_2390_));
 sky130_fd_sc_hd__a21o_1 _7023_ (.A1(net163),
    .A2(net76),
    .B1(_2333_),
    .X(_2391_));
 sky130_fd_sc_hd__and2_2 _7024_ (.A(_2334_),
    .B(_2391_),
    .X(_2392_));
 sky130_fd_sc_hd__nor2_1 _7025_ (.A(net127),
    .B(net105),
    .Y(_2393_));
 sky130_fd_sc_hd__xor2_2 _7026_ (.A(_0597_),
    .B(_2332_),
    .X(_2394_));
 sky130_fd_sc_hd__or3_2 _7027_ (.A(net166),
    .B(net110),
    .C(_2394_),
    .X(_2395_));
 sky130_fd_sc_hd__o31a_2 _7028_ (.A1(net211),
    .A2(net105),
    .A3(_2332_),
    .B1(_2395_),
    .X(_2396_));
 sky130_fd_sc_hd__and2b_1 _7029_ (.A_N(_2396_),
    .B(_2392_),
    .X(_2398_));
 sky130_fd_sc_hd__nor2_2 _7030_ (.A(net161),
    .B(net79),
    .Y(_2399_));
 sky130_fd_sc_hd__xnor2_2 _7031_ (.A(_2392_),
    .B(_2396_),
    .Y(_2400_));
 sky130_fd_sc_hd__a21oi_1 _7032_ (.A1(_2399_),
    .A2(_2400_),
    .B1(_2398_),
    .Y(_2401_));
 sky130_fd_sc_hd__or2_1 _7033_ (.A(_2390_),
    .B(_2401_),
    .X(_2402_));
 sky130_fd_sc_hd__nand2_1 _7034_ (.A(_2390_),
    .B(_2401_),
    .Y(_2403_));
 sky130_fd_sc_hd__nand2_1 _7035_ (.A(_2402_),
    .B(_2403_),
    .Y(_2404_));
 sky130_fd_sc_hd__nand3_1 _7036_ (.A(_2361_),
    .B(_2371_),
    .C(_2385_),
    .Y(_2405_));
 sky130_fd_sc_hd__nand2_1 _7037_ (.A(_2387_),
    .B(_2405_),
    .Y(_2406_));
 sky130_fd_sc_hd__or2_1 _7038_ (.A(_2404_),
    .B(_2406_),
    .X(_2407_));
 sky130_fd_sc_hd__and2_2 _7039_ (.A(_2387_),
    .B(_2407_),
    .X(_2409_));
 sky130_fd_sc_hd__a21bo_4 _7040_ (.A1(_2388_),
    .A2(_2389_),
    .B1_N(_2402_),
    .X(_2410_));
 sky130_fd_sc_hd__xnor2_4 _7041_ (.A(_2360_),
    .B(_2409_),
    .Y(_2411_));
 sky130_fd_sc_hd__and2b_1 _7042_ (.A_N(_2411_),
    .B(_2410_),
    .X(_2412_));
 sky130_fd_sc_hd__o21ba_1 _7043_ (.A1(_2360_),
    .A2(_2409_),
    .B1_N(_2412_),
    .X(_2413_));
 sky130_fd_sc_hd__nand2b_1 _7044_ (.A_N(_2413_),
    .B(_2358_),
    .Y(_2414_));
 sky130_fd_sc_hd__xnor2_1 _7045_ (.A(_2358_),
    .B(_2413_),
    .Y(_2415_));
 sky130_fd_sc_hd__or3b_2 _7046_ (.A(net138),
    .B(net200),
    .C_N(_2415_),
    .X(_2416_));
 sky130_fd_sc_hd__a21oi_2 _7047_ (.A1(_2414_),
    .A2(_2416_),
    .B1(_2357_),
    .Y(_2417_));
 sky130_fd_sc_hd__and3_1 _7048_ (.A(_2357_),
    .B(_2414_),
    .C(_2416_),
    .X(_2418_));
 sky130_fd_sc_hd__nor2_1 _7049_ (.A(_2417_),
    .B(_2418_),
    .Y(_2420_));
 sky130_fd_sc_hd__a21o_1 _7050_ (.A1(_3498_),
    .A2(net199),
    .B1(_2415_),
    .X(_2421_));
 sky130_fd_sc_hd__nand2_1 _7051_ (.A(_2416_),
    .B(_2421_),
    .Y(_2422_));
 sky130_fd_sc_hd__xor2_4 _7052_ (.A(_2410_),
    .B(_2411_),
    .X(_2423_));
 sky130_fd_sc_hd__nand2_1 _7053_ (.A(_2404_),
    .B(_2406_),
    .Y(_2424_));
 sky130_fd_sc_hd__and2_2 _7054_ (.A(_2407_),
    .B(_2424_),
    .X(_2425_));
 sky130_fd_sc_hd__xnor2_4 _7055_ (.A(_2382_),
    .B(_2384_),
    .Y(_2426_));
 sky130_fd_sc_hd__xor2_4 _7056_ (.A(_2365_),
    .B(_2369_),
    .X(_2427_));
 sky130_fd_sc_hd__nor2_1 _7057_ (.A(net144),
    .B(net79),
    .Y(_2428_));
 sky130_fd_sc_hd__nand2_2 _7058_ (.A(_3702_),
    .B(net88),
    .Y(_2429_));
 sky130_fd_sc_hd__o22a_1 _7059_ (.A1(net71),
    .A2(net174),
    .B1(net91),
    .B2(net134),
    .X(_2431_));
 sky130_fd_sc_hd__o21ba_1 _7060_ (.A1(_2305_),
    .A2(_2429_),
    .B1_N(_2431_),
    .X(_2432_));
 sky130_fd_sc_hd__and2_2 _7061_ (.A(_2428_),
    .B(_2432_),
    .X(_2433_));
 sky130_fd_sc_hd__nand2_4 _7062_ (.A(_2427_),
    .B(_2433_),
    .Y(_2434_));
 sky130_fd_sc_hd__or2_2 _7063_ (.A(_2427_),
    .B(_2433_),
    .X(_2435_));
 sky130_fd_sc_hd__nand2_4 _7064_ (.A(_2434_),
    .B(_2435_),
    .Y(_2436_));
 sky130_fd_sc_hd__a2111oi_4 _7065_ (.A1(net168),
    .A2(_0359_),
    .B1(_0362_),
    .C1(net123),
    .D1(net172),
    .Y(_2437_));
 sky130_fd_sc_hd__nor2_1 _7066_ (.A(_2258_),
    .B(_2311_),
    .Y(_2438_));
 sky130_fd_sc_hd__xor2_4 _7067_ (.A(_2258_),
    .B(_2311_),
    .X(_2439_));
 sky130_fd_sc_hd__nand2_2 _7068_ (.A(net154),
    .B(net76),
    .Y(_2440_));
 sky130_fd_sc_hd__a31o_4 _7069_ (.A1(net154),
    .A2(net76),
    .A3(_2439_),
    .B1(_2438_),
    .X(_2442_));
 sky130_fd_sc_hd__a21oi_1 _7070_ (.A1(_2377_),
    .A2(_2378_),
    .B1(_2379_),
    .Y(_2443_));
 sky130_fd_sc_hd__or2_1 _7071_ (.A(_2380_),
    .B(_2443_),
    .X(_2444_));
 sky130_fd_sc_hd__or3_1 _7072_ (.A(_2305_),
    .B(_2429_),
    .C(_2444_),
    .X(_2445_));
 sky130_fd_sc_hd__o21ai_1 _7073_ (.A1(_2305_),
    .A2(_2429_),
    .B1(_2444_),
    .Y(_2446_));
 sky130_fd_sc_hd__and2_2 _7074_ (.A(_2445_),
    .B(_2446_),
    .X(_2447_));
 sky130_fd_sc_hd__nand2_1 _7075_ (.A(_2442_),
    .B(_2447_),
    .Y(_2448_));
 sky130_fd_sc_hd__xnor2_4 _7076_ (.A(_2442_),
    .B(_2447_),
    .Y(_2449_));
 sky130_fd_sc_hd__or2_2 _7077_ (.A(_2436_),
    .B(_2449_),
    .X(_2450_));
 sky130_fd_sc_hd__a21oi_4 _7078_ (.A1(_2434_),
    .A2(_2450_),
    .B1(_2426_),
    .Y(_2451_));
 sky130_fd_sc_hd__xnor2_2 _7079_ (.A(_2399_),
    .B(_2400_),
    .Y(_2453_));
 sky130_fd_sc_hd__a21oi_1 _7080_ (.A1(_2445_),
    .A2(_2448_),
    .B1(_2453_),
    .Y(_2454_));
 sky130_fd_sc_hd__and3_1 _7081_ (.A(_2445_),
    .B(_2448_),
    .C(_2453_),
    .X(_2455_));
 sky130_fd_sc_hd__or2_4 _7082_ (.A(_2454_),
    .B(_2455_),
    .X(_2456_));
 sky130_fd_sc_hd__o21ai_2 _7083_ (.A1(net166),
    .A2(net110),
    .B1(_2394_),
    .Y(_2457_));
 sky130_fd_sc_hd__nand2_4 _7084_ (.A(_2395_),
    .B(_2457_),
    .Y(_2458_));
 sky130_fd_sc_hd__nand2_1 _7085_ (.A(net162),
    .B(_0587_),
    .Y(_2459_));
 sky130_fd_sc_hd__or2_4 _7086_ (.A(_2332_),
    .B(_2459_),
    .X(_2460_));
 sky130_fd_sc_hd__xnor2_4 _7087_ (.A(_2458_),
    .B(_2460_),
    .Y(_2461_));
 sky130_fd_sc_hd__nor2_2 _7088_ (.A(net160),
    .B(net75),
    .Y(_2462_));
 sky130_fd_sc_hd__o32a_4 _7089_ (.A1(net161),
    .A2(net75),
    .A3(_2461_),
    .B1(_2460_),
    .B2(_2458_),
    .X(_2464_));
 sky130_fd_sc_hd__xnor2_4 _7090_ (.A(_2456_),
    .B(_2464_),
    .Y(_2465_));
 sky130_fd_sc_hd__and3_1 _7091_ (.A(_2426_),
    .B(_2434_),
    .C(_2450_),
    .X(_2466_));
 sky130_fd_sc_hd__nor2_2 _7092_ (.A(_2451_),
    .B(_2466_),
    .Y(_2467_));
 sky130_fd_sc_hd__and2b_2 _7093_ (.A_N(_2465_),
    .B(_2467_),
    .X(_2468_));
 sky130_fd_sc_hd__nor2_4 _7094_ (.A(_2451_),
    .B(_2468_),
    .Y(_2469_));
 sky130_fd_sc_hd__nand2b_1 _7095_ (.A_N(_2469_),
    .B(_2425_),
    .Y(_2470_));
 sky130_fd_sc_hd__o21ba_4 _7096_ (.A1(_2456_),
    .A2(_2464_),
    .B1_N(_2454_),
    .X(_2471_));
 sky130_fd_sc_hd__xnor2_4 _7097_ (.A(_2425_),
    .B(_2469_),
    .Y(_2472_));
 sky130_fd_sc_hd__nand2b_1 _7098_ (.A_N(_2471_),
    .B(_2472_),
    .Y(_2473_));
 sky130_fd_sc_hd__and2_2 _7099_ (.A(_2470_),
    .B(_2473_),
    .X(_2475_));
 sky130_fd_sc_hd__or2_1 _7100_ (.A(_2423_),
    .B(_2475_),
    .X(_2476_));
 sky130_fd_sc_hd__or2_4 _7101_ (.A(net71),
    .B(net138),
    .X(_2477_));
 sky130_fd_sc_hd__xnor2_4 _7102_ (.A(_2423_),
    .B(_2475_),
    .Y(_2478_));
 sky130_fd_sc_hd__o21ai_2 _7103_ (.A1(_2477_),
    .A2(_2478_),
    .B1(_2476_),
    .Y(_2479_));
 sky130_fd_sc_hd__nand2b_1 _7104_ (.A_N(_2422_),
    .B(_2479_),
    .Y(_2480_));
 sky130_fd_sc_hd__nand2b_1 _7105_ (.A_N(_2479_),
    .B(_2422_),
    .Y(_2481_));
 sky130_fd_sc_hd__nand2_1 _7106_ (.A(_2480_),
    .B(_2481_),
    .Y(_2482_));
 sky130_fd_sc_hd__xnor2_4 _7107_ (.A(_2477_),
    .B(_2478_),
    .Y(_2483_));
 sky130_fd_sc_hd__xnor2_4 _7108_ (.A(_2471_),
    .B(_2472_),
    .Y(_2484_));
 sky130_fd_sc_hd__o21a_1 _7109_ (.A1(_2451_),
    .A2(_2466_),
    .B1(_2465_),
    .X(_2486_));
 sky130_fd_sc_hd__xnor2_4 _7110_ (.A(_2465_),
    .B(_2467_),
    .Y(_2487_));
 sky130_fd_sc_hd__xnor2_4 _7111_ (.A(_2436_),
    .B(_2449_),
    .Y(_2488_));
 sky130_fd_sc_hd__xnor2_1 _7112_ (.A(_2428_),
    .B(_2432_),
    .Y(_2489_));
 sky130_fd_sc_hd__or2_1 _7113_ (.A(net175),
    .B(net84),
    .X(_2490_));
 sky130_fd_sc_hd__and3_4 _7114_ (.A(_3702_),
    .B(net64),
    .C(_2304_),
    .X(_2491_));
 sky130_fd_sc_hd__o21ba_4 _7115_ (.A1(_2304_),
    .A2(_2367_),
    .B1_N(_2491_),
    .X(_2492_));
 sky130_fd_sc_hd__nor2_4 _7116_ (.A(net143),
    .B(net75),
    .Y(_2493_));
 sky130_fd_sc_hd__nand2_1 _7117_ (.A(_2492_),
    .B(_2493_),
    .Y(_2494_));
 sky130_fd_sc_hd__or2_1 _7118_ (.A(_2489_),
    .B(_2494_),
    .X(_2495_));
 sky130_fd_sc_hd__nand2_1 _7119_ (.A(_2489_),
    .B(_2494_),
    .Y(_2497_));
 sky130_fd_sc_hd__and2_1 _7120_ (.A(_2495_),
    .B(_2497_),
    .X(_2498_));
 sky130_fd_sc_hd__a2111o_4 _7121_ (.A1(net167),
    .A2(_3451_),
    .B1(net123),
    .C1(_0371_),
    .D1(net172),
    .X(_2499_));
 sky130_fd_sc_hd__or2_2 _7122_ (.A(_2376_),
    .B(_2499_),
    .X(_2500_));
 sky130_fd_sc_hd__nand2_4 _7123_ (.A(net153),
    .B(net113),
    .Y(_2501_));
 sky130_fd_sc_hd__o22a_2 _7124_ (.A1(net122),
    .A2(net91),
    .B1(net82),
    .B2(net177),
    .X(_2502_));
 sky130_fd_sc_hd__o21ba_2 _7125_ (.A1(_2376_),
    .A2(_2499_),
    .B1_N(_2502_),
    .X(_2503_));
 sky130_fd_sc_hd__o21ai_4 _7126_ (.A1(_2501_),
    .A2(_2502_),
    .B1(_2500_),
    .Y(_2504_));
 sky130_fd_sc_hd__xnor2_4 _7127_ (.A(_2439_),
    .B(_2440_),
    .Y(_2505_));
 sky130_fd_sc_hd__xnor2_4 _7128_ (.A(_2491_),
    .B(_2505_),
    .Y(_2506_));
 sky130_fd_sc_hd__and2b_1 _7129_ (.A_N(_2506_),
    .B(_2504_),
    .X(_2508_));
 sky130_fd_sc_hd__xnor2_2 _7130_ (.A(_2504_),
    .B(_2506_),
    .Y(_2509_));
 sky130_fd_sc_hd__nand2_2 _7131_ (.A(_2498_),
    .B(_2509_),
    .Y(_2510_));
 sky130_fd_sc_hd__nand2_2 _7132_ (.A(_2495_),
    .B(_2510_),
    .Y(_2511_));
 sky130_fd_sc_hd__and2b_1 _7133_ (.A_N(_2488_),
    .B(_2511_),
    .X(_2512_));
 sky130_fd_sc_hd__and3_1 _7134_ (.A(_2488_),
    .B(_2495_),
    .C(_2510_),
    .X(_2513_));
 sky130_fd_sc_hd__xnor2_4 _7135_ (.A(_2488_),
    .B(_2511_),
    .Y(_2514_));
 sky130_fd_sc_hd__nor2_2 _7136_ (.A(net164),
    .B(net106),
    .Y(_2515_));
 sky130_fd_sc_hd__o21a_2 _7137_ (.A1(_2393_),
    .A2(_2515_),
    .B1(_2460_),
    .X(_2516_));
 sky130_fd_sc_hd__nor2_2 _7138_ (.A(net160),
    .B(net110),
    .Y(_2517_));
 sky130_fd_sc_hd__and2_2 _7139_ (.A(_2516_),
    .B(_2517_),
    .X(_2519_));
 sky130_fd_sc_hd__a21o_4 _7140_ (.A1(_2491_),
    .A2(_2505_),
    .B1(_2508_),
    .X(_2520_));
 sky130_fd_sc_hd__xnor2_4 _7141_ (.A(_2461_),
    .B(_2462_),
    .Y(_2521_));
 sky130_fd_sc_hd__xor2_4 _7142_ (.A(_2520_),
    .B(_2521_),
    .X(_2522_));
 sky130_fd_sc_hd__xnor2_4 _7143_ (.A(_2519_),
    .B(_2522_),
    .Y(_2523_));
 sky130_fd_sc_hd__o21ba_4 _7144_ (.A1(_2513_),
    .A2(_2523_),
    .B1_N(_2512_),
    .X(_2524_));
 sky130_fd_sc_hd__a32o_4 _7145_ (.A1(_2516_),
    .A2(_2517_),
    .A3(_2522_),
    .B1(_2521_),
    .B2(_2520_),
    .X(_2525_));
 sky130_fd_sc_hd__xnor2_4 _7146_ (.A(_2487_),
    .B(_2524_),
    .Y(_2526_));
 sky130_fd_sc_hd__nand2_1 _7147_ (.A(_2525_),
    .B(_2526_),
    .Y(_2527_));
 sky130_fd_sc_hd__o31a_4 _7148_ (.A1(_2468_),
    .A2(_2486_),
    .A3(_2524_),
    .B1(_2527_),
    .X(_2528_));
 sky130_fd_sc_hd__nand2b_1 _7149_ (.A_N(_2528_),
    .B(_2484_),
    .Y(_2530_));
 sky130_fd_sc_hd__nor2_1 _7150_ (.A(_3499_),
    .B(net66),
    .Y(_2531_));
 sky130_fd_sc_hd__xor2_4 _7151_ (.A(_2484_),
    .B(_2528_),
    .X(_2532_));
 sky130_fd_sc_hd__o31a_2 _7152_ (.A1(_3499_),
    .A2(net66),
    .A3(_2532_),
    .B1(_2530_),
    .X(_2533_));
 sky130_fd_sc_hd__nor2_4 _7153_ (.A(_2483_),
    .B(_2533_),
    .Y(_2534_));
 sky130_fd_sc_hd__and2_1 _7154_ (.A(_2483_),
    .B(_2533_),
    .X(_2535_));
 sky130_fd_sc_hd__nor2_4 _7155_ (.A(_2534_),
    .B(_2535_),
    .Y(_2536_));
 sky130_fd_sc_hd__xnor2_2 _7156_ (.A(_2531_),
    .B(_2532_),
    .Y(_2537_));
 sky130_fd_sc_hd__xnor2_4 _7157_ (.A(_2525_),
    .B(_2526_),
    .Y(_2538_));
 sky130_fd_sc_hd__xnor2_4 _7158_ (.A(_2514_),
    .B(_2523_),
    .Y(_2539_));
 sky130_fd_sc_hd__or2_2 _7159_ (.A(_2498_),
    .B(_2509_),
    .X(_2541_));
 sky130_fd_sc_hd__nand2_4 _7160_ (.A(_2510_),
    .B(_2541_),
    .Y(_2542_));
 sky130_fd_sc_hd__xnor2_4 _7161_ (.A(_2492_),
    .B(_2493_),
    .Y(_2543_));
 sky130_fd_sc_hd__nand2_1 _7162_ (.A(net136),
    .B(net83),
    .Y(_2544_));
 sky130_fd_sc_hd__and4_4 _7163_ (.A(net136),
    .B(_3702_),
    .C(net88),
    .D(net83),
    .X(_2545_));
 sky130_fd_sc_hd__a21o_1 _7164_ (.A1(_2429_),
    .A2(_2544_),
    .B1(_2545_),
    .X(_2546_));
 sky130_fd_sc_hd__nand2_2 _7165_ (.A(net145),
    .B(net113),
    .Y(_2547_));
 sky130_fd_sc_hd__or2_4 _7166_ (.A(_2546_),
    .B(_2547_),
    .X(_2548_));
 sky130_fd_sc_hd__xnor2_4 _7167_ (.A(_2501_),
    .B(_2503_),
    .Y(_2549_));
 sky130_fd_sc_hd__nand2_1 _7168_ (.A(_2545_),
    .B(_2549_),
    .Y(_2550_));
 sky130_fd_sc_hd__xnor2_4 _7169_ (.A(_2545_),
    .B(_2549_),
    .Y(_2552_));
 sky130_fd_sc_hd__and3_2 _7170_ (.A(net170),
    .B(_1990_),
    .C(net181),
    .X(_2553_));
 sky130_fd_sc_hd__and2_1 _7171_ (.A(_2437_),
    .B(_2553_),
    .X(_2554_));
 sky130_fd_sc_hd__or2_4 _7172_ (.A(net147),
    .B(net106),
    .X(_2555_));
 sky130_fd_sc_hd__xor2_4 _7173_ (.A(_2437_),
    .B(_2553_),
    .X(_2556_));
 sky130_fd_sc_hd__a31o_4 _7174_ (.A1(net153),
    .A2(net73),
    .A3(_2556_),
    .B1(_2554_),
    .X(_2557_));
 sky130_fd_sc_hd__nand2b_1 _7175_ (.A_N(_2552_),
    .B(_2557_),
    .Y(_2558_));
 sky130_fd_sc_hd__xor2_4 _7176_ (.A(_2552_),
    .B(_2557_),
    .X(_2559_));
 sky130_fd_sc_hd__xor2_4 _7177_ (.A(_2543_),
    .B(_2548_),
    .X(_2560_));
 sky130_fd_sc_hd__nand2b_2 _7178_ (.A_N(_2559_),
    .B(_2560_),
    .Y(_2561_));
 sky130_fd_sc_hd__o21ai_4 _7179_ (.A1(_2543_),
    .A2(_2548_),
    .B1(_2561_),
    .Y(_2563_));
 sky130_fd_sc_hd__and2b_1 _7180_ (.A_N(_2542_),
    .B(_2563_),
    .X(_2564_));
 sky130_fd_sc_hd__xor2_4 _7181_ (.A(_2542_),
    .B(_2563_),
    .X(_2565_));
 sky130_fd_sc_hd__xnor2_1 _7182_ (.A(_2516_),
    .B(_2517_),
    .Y(_2566_));
 sky130_fd_sc_hd__a21oi_1 _7183_ (.A1(_2550_),
    .A2(_2558_),
    .B1(_2566_),
    .Y(_2567_));
 sky130_fd_sc_hd__and3_1 _7184_ (.A(_2550_),
    .B(_2558_),
    .C(_2566_),
    .X(_2568_));
 sky130_fd_sc_hd__or2_4 _7185_ (.A(_2567_),
    .B(_2568_),
    .X(_2569_));
 sky130_fd_sc_hd__nor2_4 _7186_ (.A(net160),
    .B(net104),
    .Y(_2570_));
 sky130_fd_sc_hd__nand2_4 _7187_ (.A(_2515_),
    .B(_2570_),
    .Y(_2571_));
 sky130_fd_sc_hd__xnor2_4 _7188_ (.A(_2569_),
    .B(_2571_),
    .Y(_2572_));
 sky130_fd_sc_hd__o21bai_4 _7189_ (.A1(_2565_),
    .A2(_2572_),
    .B1_N(_2564_),
    .Y(_2574_));
 sky130_fd_sc_hd__xnor2_4 _7190_ (.A(_2539_),
    .B(_2574_),
    .Y(_2575_));
 sky130_fd_sc_hd__o21ba_4 _7191_ (.A1(_2569_),
    .A2(_2571_),
    .B1_N(_2567_),
    .X(_2576_));
 sky130_fd_sc_hd__nor2_1 _7192_ (.A(_2575_),
    .B(_2576_),
    .Y(_2577_));
 sky130_fd_sc_hd__a21oi_4 _7193_ (.A1(_2539_),
    .A2(_2574_),
    .B1(_2577_),
    .Y(_2578_));
 sky130_fd_sc_hd__xor2_2 _7194_ (.A(_2538_),
    .B(_2578_),
    .X(_2579_));
 sky130_fd_sc_hd__and3_2 _7195_ (.A(net140),
    .B(net88),
    .C(_2579_),
    .X(_2580_));
 sky130_fd_sc_hd__o21ba_1 _7196_ (.A1(_2538_),
    .A2(_2578_),
    .B1_N(_2580_),
    .X(_2581_));
 sky130_fd_sc_hd__nand2b_4 _7197_ (.A_N(_2581_),
    .B(_2537_),
    .Y(_2582_));
 sky130_fd_sc_hd__nand2b_1 _7198_ (.A_N(_2537_),
    .B(_2581_),
    .Y(_2583_));
 sky130_fd_sc_hd__nand2_4 _7199_ (.A(_2582_),
    .B(_2583_),
    .Y(_2585_));
 sky130_fd_sc_hd__a21oi_2 _7200_ (.A1(net140),
    .A2(net88),
    .B1(_2579_),
    .Y(_2586_));
 sky130_fd_sc_hd__nor2_4 _7201_ (.A(_2580_),
    .B(_2586_),
    .Y(_2587_));
 sky130_fd_sc_hd__xnor2_4 _7202_ (.A(_2575_),
    .B(_2576_),
    .Y(_2588_));
 sky130_fd_sc_hd__xnor2_4 _7203_ (.A(_2565_),
    .B(_2572_),
    .Y(_2589_));
 sky130_fd_sc_hd__xnor2_4 _7204_ (.A(_2559_),
    .B(_2560_),
    .Y(_2590_));
 sky130_fd_sc_hd__xnor2_2 _7205_ (.A(_2546_),
    .B(_2547_),
    .Y(_2591_));
 sky130_fd_sc_hd__nand2_1 _7206_ (.A(net136),
    .B(net80),
    .Y(_2592_));
 sky130_fd_sc_hd__nor4_4 _7207_ (.A(net135),
    .B(net175),
    .C(net84),
    .D(net79),
    .Y(_2593_));
 sky130_fd_sc_hd__a21o_2 _7208_ (.A1(_2490_),
    .A2(_2592_),
    .B1(_2593_),
    .X(_2594_));
 sky130_fd_sc_hd__nor2_2 _7209_ (.A(net142),
    .B(net106),
    .Y(_2596_));
 sky130_fd_sc_hd__or3_2 _7210_ (.A(net142),
    .B(net106),
    .C(_2594_),
    .X(_2597_));
 sky130_fd_sc_hd__xnor2_4 _7211_ (.A(_2555_),
    .B(_2556_),
    .Y(_2598_));
 sky130_fd_sc_hd__xnor2_2 _7212_ (.A(_2593_),
    .B(_2598_),
    .Y(_2599_));
 sky130_fd_sc_hd__and3_4 _7213_ (.A(net170),
    .B(net181),
    .C(_0496_),
    .X(_2600_));
 sky130_fd_sc_hd__or3_1 _7214_ (.A(net177),
    .B(net75),
    .C(_2499_),
    .X(_2601_));
 sky130_fd_sc_hd__nor2_4 _7215_ (.A(net147),
    .B(net104),
    .Y(_2602_));
 sky130_fd_sc_hd__xnor2_4 _7216_ (.A(_2499_),
    .B(_2600_),
    .Y(_2603_));
 sky130_fd_sc_hd__a21bo_1 _7217_ (.A1(_2602_),
    .A2(_2603_),
    .B1_N(_2601_),
    .X(_2604_));
 sky130_fd_sc_hd__and2b_1 _7218_ (.A_N(_2599_),
    .B(_2604_),
    .X(_2605_));
 sky130_fd_sc_hd__xor2_1 _7219_ (.A(_2599_),
    .B(_2604_),
    .X(_2607_));
 sky130_fd_sc_hd__xnor2_1 _7220_ (.A(_2591_),
    .B(_2597_),
    .Y(_2608_));
 sky130_fd_sc_hd__nor2_1 _7221_ (.A(_2607_),
    .B(_2608_),
    .Y(_2609_));
 sky130_fd_sc_hd__o21ba_2 _7222_ (.A1(_2591_),
    .A2(_2597_),
    .B1_N(_2609_),
    .X(_2610_));
 sky130_fd_sc_hd__nand2b_1 _7223_ (.A_N(_2610_),
    .B(_2590_),
    .Y(_2611_));
 sky130_fd_sc_hd__a21o_2 _7224_ (.A1(_2593_),
    .A2(_2598_),
    .B1(_2605_),
    .X(_2612_));
 sky130_fd_sc_hd__o21ai_2 _7225_ (.A1(net160),
    .A2(net106),
    .B1(_2459_),
    .Y(_2613_));
 sky130_fd_sc_hd__nand2_2 _7226_ (.A(_2571_),
    .B(_2613_),
    .Y(_2614_));
 sky130_fd_sc_hd__and3_4 _7227_ (.A(_2571_),
    .B(_2612_),
    .C(_2613_),
    .X(_2615_));
 sky130_fd_sc_hd__xnor2_4 _7228_ (.A(_2612_),
    .B(_2614_),
    .Y(_2616_));
 sky130_fd_sc_hd__xnor2_4 _7229_ (.A(_2590_),
    .B(_2610_),
    .Y(_2618_));
 sky130_fd_sc_hd__a21bo_4 _7230_ (.A1(_2616_),
    .A2(_2618_),
    .B1_N(_2611_),
    .X(_2619_));
 sky130_fd_sc_hd__nand2b_1 _7231_ (.A_N(_2589_),
    .B(_2619_),
    .Y(_2620_));
 sky130_fd_sc_hd__xnor2_4 _7232_ (.A(_2589_),
    .B(_2619_),
    .Y(_2621_));
 sky130_fd_sc_hd__a21boi_4 _7233_ (.A1(_2615_),
    .A2(_2621_),
    .B1_N(_2620_),
    .Y(_2622_));
 sky130_fd_sc_hd__xor2_4 _7234_ (.A(_2588_),
    .B(_2622_),
    .X(_2623_));
 sky130_fd_sc_hd__nor2_2 _7235_ (.A(net138),
    .B(net84),
    .Y(_2624_));
 sky130_fd_sc_hd__o2bb2a_2 _7236_ (.A1_N(_2623_),
    .A2_N(_2624_),
    .B1(_2588_),
    .B2(_2622_),
    .X(_2625_));
 sky130_fd_sc_hd__and2b_1 _7237_ (.A_N(_2625_),
    .B(_2587_),
    .X(_2626_));
 sky130_fd_sc_hd__xnor2_4 _7238_ (.A(_2587_),
    .B(_2625_),
    .Y(_2627_));
 sky130_fd_sc_hd__xor2_4 _7239_ (.A(_2623_),
    .B(_2624_),
    .X(_2629_));
 sky130_fd_sc_hd__xnor2_4 _7240_ (.A(_2615_),
    .B(_2621_),
    .Y(_2630_));
 sky130_fd_sc_hd__xnor2_4 _7241_ (.A(_2616_),
    .B(_2618_),
    .Y(_2631_));
 sky130_fd_sc_hd__and2_1 _7242_ (.A(_2607_),
    .B(_2608_),
    .X(_2632_));
 sky130_fd_sc_hd__or2_4 _7243_ (.A(_2609_),
    .B(_2632_),
    .X(_2633_));
 sky130_fd_sc_hd__xnor2_4 _7244_ (.A(_2594_),
    .B(_2596_),
    .Y(_2634_));
 sky130_fd_sc_hd__nor2_4 _7245_ (.A(net142),
    .B(net105),
    .Y(_2635_));
 sky130_fd_sc_hd__o22a_1 _7246_ (.A1(net175),
    .A2(net82),
    .B1(net75),
    .B2(net134),
    .X(_2636_));
 sky130_fd_sc_hd__or4_4 _7247_ (.A(net134),
    .B(net175),
    .C(net82),
    .D(net75),
    .X(_2637_));
 sky130_fd_sc_hd__and2b_2 _7248_ (.A_N(_2636_),
    .B(_2637_),
    .X(_2638_));
 sky130_fd_sc_hd__and2_2 _7249_ (.A(_2635_),
    .B(_2638_),
    .X(_2640_));
 sky130_fd_sc_hd__nand2_1 _7250_ (.A(_2634_),
    .B(_2640_),
    .Y(_2641_));
 sky130_fd_sc_hd__xnor2_4 _7251_ (.A(_2602_),
    .B(_2603_),
    .Y(_2642_));
 sky130_fd_sc_hd__xnor2_4 _7252_ (.A(_2637_),
    .B(_2642_),
    .Y(_2643_));
 sky130_fd_sc_hd__nand2_2 _7253_ (.A(net124),
    .B(net113),
    .Y(_2644_));
 sky130_fd_sc_hd__or3_4 _7254_ (.A(net178),
    .B(net79),
    .C(_2644_),
    .X(_2645_));
 sky130_fd_sc_hd__or2_1 _7255_ (.A(_2643_),
    .B(_2645_),
    .X(_2646_));
 sky130_fd_sc_hd__xnor2_4 _7256_ (.A(_2643_),
    .B(_2645_),
    .Y(_2647_));
 sky130_fd_sc_hd__xnor2_4 _7257_ (.A(_2634_),
    .B(_2640_),
    .Y(_2648_));
 sky130_fd_sc_hd__o21ai_4 _7258_ (.A1(_2647_),
    .A2(_2648_),
    .B1(_2641_),
    .Y(_2649_));
 sky130_fd_sc_hd__and2b_1 _7259_ (.A_N(_2633_),
    .B(_2649_),
    .X(_2651_));
 sky130_fd_sc_hd__o21a_2 _7260_ (.A1(_2637_),
    .A2(_2642_),
    .B1(_2646_),
    .X(_2652_));
 sky130_fd_sc_hd__or3_4 _7261_ (.A(net160),
    .B(net104),
    .C(_2652_),
    .X(_2653_));
 sky130_fd_sc_hd__xnor2_4 _7262_ (.A(_2570_),
    .B(_2652_),
    .Y(_2654_));
 sky130_fd_sc_hd__xnor2_4 _7263_ (.A(_2633_),
    .B(_2649_),
    .Y(_2655_));
 sky130_fd_sc_hd__a21oi_2 _7264_ (.A1(_2654_),
    .A2(_2655_),
    .B1(_2651_),
    .Y(_2656_));
 sky130_fd_sc_hd__or2_1 _7265_ (.A(_2631_),
    .B(_2656_),
    .X(_2657_));
 sky130_fd_sc_hd__xnor2_2 _7266_ (.A(_2631_),
    .B(_2656_),
    .Y(_2658_));
 sky130_fd_sc_hd__o21a_2 _7267_ (.A1(_2653_),
    .A2(_2658_),
    .B1(_2657_),
    .X(_2659_));
 sky130_fd_sc_hd__xnor2_4 _7268_ (.A(_2630_),
    .B(_2659_),
    .Y(_2660_));
 sky130_fd_sc_hd__nand2_2 _7269_ (.A(net140),
    .B(net83),
    .Y(_2662_));
 sky130_fd_sc_hd__o32a_1 _7270_ (.A1(net138),
    .A2(net82),
    .A3(_2660_),
    .B1(_2659_),
    .B2(_2630_),
    .X(_2663_));
 sky130_fd_sc_hd__nand2b_4 _7271_ (.A_N(_2663_),
    .B(_2629_),
    .Y(_2664_));
 sky130_fd_sc_hd__nand2b_1 _7272_ (.A_N(_2629_),
    .B(_2663_),
    .Y(_2665_));
 sky130_fd_sc_hd__nand2_4 _7273_ (.A(_2664_),
    .B(_2665_),
    .Y(_2666_));
 sky130_fd_sc_hd__xnor2_4 _7274_ (.A(_2660_),
    .B(_2662_),
    .Y(_2667_));
 sky130_fd_sc_hd__xor2_2 _7275_ (.A(_2653_),
    .B(_2658_),
    .X(_2668_));
 sky130_fd_sc_hd__xnor2_4 _7276_ (.A(_2654_),
    .B(_2655_),
    .Y(_2669_));
 sky130_fd_sc_hd__xnor2_4 _7277_ (.A(_2647_),
    .B(_2648_),
    .Y(_2670_));
 sky130_fd_sc_hd__xnor2_4 _7278_ (.A(_2635_),
    .B(_2638_),
    .Y(_2671_));
 sky130_fd_sc_hd__a32o_1 _7279_ (.A1(net170),
    .A2(_1990_),
    .A3(net124),
    .B1(net113),
    .B2(net181),
    .X(_2673_));
 sky130_fd_sc_hd__o31a_4 _7280_ (.A1(net178),
    .A2(net79),
    .A3(_2644_),
    .B1(_2673_),
    .X(_2674_));
 sky130_fd_sc_hd__and4_4 _7281_ (.A(net136),
    .B(_3702_),
    .C(net80),
    .D(net113),
    .X(_2675_));
 sky130_fd_sc_hd__nand2_1 _7282_ (.A(_2674_),
    .B(_2675_),
    .Y(_2676_));
 sky130_fd_sc_hd__xor2_4 _7283_ (.A(_2674_),
    .B(_2675_),
    .X(_2677_));
 sky130_fd_sc_hd__or2_2 _7284_ (.A(net123),
    .B(net106),
    .X(_2678_));
 sky130_fd_sc_hd__and3_2 _7285_ (.A(net124),
    .B(net73),
    .C(_2600_),
    .X(_2679_));
 sky130_fd_sc_hd__xnor2_4 _7286_ (.A(_2677_),
    .B(_2679_),
    .Y(_2680_));
 sky130_fd_sc_hd__or2_4 _7287_ (.A(_2671_),
    .B(_2680_),
    .X(_2681_));
 sky130_fd_sc_hd__nor2_1 _7288_ (.A(_2670_),
    .B(_2681_),
    .Y(_2682_));
 sky130_fd_sc_hd__a21bo_2 _7289_ (.A1(_2677_),
    .A2(_2679_),
    .B1_N(_2676_),
    .X(_2684_));
 sky130_fd_sc_hd__xor2_4 _7290_ (.A(_2670_),
    .B(_2681_),
    .X(_2685_));
 sky130_fd_sc_hd__a21o_2 _7291_ (.A1(_2684_),
    .A2(_2685_),
    .B1(_2682_),
    .X(_2686_));
 sky130_fd_sc_hd__and2b_1 _7292_ (.A_N(_2669_),
    .B(_2686_),
    .X(_2687_));
 sky130_fd_sc_hd__xnor2_1 _7293_ (.A(_2668_),
    .B(_2687_),
    .Y(_2688_));
 sky130_fd_sc_hd__or3_1 _7294_ (.A(net138),
    .B(net79),
    .C(_2688_),
    .X(_2689_));
 sky130_fd_sc_hd__a21bo_2 _7295_ (.A1(_2668_),
    .A2(_2687_),
    .B1_N(_2689_),
    .X(_2690_));
 sky130_fd_sc_hd__and2b_1 _7296_ (.A_N(_2667_),
    .B(_2690_),
    .X(_2691_));
 sky130_fd_sc_hd__xnor2_4 _7297_ (.A(_2667_),
    .B(_2690_),
    .Y(_2692_));
 sky130_fd_sc_hd__o21ai_1 _7298_ (.A1(net138),
    .A2(net79),
    .B1(_2688_),
    .Y(_2693_));
 sky130_fd_sc_hd__nand2_1 _7299_ (.A(_2689_),
    .B(_2693_),
    .Y(_2695_));
 sky130_fd_sc_hd__xor2_4 _7300_ (.A(_2669_),
    .B(_2686_),
    .X(_2696_));
 sky130_fd_sc_hd__xnor2_2 _7301_ (.A(_2684_),
    .B(_2685_),
    .Y(_2697_));
 sky130_fd_sc_hd__xor2_4 _7302_ (.A(_2671_),
    .B(_2680_),
    .X(_2698_));
 sky130_fd_sc_hd__o22a_1 _7303_ (.A1(net175),
    .A2(net79),
    .B1(net110),
    .B2(net134),
    .X(_2699_));
 sky130_fd_sc_hd__or2_4 _7304_ (.A(_2675_),
    .B(_2699_),
    .X(_2700_));
 sky130_fd_sc_hd__nor2_1 _7305_ (.A(net176),
    .B(net106),
    .Y(_2701_));
 sky130_fd_sc_hd__and3_4 _7306_ (.A(net136),
    .B(net77),
    .C(_2701_),
    .X(_2702_));
 sky130_fd_sc_hd__o32a_2 _7307_ (.A1(net173),
    .A2(net123),
    .A3(_0495_),
    .B1(net106),
    .B2(net178),
    .X(_2703_));
 sky130_fd_sc_hd__a31oi_4 _7308_ (.A1(net124),
    .A2(net73),
    .A3(_2600_),
    .B1(_2703_),
    .Y(_2704_));
 sky130_fd_sc_hd__nand2_1 _7309_ (.A(_2702_),
    .B(_2704_),
    .Y(_2706_));
 sky130_fd_sc_hd__xnor2_4 _7310_ (.A(_2702_),
    .B(_2704_),
    .Y(_2707_));
 sky130_fd_sc_hd__or3_4 _7311_ (.A(net178),
    .B(net104),
    .C(_2644_),
    .X(_2708_));
 sky130_fd_sc_hd__xor2_4 _7312_ (.A(_2707_),
    .B(_2708_),
    .X(_2709_));
 sky130_fd_sc_hd__and2b_1 _7313_ (.A_N(_2700_),
    .B(_2709_),
    .X(_2710_));
 sky130_fd_sc_hd__nand2_1 _7314_ (.A(_2698_),
    .B(_2710_),
    .Y(_2711_));
 sky130_fd_sc_hd__o21a_2 _7315_ (.A1(_2707_),
    .A2(_2708_),
    .B1(_2706_),
    .X(_2712_));
 sky130_fd_sc_hd__xnor2_2 _7316_ (.A(_2698_),
    .B(_2710_),
    .Y(_2713_));
 sky130_fd_sc_hd__o21a_1 _7317_ (.A1(_2712_),
    .A2(_2713_),
    .B1(_2711_),
    .X(_2714_));
 sky130_fd_sc_hd__nor2_2 _7318_ (.A(_2697_),
    .B(_2714_),
    .Y(_2715_));
 sky130_fd_sc_hd__nand2_2 _7319_ (.A(net140),
    .B(net77),
    .Y(_2717_));
 sky130_fd_sc_hd__xnor2_2 _7320_ (.A(_2696_),
    .B(_2715_),
    .Y(_2718_));
 sky130_fd_sc_hd__nand2b_1 _7321_ (.A_N(_2717_),
    .B(_2718_),
    .Y(_2719_));
 sky130_fd_sc_hd__o31a_1 _7322_ (.A1(_2696_),
    .A2(_2697_),
    .A3(_2714_),
    .B1(_2719_),
    .X(_2720_));
 sky130_fd_sc_hd__nor2_1 _7323_ (.A(_2695_),
    .B(_2720_),
    .Y(_2721_));
 sky130_fd_sc_hd__nand2_1 _7324_ (.A(_2695_),
    .B(_2720_),
    .Y(_2722_));
 sky130_fd_sc_hd__nand2b_1 _7325_ (.A_N(_2721_),
    .B(_2722_),
    .Y(_2723_));
 sky130_fd_sc_hd__xnor2_2 _7326_ (.A(_2717_),
    .B(_2718_),
    .Y(_2724_));
 sky130_fd_sc_hd__and2_1 _7327_ (.A(_2697_),
    .B(_2714_),
    .X(_2725_));
 sky130_fd_sc_hd__or2_4 _7328_ (.A(_2715_),
    .B(_2725_),
    .X(_2726_));
 sky130_fd_sc_hd__xnor2_2 _7329_ (.A(_2712_),
    .B(_2713_),
    .Y(_2728_));
 sky130_fd_sc_hd__xnor2_4 _7330_ (.A(_2700_),
    .B(_2709_),
    .Y(_2729_));
 sky130_fd_sc_hd__o22a_1 _7331_ (.A1(net176),
    .A2(net75),
    .B1(net106),
    .B2(_3509_),
    .X(_2730_));
 sky130_fd_sc_hd__nor2_2 _7332_ (.A(_2702_),
    .B(_2730_),
    .Y(_2731_));
 sky130_fd_sc_hd__nor2_1 _7333_ (.A(net176),
    .B(net104),
    .Y(_2732_));
 sky130_fd_sc_hd__or4_4 _7334_ (.A(net135),
    .B(net174),
    .C(net110),
    .D(net104),
    .X(_2733_));
 sky130_fd_sc_hd__o21ai_1 _7335_ (.A1(net178),
    .A2(net104),
    .B1(_2644_),
    .Y(_2734_));
 sky130_fd_sc_hd__and2_4 _7336_ (.A(_2708_),
    .B(_2734_),
    .X(_2735_));
 sky130_fd_sc_hd__nand2b_4 _7337_ (.A_N(_2733_),
    .B(_2735_),
    .Y(_2736_));
 sky130_fd_sc_hd__xnor2_4 _7338_ (.A(_2733_),
    .B(_2735_),
    .Y(_2737_));
 sky130_fd_sc_hd__nand2_4 _7339_ (.A(_2731_),
    .B(_2737_),
    .Y(_2739_));
 sky130_fd_sc_hd__xnor2_4 _7340_ (.A(_2729_),
    .B(_2739_),
    .Y(_2740_));
 sky130_fd_sc_hd__a21boi_4 _7341_ (.A1(_2736_),
    .A2(_2739_),
    .B1_N(_2729_),
    .Y(_2741_));
 sky130_fd_sc_hd__and2b_2 _7342_ (.A_N(_2728_),
    .B(_2741_),
    .X(_2742_));
 sky130_fd_sc_hd__and2b_1 _7343_ (.A_N(_2726_),
    .B(_2742_),
    .X(_2743_));
 sky130_fd_sc_hd__nor2_2 _7344_ (.A(net138),
    .B(net110),
    .Y(_2744_));
 sky130_fd_sc_hd__xnor2_4 _7345_ (.A(_2726_),
    .B(_2742_),
    .Y(_2745_));
 sky130_fd_sc_hd__a21oi_2 _7346_ (.A1(_2744_),
    .A2(_2745_),
    .B1(_2743_),
    .Y(_2746_));
 sky130_fd_sc_hd__and2b_1 _7347_ (.A_N(_2746_),
    .B(_2724_),
    .X(_2747_));
 sky130_fd_sc_hd__xnor2_2 _7348_ (.A(_2724_),
    .B(_2746_),
    .Y(_2748_));
 sky130_fd_sc_hd__xnor2_2 _7349_ (.A(_2744_),
    .B(_2745_),
    .Y(_2750_));
 sky130_fd_sc_hd__xnor2_2 _7350_ (.A(_2728_),
    .B(_2741_),
    .Y(_2751_));
 sky130_fd_sc_hd__xnor2_4 _7351_ (.A(_2736_),
    .B(_2740_),
    .Y(_2752_));
 sky130_fd_sc_hd__xnor2_2 _7352_ (.A(_2731_),
    .B(_2737_),
    .Y(_2753_));
 sky130_fd_sc_hd__a22o_1 _7353_ (.A1(_3702_),
    .A2(net113),
    .B1(_0587_),
    .B2(net137),
    .X(_2754_));
 sky130_fd_sc_hd__nand2_2 _7354_ (.A(_2733_),
    .B(_2754_),
    .Y(_2755_));
 sky130_fd_sc_hd__or3_1 _7355_ (.A(_2678_),
    .B(_2753_),
    .C(_2755_),
    .X(_2756_));
 sky130_fd_sc_hd__inv_2 _7356_ (.A(_2756_),
    .Y(_2757_));
 sky130_fd_sc_hd__nand2_1 _7357_ (.A(_2752_),
    .B(_2757_),
    .Y(_2758_));
 sky130_fd_sc_hd__or2_1 _7358_ (.A(net138),
    .B(net107),
    .X(_2759_));
 sky130_fd_sc_hd__xor2_1 _7359_ (.A(_2751_),
    .B(_2758_),
    .X(_2761_));
 sky130_fd_sc_hd__nor2_1 _7360_ (.A(_2759_),
    .B(_2761_),
    .Y(_2762_));
 sky130_fd_sc_hd__a31o_2 _7361_ (.A1(_2751_),
    .A2(_2752_),
    .A3(_2757_),
    .B1(_2762_),
    .X(_2763_));
 sky130_fd_sc_hd__and2b_1 _7362_ (.A_N(_2750_),
    .B(_2763_),
    .X(_2764_));
 sky130_fd_sc_hd__and2_1 _7363_ (.A(_2759_),
    .B(_2761_),
    .X(_2765_));
 sky130_fd_sc_hd__or2_1 _7364_ (.A(_2762_),
    .B(_2765_),
    .X(_2766_));
 sky130_fd_sc_hd__xor2_1 _7365_ (.A(_2678_),
    .B(_2755_),
    .X(_2767_));
 sky130_fd_sc_hd__or4b_1 _7366_ (.A(net176),
    .B(net104),
    .C(_2678_),
    .D_N(_2767_),
    .X(_2768_));
 sky130_fd_sc_hd__nor2_1 _7367_ (.A(_2753_),
    .B(_2768_),
    .Y(_2769_));
 sky130_fd_sc_hd__nand2_1 _7368_ (.A(_2752_),
    .B(_2769_),
    .Y(_2770_));
 sky130_fd_sc_hd__or2_1 _7369_ (.A(_2757_),
    .B(_2769_),
    .X(_2772_));
 sky130_fd_sc_hd__xnor2_1 _7370_ (.A(_2752_),
    .B(_2772_),
    .Y(_2773_));
 sky130_fd_sc_hd__or3_1 _7371_ (.A(net138),
    .B(net104),
    .C(_2773_),
    .X(_2774_));
 sky130_fd_sc_hd__a21o_1 _7372_ (.A1(_2770_),
    .A2(_2774_),
    .B1(_2766_),
    .X(_2775_));
 sky130_fd_sc_hd__inv_2 _7373_ (.A(_2775_),
    .Y(_2776_));
 sky130_fd_sc_hd__xnor2_2 _7374_ (.A(_2750_),
    .B(_2763_),
    .Y(_2777_));
 sky130_fd_sc_hd__a21o_1 _7375_ (.A1(_2776_),
    .A2(_2777_),
    .B1(_2764_),
    .X(_2778_));
 sky130_fd_sc_hd__a21o_1 _7376_ (.A1(_2748_),
    .A2(_2778_),
    .B1(_2747_),
    .X(_2779_));
 sky130_fd_sc_hd__a21o_2 _7377_ (.A1(_2722_),
    .A2(_2779_),
    .B1(_2721_),
    .X(_2780_));
 sky130_fd_sc_hd__a21oi_4 _7378_ (.A1(_2692_),
    .A2(_2780_),
    .B1(_2691_),
    .Y(_2781_));
 sky130_fd_sc_hd__o21ai_4 _7379_ (.A1(_2666_),
    .A2(_2781_),
    .B1(_2664_),
    .Y(_2783_));
 sky130_fd_sc_hd__a21oi_4 _7380_ (.A1(_2627_),
    .A2(_2783_),
    .B1(_2626_),
    .Y(_2784_));
 sky130_fd_sc_hd__o21ai_4 _7381_ (.A1(_2585_),
    .A2(_2784_),
    .B1(_2582_),
    .Y(_2785_));
 sky130_fd_sc_hd__a21oi_4 _7382_ (.A1(_2536_),
    .A2(_2785_),
    .B1(_2534_),
    .Y(_2786_));
 sky130_fd_sc_hd__o21ai_2 _7383_ (.A1(_2482_),
    .A2(_2786_),
    .B1(_2480_),
    .Y(_2787_));
 sky130_fd_sc_hd__a21oi_2 _7384_ (.A1(_2420_),
    .A2(_2787_),
    .B1(_2417_),
    .Y(_2788_));
 sky130_fd_sc_hd__o21bai_2 _7385_ (.A1(_2355_),
    .A2(_2788_),
    .B1_N(_2354_),
    .Y(_2789_));
 sky130_fd_sc_hd__a21oi_1 _7386_ (.A1(_2297_),
    .A2(_2789_),
    .B1(_2294_),
    .Y(_2790_));
 sky130_fd_sc_hd__and2b_1 _7387_ (.A_N(_2790_),
    .B(_2247_),
    .X(_2791_));
 sky130_fd_sc_hd__o21bai_2 _7388_ (.A1(_2213_),
    .A2(_2246_),
    .B1_N(_2791_),
    .Y(_2792_));
 sky130_fd_sc_hd__a21oi_2 _7389_ (.A1(_2163_),
    .A2(_2212_),
    .B1(_2170_),
    .Y(_2794_));
 sky130_fd_sc_hd__a31oi_4 _7390_ (.A1(_2163_),
    .A2(_2170_),
    .A3(_2212_),
    .B1(_2794_),
    .Y(_2795_));
 sky130_fd_sc_hd__a2bb2o_1 _7391_ (.A1_N(_2170_),
    .A2_N(_2212_),
    .B1(_2792_),
    .B2(_2795_),
    .X(_2796_));
 sky130_fd_sc_hd__or3_1 _7392_ (.A(_2173_),
    .B(_2175_),
    .C(_2176_),
    .X(_2797_));
 sky130_fd_sc_hd__a21o_1 _7393_ (.A1(_2171_),
    .A2(_2179_),
    .B1(_2797_),
    .X(_2798_));
 sky130_fd_sc_hd__a21o_1 _7394_ (.A1(_2180_),
    .A2(_2796_),
    .B1(_2798_),
    .X(_2799_));
 sky130_fd_sc_hd__a21o_1 _7395_ (.A1(_1652_),
    .A2(net40),
    .B1(_1650_),
    .X(_2800_));
 sky130_fd_sc_hd__a21o_2 _7396_ (.A1(_1607_),
    .A2(_2800_),
    .B1(_1606_),
    .X(_2801_));
 sky130_fd_sc_hd__a21o_4 _7397_ (.A1(_1271_),
    .A2(_2801_),
    .B1(_1272_),
    .X(_2802_));
 sky130_fd_sc_hd__xnor2_4 _7398_ (.A(_1266_),
    .B(_2802_),
    .Y(_2803_));
 sky130_fd_sc_hd__clkinv_2 _7399_ (.A(_2803_),
    .Y(_2805_));
 sky130_fd_sc_hd__xnor2_2 _7400_ (.A(_1273_),
    .B(_2801_),
    .Y(_2806_));
 sky130_fd_sc_hd__xor2_2 _7401_ (.A(_1607_),
    .B(_2800_),
    .X(_2807_));
 sky130_fd_sc_hd__xnor2_4 _7402_ (.A(_1651_),
    .B(net40),
    .Y(_2808_));
 sky130_fd_sc_hd__or4_4 _7403_ (.A(_2803_),
    .B(_2806_),
    .C(_2807_),
    .D(_2808_),
    .X(_2809_));
 sky130_fd_sc_hd__inv_2 _7404_ (.A(_2809_),
    .Y(_2810_));
 sky130_fd_sc_hd__a21oi_4 _7405_ (.A1(_1262_),
    .A2(_2802_),
    .B1(_1263_),
    .Y(_2811_));
 sky130_fd_sc_hd__o21bai_4 _7406_ (.A1(_1293_),
    .A2(_2811_),
    .B1_N(_1290_),
    .Y(_2812_));
 sky130_fd_sc_hd__a21o_2 _7407_ (.A1(_1309_),
    .A2(_2812_),
    .B1(_1305_),
    .X(_2813_));
 sky130_fd_sc_hd__a21o_2 _7408_ (.A1(_1327_),
    .A2(_2813_),
    .B1(_1324_),
    .X(_2814_));
 sky130_fd_sc_hd__o32a_4 _7409_ (.A1(net212),
    .A2(net201),
    .A3(_1333_),
    .B1(_1335_),
    .B2(_2814_),
    .X(_2816_));
 sky130_fd_sc_hd__inv_2 _7410_ (.A(_2816_),
    .Y(_2817_));
 sky130_fd_sc_hd__xnor2_4 _7411_ (.A(_2805_),
    .B(_2816_),
    .Y(_2818_));
 sky130_fd_sc_hd__nor2_2 _7412_ (.A(_2810_),
    .B(_2818_),
    .Y(_2819_));
 sky130_fd_sc_hd__xor2_4 _7413_ (.A(_1293_),
    .B(_2811_),
    .X(_2820_));
 sky130_fd_sc_hd__or2_4 _7414_ (.A(_2810_),
    .B(_2816_),
    .X(_2821_));
 sky130_fd_sc_hd__xnor2_4 _7415_ (.A(_2820_),
    .B(_2821_),
    .Y(_2822_));
 sky130_fd_sc_hd__xnor2_4 _7416_ (.A(_1310_),
    .B(_2812_),
    .Y(_2823_));
 sky130_fd_sc_hd__o21a_1 _7417_ (.A1(_2809_),
    .A2(_2820_),
    .B1(_2817_),
    .X(_2824_));
 sky130_fd_sc_hd__xnor2_2 _7418_ (.A(_2823_),
    .B(_2824_),
    .Y(_2825_));
 sky130_fd_sc_hd__or4b_4 _7419_ (.A(_2810_),
    .B(_2825_),
    .C(_2818_),
    .D_N(_2822_),
    .X(_2827_));
 sky130_fd_sc_hd__xnor2_4 _7420_ (.A(_1327_),
    .B(_2813_),
    .Y(_2828_));
 sky130_fd_sc_hd__nor3_2 _7421_ (.A(_2809_),
    .B(_2820_),
    .C(_2823_),
    .Y(_2829_));
 sky130_fd_sc_hd__or2_4 _7422_ (.A(_2816_),
    .B(_2829_),
    .X(_2830_));
 sky130_fd_sc_hd__xnor2_4 _7423_ (.A(_2828_),
    .B(_2830_),
    .Y(_2831_));
 sky130_fd_sc_hd__nand2_4 _7424_ (.A(_2827_),
    .B(_2831_),
    .Y(_2832_));
 sky130_fd_sc_hd__a21bo_1 _7425_ (.A1(_2828_),
    .A2(_2829_),
    .B1_N(_1334_),
    .X(_2833_));
 sky130_fd_sc_hd__nand3_2 _7426_ (.A(_1337_),
    .B(_2814_),
    .C(_2833_),
    .Y(_2834_));
 sky130_fd_sc_hd__a2111o_2 _7427_ (.A1(_2828_),
    .A2(_2829_),
    .B1(_1336_),
    .C1(_2814_),
    .D1(_2816_),
    .X(_2835_));
 sky130_fd_sc_hd__nand2_4 _7428_ (.A(_2834_),
    .B(_2835_),
    .Y(_2836_));
 sky130_fd_sc_hd__nor2_8 _7429_ (.A(_2832_),
    .B(_2836_),
    .Y(_2838_));
 sky130_fd_sc_hd__or2_1 _7430_ (.A(_2832_),
    .B(_2836_),
    .X(_2839_));
 sky130_fd_sc_hd__a21bo_1 _7431_ (.A1(_2819_),
    .A2(_2822_),
    .B1_N(_2825_),
    .X(_2840_));
 sky130_fd_sc_hd__o21bai_4 _7432_ (.A1(_2827_),
    .A2(_2831_),
    .B1_N(_2836_),
    .Y(_2841_));
 sky130_fd_sc_hd__a21o_1 _7433_ (.A1(_2827_),
    .A2(_2840_),
    .B1(_2841_),
    .X(_2842_));
 sky130_fd_sc_hd__clkinv_4 _7434_ (.A(net31),
    .Y(_2843_));
 sky130_fd_sc_hd__a32o_1 _7435_ (.A1(_2818_),
    .A2(_2822_),
    .A3(_2832_),
    .B1(net32),
    .B2(net31),
    .X(_2844_));
 sky130_fd_sc_hd__xor2_2 _7436_ (.A(_2819_),
    .B(_2822_),
    .X(_2845_));
 sky130_fd_sc_hd__nor2_1 _7437_ (.A(_2841_),
    .B(_2845_),
    .Y(_2846_));
 sky130_fd_sc_hd__or2_1 _7438_ (.A(_2818_),
    .B(_2841_),
    .X(_2847_));
 sky130_fd_sc_hd__xor2_1 _7439_ (.A(_2482_),
    .B(_2786_),
    .X(_2849_));
 sky130_fd_sc_hd__xor2_1 _7440_ (.A(_2420_),
    .B(_2787_),
    .X(_2850_));
 sky130_fd_sc_hd__mux2_1 _7441_ (.A0(_2849_),
    .A1(_2850_),
    .S(net41),
    .X(_2851_));
 sky130_fd_sc_hd__xor2_1 _7442_ (.A(_2355_),
    .B(_2788_),
    .X(_2852_));
 sky130_fd_sc_hd__mux2_1 _7443_ (.A0(_2850_),
    .A1(_2852_),
    .S(net41),
    .X(_2853_));
 sky130_fd_sc_hd__mux2_1 _7444_ (.A0(_2851_),
    .A1(_2853_),
    .S(net27),
    .X(_2854_));
 sky130_fd_sc_hd__xnor2_1 _7445_ (.A(_2296_),
    .B(_2789_),
    .Y(_2855_));
 sky130_fd_sc_hd__mux2_1 _7446_ (.A0(_2852_),
    .A1(_2855_),
    .S(net41),
    .X(_2856_));
 sky130_fd_sc_hd__and2b_1 _7447_ (.A_N(_2247_),
    .B(_2790_),
    .X(_2857_));
 sky130_fd_sc_hd__nor2_1 _7448_ (.A(_2791_),
    .B(_2857_),
    .Y(_2858_));
 sky130_fd_sc_hd__mux2_1 _7449_ (.A0(_2855_),
    .A1(_2858_),
    .S(net41),
    .X(_2860_));
 sky130_fd_sc_hd__mux2_1 _7450_ (.A0(_2856_),
    .A1(_2860_),
    .S(net27),
    .X(_2861_));
 sky130_fd_sc_hd__mux2_1 _7451_ (.A0(_2861_),
    .A1(_2854_),
    .S(net28),
    .X(_2862_));
 sky130_fd_sc_hd__xor2_1 _7452_ (.A(_2792_),
    .B(_2795_),
    .X(_2863_));
 sky130_fd_sc_hd__mux2_1 _7453_ (.A0(_2858_),
    .A1(_2863_),
    .S(net41),
    .X(_2864_));
 sky130_fd_sc_hd__or2_1 _7454_ (.A(_2180_),
    .B(_2796_),
    .X(_2865_));
 sky130_fd_sc_hd__mux2_1 _7455_ (.A0(_2863_),
    .A1(_2865_),
    .S(_2798_),
    .X(_2866_));
 sky130_fd_sc_hd__mux2_1 _7456_ (.A0(_2864_),
    .A1(_2866_),
    .S(net27),
    .X(_2867_));
 sky130_fd_sc_hd__nand2b_1 _7457_ (.A_N(_2807_),
    .B(net27),
    .Y(_2868_));
 sky130_fd_sc_hd__o21ai_2 _7458_ (.A1(_2808_),
    .A2(net27),
    .B1(_2868_),
    .Y(_2869_));
 sky130_fd_sc_hd__inv_2 _7459_ (.A(_2869_),
    .Y(_2871_));
 sky130_fd_sc_hd__mux2_2 _7460_ (.A0(_2871_),
    .A1(_2867_),
    .S(net29),
    .X(_2872_));
 sky130_fd_sc_hd__mux2_1 _7461_ (.A0(_2862_),
    .A1(_2872_),
    .S(net30),
    .X(_2873_));
 sky130_fd_sc_hd__inv_2 _7462_ (.A(_2873_),
    .Y(_2874_));
 sky130_fd_sc_hd__mux2_1 _7463_ (.A0(_2853_),
    .A1(_2856_),
    .S(net27),
    .X(_2875_));
 sky130_fd_sc_hd__mux2_1 _7464_ (.A0(_2860_),
    .A1(_2864_),
    .S(net27),
    .X(_2876_));
 sky130_fd_sc_hd__mux2_1 _7465_ (.A0(_2876_),
    .A1(_2875_),
    .S(net29),
    .X(_2877_));
 sky130_fd_sc_hd__mux2_1 _7466_ (.A0(_2866_),
    .A1(_2808_),
    .S(net27),
    .X(_2878_));
 sky130_fd_sc_hd__mux2_1 _7467_ (.A0(_2807_),
    .A1(_2806_),
    .S(net26),
    .X(_2879_));
 sky130_fd_sc_hd__mux2_1 _7468_ (.A0(_2879_),
    .A1(_2878_),
    .S(net29),
    .X(_2880_));
 sky130_fd_sc_hd__mux2_1 _7469_ (.A0(_2877_),
    .A1(_2880_),
    .S(net30),
    .X(_2882_));
 sky130_fd_sc_hd__inv_2 _7470_ (.A(_2882_),
    .Y(_2883_));
 sky130_fd_sc_hd__xor2_2 _7471_ (.A(_2666_),
    .B(_2781_),
    .X(_2884_));
 sky130_fd_sc_hd__xor2_2 _7472_ (.A(_2627_),
    .B(_2783_),
    .X(_2885_));
 sky130_fd_sc_hd__mux2_1 _7473_ (.A0(_2884_),
    .A1(_2885_),
    .S(net40),
    .X(_2886_));
 sky130_fd_sc_hd__xor2_2 _7474_ (.A(_2585_),
    .B(_2784_),
    .X(_2887_));
 sky130_fd_sc_hd__mux2_1 _7475_ (.A0(_2885_),
    .A1(_2887_),
    .S(net40),
    .X(_2888_));
 sky130_fd_sc_hd__mux2_1 _7476_ (.A0(_2886_),
    .A1(_2888_),
    .S(net25),
    .X(_2889_));
 sky130_fd_sc_hd__xor2_2 _7477_ (.A(_2536_),
    .B(_2785_),
    .X(_2890_));
 sky130_fd_sc_hd__mux2_1 _7478_ (.A0(_2887_),
    .A1(_2890_),
    .S(net40),
    .X(_2891_));
 sky130_fd_sc_hd__mux2_1 _7479_ (.A0(_2890_),
    .A1(_2849_),
    .S(net40),
    .X(_2893_));
 sky130_fd_sc_hd__mux2_1 _7480_ (.A0(_2891_),
    .A1(_2893_),
    .S(net25),
    .X(_2894_));
 sky130_fd_sc_hd__mux2_1 _7481_ (.A0(_2894_),
    .A1(_2889_),
    .S(net28),
    .X(_2895_));
 sky130_fd_sc_hd__mux2_1 _7482_ (.A0(_2862_),
    .A1(_2895_),
    .S(_2843_),
    .X(_2896_));
 sky130_fd_sc_hd__mux2_1 _7483_ (.A0(_2893_),
    .A1(_2851_),
    .S(net25),
    .X(_2897_));
 sky130_fd_sc_hd__mux2_1 _7484_ (.A0(_2875_),
    .A1(_2897_),
    .S(net29),
    .X(_2898_));
 sky130_fd_sc_hd__mux2_1 _7485_ (.A0(_2878_),
    .A1(_2876_),
    .S(net28),
    .X(_2899_));
 sky130_fd_sc_hd__mux2_1 _7486_ (.A0(_2898_),
    .A1(_2899_),
    .S(net30),
    .X(_2900_));
 sky130_fd_sc_hd__xnor2_1 _7487_ (.A(_2723_),
    .B(_2779_),
    .Y(_2901_));
 sky130_fd_sc_hd__xor2_1 _7488_ (.A(_2692_),
    .B(_2780_),
    .X(_2902_));
 sky130_fd_sc_hd__mux2_1 _7489_ (.A0(_2901_),
    .A1(_2902_),
    .S(net40),
    .X(_2904_));
 sky130_fd_sc_hd__mux2_1 _7490_ (.A0(_2902_),
    .A1(_2884_),
    .S(net40),
    .X(_2905_));
 sky130_fd_sc_hd__mux2_1 _7491_ (.A0(_2904_),
    .A1(_2905_),
    .S(net25),
    .X(_2906_));
 sky130_fd_sc_hd__mux2_1 _7492_ (.A0(_2889_),
    .A1(_2906_),
    .S(net28),
    .X(_2907_));
 sky130_fd_sc_hd__mux2_1 _7493_ (.A0(_2854_),
    .A1(_2894_),
    .S(net28),
    .X(_2908_));
 sky130_fd_sc_hd__mux2_1 _7494_ (.A0(_2907_),
    .A1(_2908_),
    .S(net31),
    .X(_2909_));
 sky130_fd_sc_hd__inv_2 _7495_ (.A(_2909_),
    .Y(_2910_));
 sky130_fd_sc_hd__mux2_1 _7496_ (.A0(_2888_),
    .A1(_2891_),
    .S(net26),
    .X(_2911_));
 sky130_fd_sc_hd__mux2_1 _7497_ (.A0(_2897_),
    .A1(_2911_),
    .S(net28),
    .X(_2912_));
 sky130_fd_sc_hd__mux2_2 _7498_ (.A0(_2877_),
    .A1(_2912_),
    .S(_2843_),
    .X(_2913_));
 sky130_fd_sc_hd__mux2_1 _7499_ (.A0(_2867_),
    .A1(_2861_),
    .S(net29),
    .X(_2915_));
 sky130_fd_sc_hd__inv_2 _7500_ (.A(_2915_),
    .Y(_2916_));
 sky130_fd_sc_hd__mux2_2 _7501_ (.A0(_2908_),
    .A1(_2915_),
    .S(net30),
    .X(_2917_));
 sky130_fd_sc_hd__nand2_1 _7502_ (.A(_2816_),
    .B(net26),
    .Y(_2918_));
 sky130_fd_sc_hd__o31ai_1 _7503_ (.A1(_2803_),
    .A2(_2816_),
    .A3(_2841_),
    .B1(_2918_),
    .Y(_2919_));
 sky130_fd_sc_hd__mux2_1 _7504_ (.A0(_2919_),
    .A1(_2879_),
    .S(net29),
    .X(_2920_));
 sky130_fd_sc_hd__mux2_2 _7505_ (.A0(_2899_),
    .A1(_2920_),
    .S(net30),
    .X(_2921_));
 sky130_fd_sc_hd__mux2_1 _7506_ (.A0(_2905_),
    .A1(_2886_),
    .S(net25),
    .X(_2922_));
 sky130_fd_sc_hd__mux2_1 _7507_ (.A0(_2911_),
    .A1(_2922_),
    .S(net28),
    .X(_2923_));
 sky130_fd_sc_hd__xor2_1 _7508_ (.A(_2748_),
    .B(_2778_),
    .X(_2924_));
 sky130_fd_sc_hd__mux2_1 _7509_ (.A0(_2924_),
    .A1(_2901_),
    .S(net40),
    .X(_2926_));
 sky130_fd_sc_hd__mux2_1 _7510_ (.A0(_2926_),
    .A1(_2904_),
    .S(net25),
    .X(_2927_));
 sky130_fd_sc_hd__mux2_1 _7511_ (.A0(_2922_),
    .A1(_2927_),
    .S(net28),
    .X(_2928_));
 sky130_fd_sc_hd__xnor2_1 _7512_ (.A(_2775_),
    .B(_2777_),
    .Y(_2929_));
 sky130_fd_sc_hd__mux2_1 _7513_ (.A0(_2929_),
    .A1(_2924_),
    .S(net41),
    .X(_2930_));
 sky130_fd_sc_hd__mux2_1 _7514_ (.A0(_2930_),
    .A1(_2926_),
    .S(net25),
    .X(_2931_));
 sky130_fd_sc_hd__mux2_1 _7515_ (.A0(_2906_),
    .A1(_2931_),
    .S(net28),
    .X(_2932_));
 sky130_fd_sc_hd__and3_1 _7516_ (.A(_2766_),
    .B(_2770_),
    .C(_2774_),
    .X(_2933_));
 sky130_fd_sc_hd__nor2_1 _7517_ (.A(_2776_),
    .B(_2933_),
    .Y(_2934_));
 sky130_fd_sc_hd__o21ai_1 _7518_ (.A1(net138),
    .A2(net104),
    .B1(_2773_),
    .Y(_2935_));
 sky130_fd_sc_hd__o211a_1 _7519_ (.A1(_2678_),
    .A2(_2755_),
    .B1(_2768_),
    .C1(_2753_),
    .X(_2937_));
 sky130_fd_sc_hd__a2111oi_1 _7520_ (.A1(_3510_),
    .A2(_0587_),
    .B1(_2701_),
    .C1(_2732_),
    .D1(_2767_),
    .Y(_2938_));
 sky130_fd_sc_hd__o21ai_1 _7521_ (.A1(_2772_),
    .A2(_2937_),
    .B1(_2938_),
    .Y(_2939_));
 sky130_fd_sc_hd__a21o_1 _7522_ (.A1(_2774_),
    .A2(_2935_),
    .B1(_2939_),
    .X(_2940_));
 sky130_fd_sc_hd__a211o_1 _7523_ (.A1(net40),
    .A2(_2929_),
    .B1(_2934_),
    .C1(_2940_),
    .X(_2941_));
 sky130_fd_sc_hd__nand2_1 _7524_ (.A(_2843_),
    .B(_2845_),
    .Y(_2942_));
 sky130_fd_sc_hd__inv_2 _7525_ (.A(_2942_),
    .Y(_2943_));
 sky130_fd_sc_hd__o21ba_1 _7526_ (.A1(_2927_),
    .A2(_2931_),
    .B1_N(net28),
    .X(_2944_));
 sky130_fd_sc_hd__mux2_1 _7527_ (.A0(_2941_),
    .A1(_2930_),
    .S(net25),
    .X(_2945_));
 sky130_fd_sc_hd__a21o_1 _7528_ (.A1(net25),
    .A2(_2930_),
    .B1(_2941_),
    .X(_2946_));
 sky130_fd_sc_hd__or2_1 _7529_ (.A(net31),
    .B(_2946_),
    .X(_2948_));
 sky130_fd_sc_hd__a21o_1 _7530_ (.A1(_2942_),
    .A2(_2948_),
    .B1(_2944_),
    .X(_2949_));
 sky130_fd_sc_hd__or4_1 _7531_ (.A(_2843_),
    .B(_2907_),
    .C(_2923_),
    .D(_2928_),
    .X(_2950_));
 sky130_fd_sc_hd__a22o_1 _7532_ (.A1(_2943_),
    .A2(_2945_),
    .B1(_2949_),
    .B2(_2950_),
    .X(_2951_));
 sky130_fd_sc_hd__mux2_1 _7533_ (.A0(_2895_),
    .A1(_2932_),
    .S(_2843_),
    .X(_2952_));
 sky130_fd_sc_hd__and2_1 _7534_ (.A(_2843_),
    .B(_2928_),
    .X(_2953_));
 sky130_fd_sc_hd__and2_1 _7535_ (.A(net31),
    .B(_2912_),
    .X(_2954_));
 sky130_fd_sc_hd__or4_1 _7536_ (.A(net33),
    .B(_2952_),
    .C(_2953_),
    .D(_2954_),
    .X(_2955_));
 sky130_fd_sc_hd__or4_1 _7537_ (.A(_2838_),
    .B(_2873_),
    .C(_2882_),
    .D(_2951_),
    .X(_2956_));
 sky130_fd_sc_hd__mux2_1 _7538_ (.A0(_2898_),
    .A1(_2923_),
    .S(_2843_),
    .X(_2957_));
 sky130_fd_sc_hd__or2_2 _7539_ (.A(net33),
    .B(_2957_),
    .X(_2959_));
 sky130_fd_sc_hd__o21ai_4 _7540_ (.A1(_2838_),
    .A2(_2921_),
    .B1(_2959_),
    .Y(_2960_));
 sky130_fd_sc_hd__o21ai_1 _7541_ (.A1(_2944_),
    .A2(_2946_),
    .B1(net31),
    .Y(_2961_));
 sky130_fd_sc_hd__or4_1 _7542_ (.A(_2909_),
    .B(_2917_),
    .C(_2952_),
    .D(_2957_),
    .X(_2962_));
 sky130_fd_sc_hd__or4_1 _7543_ (.A(_2838_),
    .B(_2953_),
    .C(_2954_),
    .D(_2962_),
    .X(_2963_));
 sky130_fd_sc_hd__or4_1 _7544_ (.A(_2896_),
    .B(_2900_),
    .C(_2913_),
    .D(_2963_),
    .X(_2964_));
 sky130_fd_sc_hd__a32o_1 _7545_ (.A1(net25),
    .A2(_2941_),
    .A3(_2943_),
    .B1(_2932_),
    .B2(net31),
    .X(_2965_));
 sky130_fd_sc_hd__o31a_1 _7546_ (.A1(net33),
    .A2(_2951_),
    .A3(_2965_),
    .B1(_2964_),
    .X(_2966_));
 sky130_fd_sc_hd__a21oi_1 _7547_ (.A1(_2955_),
    .A2(_2956_),
    .B1(_2966_),
    .Y(_2967_));
 sky130_fd_sc_hd__a31o_1 _7548_ (.A1(_2960_),
    .A2(_2961_),
    .A3(_2967_),
    .B1(_2844_),
    .X(_2968_));
 sky130_fd_sc_hd__o21ai_1 _7549_ (.A1(_2806_),
    .A2(net26),
    .B1(_2918_),
    .Y(_2970_));
 sky130_fd_sc_hd__mux2_1 _7550_ (.A0(_2970_),
    .A1(_2869_),
    .S(net29),
    .X(_2971_));
 sky130_fd_sc_hd__mux2_1 _7551_ (.A0(_2916_),
    .A1(_2971_),
    .S(net30),
    .X(_2972_));
 sky130_fd_sc_hd__mux2_2 _7552_ (.A0(_2910_),
    .A1(_2972_),
    .S(net32),
    .X(_2973_));
 sky130_fd_sc_hd__and2b_1 _7553_ (.A_N(_2973_),
    .B(_2968_),
    .X(_2974_));
 sky130_fd_sc_hd__or3_4 _7554_ (.A(_2844_),
    .B(_2960_),
    .C(_2973_),
    .X(_2975_));
 sky130_fd_sc_hd__o21ai_1 _7555_ (.A1(_2968_),
    .A2(_2973_),
    .B1(_2960_),
    .Y(_2976_));
 sky130_fd_sc_hd__and2_1 _7556_ (.A(_2975_),
    .B(_2976_),
    .X(_2977_));
 sky130_fd_sc_hd__a21oi_1 _7557_ (.A1(net222),
    .A2(_2974_),
    .B1(_2977_),
    .Y(_2978_));
 sky130_fd_sc_hd__or3b_2 _7558_ (.A(_1216_),
    .B(\cmd[7] ),
    .C_N(\cmd[6] ),
    .X(_2979_));
 sky130_fd_sc_hd__and3b_1 _7559_ (.A_N(_2960_),
    .B(_2974_),
    .C(net223),
    .X(_2981_));
 sky130_fd_sc_hd__o31a_1 _7560_ (.A1(_1559_),
    .A2(_1562_),
    .A3(_1563_),
    .B1(_2119_),
    .X(_2982_));
 sky130_fd_sc_hd__o31a_1 _7561_ (.A1(_2978_),
    .A2(net182),
    .A3(_2981_),
    .B1(_2982_),
    .X(_2983_));
 sky130_fd_sc_hd__and2b_1 _7562_ (.A_N(net228),
    .B(net239),
    .X(_2984_));
 sky130_fd_sc_hd__inv_2 _7563_ (.A(net220),
    .Y(_2985_));
 sky130_fd_sc_hd__o2bb2a_1 _7564_ (.A1_N(\out_reg[0] ),
    .A2_N(net219),
    .B1(_2983_),
    .B2(net239),
    .X(_2986_));
 sky130_fd_sc_hd__nor2_1 _7565_ (.A(net236),
    .B(_2986_),
    .Y(_0020_));
 sky130_fd_sc_hd__o211a_4 _7566_ (.A1(_1384_),
    .A2(_1556_),
    .B1(_1557_),
    .C1(_1552_),
    .X(_2987_));
 sky130_fd_sc_hd__nand2_8 _7567_ (.A(_1470_),
    .B(_2987_),
    .Y(_2988_));
 sky130_fd_sc_hd__or2_2 _7568_ (.A(_1470_),
    .B(_1558_),
    .X(_2989_));
 sky130_fd_sc_hd__and3_1 _7569_ (.A(net225),
    .B(_2988_),
    .C(_2989_),
    .X(_2991_));
 sky130_fd_sc_hd__nand2_1 _7570_ (.A(_1350_),
    .B(net11),
    .Y(_2992_));
 sky130_fd_sc_hd__o21a_2 _7571_ (.A1(net11),
    .A2(_1554_),
    .B1(_2992_),
    .X(_2993_));
 sky130_fd_sc_hd__o211a_1 _7572_ (.A1(net11),
    .A2(_1554_),
    .B1(_2992_),
    .C1(net6),
    .X(_2994_));
 sky130_fd_sc_hd__a211o_1 _7573_ (.A1(_1412_),
    .A2(_1503_),
    .B1(_2994_),
    .C1(_1384_),
    .X(_2995_));
 sky130_fd_sc_hd__a21boi_4 _7574_ (.A1(_1384_),
    .A2(_1490_),
    .B1_N(_2995_),
    .Y(_2996_));
 sky130_fd_sc_hd__nand3_4 _7575_ (.A(_1470_),
    .B(_2987_),
    .C(_2996_),
    .Y(_2997_));
 sky130_fd_sc_hd__xnor2_4 _7576_ (.A(_2988_),
    .B(_2996_),
    .Y(_2998_));
 sky130_fd_sc_hd__nand2_1 _7577_ (.A(_2991_),
    .B(_2996_),
    .Y(_2999_));
 sky130_fd_sc_hd__o211a_2 _7578_ (.A1(_2991_),
    .A2(_2998_),
    .B1(_2999_),
    .C1(_1560_),
    .X(_3000_));
 sky130_fd_sc_hd__and2_2 _7579_ (.A(_2107_),
    .B(_2110_),
    .X(_3002_));
 sky130_fd_sc_hd__and3b_1 _7580_ (.A_N(_2106_),
    .B(_1970_),
    .C(_2101_),
    .X(_3003_));
 sky130_fd_sc_hd__mux2_1 _7581_ (.A0(_2103_),
    .A1(_1930_),
    .S(net24),
    .X(_3004_));
 sky130_fd_sc_hd__inv_2 _7582_ (.A(_3004_),
    .Y(_3005_));
 sky130_fd_sc_hd__mux2_1 _7583_ (.A0(_2074_),
    .A1(_3005_),
    .S(net19),
    .X(_3006_));
 sky130_fd_sc_hd__mux2_1 _7584_ (.A0(_2038_),
    .A1(_3006_),
    .S(net16),
    .X(_3007_));
 sky130_fd_sc_hd__nand2_1 _7585_ (.A(_3003_),
    .B(_3007_),
    .Y(_3008_));
 sky130_fd_sc_hd__or2_1 _7586_ (.A(_3003_),
    .B(_3007_),
    .X(_3009_));
 sky130_fd_sc_hd__nand2_1 _7587_ (.A(_3008_),
    .B(_3009_),
    .Y(_3010_));
 sky130_fd_sc_hd__or3_1 _7588_ (.A(_2108_),
    .B(_3002_),
    .C(_3010_),
    .X(_3011_));
 sky130_fd_sc_hd__o21ai_1 _7589_ (.A1(net72),
    .A2(_3002_),
    .B1(_3010_),
    .Y(_3013_));
 sky130_fd_sc_hd__or2_1 _7590_ (.A(_2974_),
    .B(_2977_),
    .X(_3014_));
 sky130_fd_sc_hd__mux2_1 _7591_ (.A0(_2817_),
    .A1(_2970_),
    .S(net29),
    .X(_3015_));
 sky130_fd_sc_hd__nand2_1 _7592_ (.A(net30),
    .B(_3015_),
    .Y(_3016_));
 sky130_fd_sc_hd__o21ai_4 _7593_ (.A1(net30),
    .A2(_2872_),
    .B1(_3016_),
    .Y(_3017_));
 sky130_fd_sc_hd__inv_2 _7594_ (.A(_3017_),
    .Y(_3018_));
 sky130_fd_sc_hd__mux2_4 _7595_ (.A0(_2896_),
    .A1(_3018_),
    .S(net33),
    .X(_3019_));
 sky130_fd_sc_hd__nand2b_2 _7596_ (.A_N(_2975_),
    .B(_3019_),
    .Y(_3020_));
 sky130_fd_sc_hd__xnor2_2 _7597_ (.A(_2975_),
    .B(_3019_),
    .Y(_3021_));
 sky130_fd_sc_hd__and3_1 _7598_ (.A(net222),
    .B(_3014_),
    .C(_3021_),
    .X(_3022_));
 sky130_fd_sc_hd__a21oi_1 _7599_ (.A1(net222),
    .A2(_3014_),
    .B1(_3021_),
    .Y(_3024_));
 sky130_fd_sc_hd__nor3_1 _7600_ (.A(net182),
    .B(_3022_),
    .C(_3024_),
    .Y(_3025_));
 sky130_fd_sc_hd__a31o_1 _7601_ (.A1(_2116_),
    .A2(_3011_),
    .A3(_3013_),
    .B1(net241),
    .X(_3026_));
 sky130_fd_sc_hd__a21bo_1 _7602_ (.A1(\out_reg[0] ),
    .A2(_0775_),
    .B1_N(net239),
    .X(_3027_));
 sky130_fd_sc_hd__o31a_1 _7603_ (.A1(_3000_),
    .A2(_3025_),
    .A3(_3026_),
    .B1(_3027_),
    .X(_3028_));
 sky130_fd_sc_hd__a21oi_1 _7604_ (.A1(\out_reg[1] ),
    .A2(net219),
    .B1(_3028_),
    .Y(_3029_));
 sky130_fd_sc_hd__nor2_1 _7605_ (.A(net236),
    .B(_3029_),
    .Y(_0021_));
 sky130_fd_sc_hd__a21o_1 _7606_ (.A1(_2988_),
    .A2(_2989_),
    .B1(_2998_),
    .X(_3030_));
 sky130_fd_sc_hd__and2_1 _7607_ (.A(net225),
    .B(_3030_),
    .X(_3031_));
 sky130_fd_sc_hd__o21ai_1 _7608_ (.A1(_1270_),
    .A2(net11),
    .B1(_2992_),
    .Y(_3032_));
 sky130_fd_sc_hd__mux2_1 _7609_ (.A0(_1510_),
    .A1(_3032_),
    .S(net6),
    .X(_3034_));
 sky130_fd_sc_hd__mux2_4 _7610_ (.A0(_1513_),
    .A1(_3034_),
    .S(net14),
    .X(_3035_));
 sky130_fd_sc_hd__and4b_4 _7611_ (.A_N(_3035_),
    .B(_2996_),
    .C(_2987_),
    .D(_1470_),
    .X(_3036_));
 sky130_fd_sc_hd__xor2_4 _7612_ (.A(_2997_),
    .B(_3035_),
    .X(_3037_));
 sky130_fd_sc_hd__o21ai_1 _7613_ (.A1(_3031_),
    .A2(_3037_),
    .B1(_1560_),
    .Y(_3038_));
 sky130_fd_sc_hd__a21oi_2 _7614_ (.A1(_3031_),
    .A2(_3037_),
    .B1(_3038_),
    .Y(_3039_));
 sky130_fd_sc_hd__and2_1 _7615_ (.A(_3002_),
    .B(_3010_),
    .X(_3040_));
 sky130_fd_sc_hd__mux2_2 _7616_ (.A0(_1961_),
    .A1(_2063_),
    .S(_1959_),
    .X(_3041_));
 sky130_fd_sc_hd__inv_2 _7617_ (.A(_3041_),
    .Y(_3042_));
 sky130_fd_sc_hd__mux2_1 _7618_ (.A0(_2054_),
    .A1(_3042_),
    .S(net16),
    .X(_3043_));
 sky130_fd_sc_hd__and3_4 _7619_ (.A(_3003_),
    .B(_3007_),
    .C(_3043_),
    .X(_3045_));
 sky130_fd_sc_hd__xor2_1 _7620_ (.A(_3008_),
    .B(_3043_),
    .X(_3046_));
 sky130_fd_sc_hd__o21ai_1 _7621_ (.A1(_2108_),
    .A2(_3040_),
    .B1(_3046_),
    .Y(_3047_));
 sky130_fd_sc_hd__or3_1 _7622_ (.A(net72),
    .B(_3040_),
    .C(_3046_),
    .X(_3048_));
 sky130_fd_sc_hd__nor2_1 _7623_ (.A(_3014_),
    .B(_3021_),
    .Y(_3049_));
 sky130_fd_sc_hd__mux2_1 _7624_ (.A0(_2816_),
    .A1(_2805_),
    .S(net29),
    .X(_3050_));
 sky130_fd_sc_hd__mux2_1 _7625_ (.A0(_2880_),
    .A1(_3050_),
    .S(net31),
    .X(_3051_));
 sky130_fd_sc_hd__or2_2 _7626_ (.A(_2838_),
    .B(_3051_),
    .X(_3052_));
 sky130_fd_sc_hd__o21ai_4 _7627_ (.A1(net33),
    .A2(_2913_),
    .B1(_3052_),
    .Y(_3053_));
 sky130_fd_sc_hd__nor2_4 _7628_ (.A(_3020_),
    .B(_3053_),
    .Y(_3054_));
 sky130_fd_sc_hd__and2_1 _7629_ (.A(_3020_),
    .B(_3053_),
    .X(_3056_));
 sky130_fd_sc_hd__or2_1 _7630_ (.A(_3054_),
    .B(_3056_),
    .X(_3057_));
 sky130_fd_sc_hd__o21a_1 _7631_ (.A1(net221),
    .A2(_3049_),
    .B1(_3057_),
    .X(_3058_));
 sky130_fd_sc_hd__nor2_1 _7632_ (.A(net182),
    .B(_3058_),
    .Y(_3059_));
 sky130_fd_sc_hd__o31a_1 _7633_ (.A1(net221),
    .A2(_3049_),
    .A3(_3057_),
    .B1(_3059_),
    .X(_3060_));
 sky130_fd_sc_hd__a31o_1 _7634_ (.A1(_2116_),
    .A2(_3047_),
    .A3(_3048_),
    .B1(net241),
    .X(_3061_));
 sky130_fd_sc_hd__a21bo_1 _7635_ (.A1(\out_reg[1] ),
    .A2(_0775_),
    .B1_N(net239),
    .X(_3062_));
 sky130_fd_sc_hd__o31a_2 _7636_ (.A1(_3039_),
    .A2(_3060_),
    .A3(_3061_),
    .B1(_3062_),
    .X(_3063_));
 sky130_fd_sc_hd__a21oi_1 _7637_ (.A1(\out_reg[2] ),
    .A2(net219),
    .B1(_3063_),
    .Y(_3064_));
 sky130_fd_sc_hd__nor2_1 _7638_ (.A(net236),
    .B(_3064_),
    .Y(_0022_));
 sky130_fd_sc_hd__nand2_4 _7639_ (.A(_1350_),
    .B(net6),
    .Y(_3066_));
 sky130_fd_sc_hd__o21a_2 _7640_ (.A1(net6),
    .A2(_1555_),
    .B1(_3066_),
    .X(_3067_));
 sky130_fd_sc_hd__inv_2 _7641_ (.A(_3067_),
    .Y(_3068_));
 sky130_fd_sc_hd__mux2_8 _7642_ (.A0(_1483_),
    .A1(_3068_),
    .S(net15),
    .X(_3069_));
 sky130_fd_sc_hd__or3_4 _7643_ (.A(_2997_),
    .B(_3035_),
    .C(_3069_),
    .X(_3070_));
 sky130_fd_sc_hd__xnor2_4 _7644_ (.A(_3036_),
    .B(_3069_),
    .Y(_3071_));
 sky130_fd_sc_hd__o21a_1 _7645_ (.A1(_3030_),
    .A2(_3037_),
    .B1(net225),
    .X(_3072_));
 sky130_fd_sc_hd__a21oi_1 _7646_ (.A1(_3071_),
    .A2(_3072_),
    .B1(_1562_),
    .Y(_3073_));
 sky130_fd_sc_hd__o21ai_2 _7647_ (.A1(_3071_),
    .A2(_3072_),
    .B1(_3073_),
    .Y(_3074_));
 sky130_fd_sc_hd__and3_1 _7648_ (.A(_3002_),
    .B(_3010_),
    .C(_3046_),
    .X(_3075_));
 sky130_fd_sc_hd__or2_1 _7649_ (.A(net72),
    .B(_3075_),
    .X(_3077_));
 sky130_fd_sc_hd__a21o_1 _7650_ (.A1(_1959_),
    .A2(_2104_),
    .B1(_1960_),
    .X(_3078_));
 sky130_fd_sc_hd__inv_2 _7651_ (.A(_3078_),
    .Y(_3079_));
 sky130_fd_sc_hd__mux2_4 _7652_ (.A0(_2070_),
    .A1(_3079_),
    .S(net16),
    .X(_3080_));
 sky130_fd_sc_hd__xnor2_2 _7653_ (.A(_3045_),
    .B(_3080_),
    .Y(_3081_));
 sky130_fd_sc_hd__nor2_1 _7654_ (.A(_3077_),
    .B(_3081_),
    .Y(_3082_));
 sky130_fd_sc_hd__a211o_1 _7655_ (.A1(_3077_),
    .A2(_3081_),
    .B1(_3082_),
    .C1(_2117_),
    .X(_3083_));
 sky130_fd_sc_hd__nand2_1 _7656_ (.A(_3049_),
    .B(_3057_),
    .Y(_3084_));
 sky130_fd_sc_hd__nand2_1 _7657_ (.A(_2817_),
    .B(net30),
    .Y(_3085_));
 sky130_fd_sc_hd__a21boi_2 _7658_ (.A1(_2843_),
    .A2(_2971_),
    .B1_N(_3085_),
    .Y(_3086_));
 sky130_fd_sc_hd__mux2_4 _7659_ (.A0(_2917_),
    .A1(_3086_),
    .S(net32),
    .X(_3088_));
 sky130_fd_sc_hd__xor2_2 _7660_ (.A(_3054_),
    .B(_3088_),
    .X(_3089_));
 sky130_fd_sc_hd__a21oi_1 _7661_ (.A1(net223),
    .A2(_3084_),
    .B1(_3089_),
    .Y(_3090_));
 sky130_fd_sc_hd__a31o_1 _7662_ (.A1(net223),
    .A2(_3084_),
    .A3(_3089_),
    .B1(net183),
    .X(_3091_));
 sky130_fd_sc_hd__or2_1 _7663_ (.A(_3090_),
    .B(_3091_),
    .X(_3092_));
 sky130_fd_sc_hd__a31o_2 _7664_ (.A1(_3074_),
    .A2(_3083_),
    .A3(_3092_),
    .B1(net241),
    .X(_3093_));
 sky130_fd_sc_hd__a22oi_1 _7665_ (.A1(\out_reg[2] ),
    .A2(_0786_),
    .B1(net219),
    .B2(\out_reg[3] ),
    .Y(_3094_));
 sky130_fd_sc_hd__a21oi_1 _7666_ (.A1(_3093_),
    .A2(_3094_),
    .B1(net236),
    .Y(_0023_));
 sky130_fd_sc_hd__o21ai_2 _7667_ (.A1(net6),
    .A2(_1453_),
    .B1(_3066_),
    .Y(_3095_));
 sky130_fd_sc_hd__o211a_1 _7668_ (.A1(net6),
    .A2(_1453_),
    .B1(_3066_),
    .C1(net14),
    .X(_3096_));
 sky130_fd_sc_hd__a21oi_4 _7669_ (.A1(_1384_),
    .A2(_1514_),
    .B1(_3096_),
    .Y(_3098_));
 sky130_fd_sc_hd__or3b_4 _7670_ (.A(_3069_),
    .B(_3098_),
    .C_N(_3036_),
    .X(_3099_));
 sky130_fd_sc_hd__xor2_4 _7671_ (.A(_3070_),
    .B(_3098_),
    .X(_3100_));
 sky130_fd_sc_hd__a2111oi_4 _7672_ (.A1(_2988_),
    .A2(_2989_),
    .B1(_2998_),
    .C1(_3037_),
    .D1(_3071_),
    .Y(_3101_));
 sky130_fd_sc_hd__or2_4 _7673_ (.A(net221),
    .B(_3101_),
    .X(_3102_));
 sky130_fd_sc_hd__xnor2_4 _7674_ (.A(_3100_),
    .B(_3102_),
    .Y(_3103_));
 sky130_fd_sc_hd__o21ba_1 _7675_ (.A1(net19),
    .A2(_2088_),
    .B1_N(_1960_),
    .X(_3104_));
 sky130_fd_sc_hd__mux2_2 _7676_ (.A0(_2087_),
    .A1(_3104_),
    .S(net16),
    .X(_3105_));
 sky130_fd_sc_hd__nand3_4 _7677_ (.A(_3045_),
    .B(_3080_),
    .C(_3105_),
    .Y(_3106_));
 sky130_fd_sc_hd__a21o_1 _7678_ (.A1(_3045_),
    .A2(_3080_),
    .B1(_3105_),
    .X(_3107_));
 sky130_fd_sc_hd__and2_1 _7679_ (.A(_3106_),
    .B(_3107_),
    .X(_3109_));
 sky130_fd_sc_hd__a21oi_1 _7680_ (.A1(_3075_),
    .A2(_3081_),
    .B1(net72),
    .Y(_3110_));
 sky130_fd_sc_hd__nand2_1 _7681_ (.A(_3109_),
    .B(_3110_),
    .Y(_3111_));
 sky130_fd_sc_hd__or2_1 _7682_ (.A(_3109_),
    .B(_3110_),
    .X(_3112_));
 sky130_fd_sc_hd__and3_1 _7683_ (.A(_2116_),
    .B(_3111_),
    .C(_3112_),
    .X(_3113_));
 sky130_fd_sc_hd__nor2_1 _7684_ (.A(_3084_),
    .B(_3089_),
    .Y(_3114_));
 sky130_fd_sc_hd__o21a_2 _7685_ (.A1(net30),
    .A2(_2920_),
    .B1(_3085_),
    .X(_3115_));
 sky130_fd_sc_hd__mux2_2 _7686_ (.A0(_2900_),
    .A1(_3115_),
    .S(net32),
    .X(_3116_));
 sky130_fd_sc_hd__nand3_2 _7687_ (.A(_3054_),
    .B(_3088_),
    .C(_3116_),
    .Y(_3117_));
 sky130_fd_sc_hd__a21o_1 _7688_ (.A1(_3054_),
    .A2(_3088_),
    .B1(_3116_),
    .X(_3118_));
 sky130_fd_sc_hd__nand2_1 _7689_ (.A(_3117_),
    .B(_3118_),
    .Y(_3120_));
 sky130_fd_sc_hd__o21a_1 _7690_ (.A1(net221),
    .A2(_3114_),
    .B1(_3120_),
    .X(_3121_));
 sky130_fd_sc_hd__nor2_1 _7691_ (.A(net182),
    .B(_3121_),
    .Y(_3122_));
 sky130_fd_sc_hd__o31a_2 _7692_ (.A1(net221),
    .A2(_3114_),
    .A3(_3120_),
    .B1(_3122_),
    .X(_3123_));
 sky130_fd_sc_hd__a2111oi_4 _7693_ (.A1(_1560_),
    .A2(_3103_),
    .B1(_3113_),
    .C1(_3123_),
    .D1(net241),
    .Y(_3124_));
 sky130_fd_sc_hd__a21boi_1 _7694_ (.A1(\out_reg[3] ),
    .A2(net228),
    .B1_N(net239),
    .Y(_3125_));
 sky130_fd_sc_hd__o2bb2a_1 _7695_ (.A1_N(\out_reg[4] ),
    .A2_N(net219),
    .B1(_3124_),
    .B2(_3125_),
    .X(_3126_));
 sky130_fd_sc_hd__nor2_1 _7696_ (.A(net236),
    .B(_3126_),
    .Y(_0024_));
 sky130_fd_sc_hd__nand2b_1 _7697_ (.A_N(_3100_),
    .B(_3101_),
    .Y(_3127_));
 sky130_fd_sc_hd__o21a_1 _7698_ (.A1(net6),
    .A2(_2993_),
    .B1(_3066_),
    .X(_3128_));
 sky130_fd_sc_hd__o211ai_4 _7699_ (.A1(net6),
    .A2(_2993_),
    .B1(_3066_),
    .C1(net14),
    .Y(_3130_));
 sky130_fd_sc_hd__o21ai_4 _7700_ (.A1(net14),
    .A2(_1505_),
    .B1(_3130_),
    .Y(_3131_));
 sky130_fd_sc_hd__nand2b_1 _7701_ (.A_N(_3098_),
    .B(_3131_),
    .Y(_3132_));
 sky130_fd_sc_hd__or3b_1 _7702_ (.A(_3069_),
    .B(_3132_),
    .C_N(_3036_),
    .X(_3133_));
 sky130_fd_sc_hd__xnor2_4 _7703_ (.A(_3099_),
    .B(_3131_),
    .Y(_3134_));
 sky130_fd_sc_hd__a21oi_1 _7704_ (.A1(net224),
    .A2(_3127_),
    .B1(_3134_),
    .Y(_3135_));
 sky130_fd_sc_hd__a31o_1 _7705_ (.A1(net225),
    .A2(_3127_),
    .A3(_3134_),
    .B1(_1562_),
    .X(_3136_));
 sky130_fd_sc_hd__or2_1 _7706_ (.A(_3135_),
    .B(_3136_),
    .X(_3137_));
 sky130_fd_sc_hd__nand2_1 _7707_ (.A(_3114_),
    .B(_3120_),
    .Y(_3138_));
 sky130_fd_sc_hd__a21boi_1 _7708_ (.A1(_2843_),
    .A2(_3015_),
    .B1_N(_3085_),
    .Y(_3139_));
 sky130_fd_sc_hd__inv_2 _7709_ (.A(_3139_),
    .Y(_3141_));
 sky130_fd_sc_hd__mux2_2 _7710_ (.A0(_2874_),
    .A1(_3141_),
    .S(net32),
    .X(_3142_));
 sky130_fd_sc_hd__nor2_2 _7711_ (.A(_3117_),
    .B(_3142_),
    .Y(_3143_));
 sky130_fd_sc_hd__and2_1 _7712_ (.A(_3117_),
    .B(_3142_),
    .X(_3144_));
 sky130_fd_sc_hd__nor2_1 _7713_ (.A(_3143_),
    .B(_3144_),
    .Y(_3145_));
 sky130_fd_sc_hd__a21oi_1 _7714_ (.A1(net223),
    .A2(_3138_),
    .B1(_3145_),
    .Y(_3146_));
 sky130_fd_sc_hd__a311o_1 _7715_ (.A1(net223),
    .A2(_3138_),
    .A3(_3145_),
    .B1(_3146_),
    .C1(net182),
    .X(_3147_));
 sky130_fd_sc_hd__a21o_1 _7716_ (.A1(_1959_),
    .A2(_3004_),
    .B1(_1960_),
    .X(_3148_));
 sky130_fd_sc_hd__inv_2 _7717_ (.A(_3148_),
    .Y(_3149_));
 sky130_fd_sc_hd__mux2_2 _7718_ (.A0(_2075_),
    .A1(_3149_),
    .S(net17),
    .X(_3150_));
 sky130_fd_sc_hd__and2b_1 _7719_ (.A_N(_3106_),
    .B(_3150_),
    .X(_3152_));
 sky130_fd_sc_hd__xnor2_2 _7720_ (.A(_3106_),
    .B(_3150_),
    .Y(_3153_));
 sky130_fd_sc_hd__and2_1 _7721_ (.A(_2109_),
    .B(_3112_),
    .X(_3154_));
 sky130_fd_sc_hd__o21ai_1 _7722_ (.A1(_3153_),
    .A2(_3154_),
    .B1(_2116_),
    .Y(_3155_));
 sky130_fd_sc_hd__a21o_1 _7723_ (.A1(_3153_),
    .A2(_3154_),
    .B1(_3155_),
    .X(_3156_));
 sky130_fd_sc_hd__a31o_2 _7724_ (.A1(_3137_),
    .A2(_3147_),
    .A3(_3156_),
    .B1(net241),
    .X(_3157_));
 sky130_fd_sc_hd__a22oi_1 _7725_ (.A1(\out_reg[4] ),
    .A2(_0786_),
    .B1(net219),
    .B2(\out_reg[5] ),
    .Y(_3158_));
 sky130_fd_sc_hd__a21oi_1 _7726_ (.A1(_3157_),
    .A2(_3158_),
    .B1(net236),
    .Y(_0025_));
 sky130_fd_sc_hd__or3b_1 _7727_ (.A(_3100_),
    .B(_3134_),
    .C_N(_3101_),
    .X(_3159_));
 sky130_fd_sc_hd__nand2_1 _7728_ (.A(net225),
    .B(_3159_),
    .Y(_3160_));
 sky130_fd_sc_hd__a21bo_1 _7729_ (.A1(_1412_),
    .A2(_3032_),
    .B1_N(_3066_),
    .X(_3162_));
 sky130_fd_sc_hd__mux2_1 _7730_ (.A0(_1511_),
    .A1(_3162_),
    .S(net15),
    .X(_3163_));
 sky130_fd_sc_hd__nor3b_1 _7731_ (.A(_3098_),
    .B(_3163_),
    .C_N(_3131_),
    .Y(_3164_));
 sky130_fd_sc_hd__and3b_1 _7732_ (.A_N(_3069_),
    .B(_3164_),
    .C(_3036_),
    .X(_3165_));
 sky130_fd_sc_hd__a21o_2 _7733_ (.A1(_3133_),
    .A2(_3163_),
    .B1(_3165_),
    .X(_3166_));
 sky130_fd_sc_hd__a21oi_1 _7734_ (.A1(_3160_),
    .A2(_3166_),
    .B1(_1562_),
    .Y(_3167_));
 sky130_fd_sc_hd__o21ai_2 _7735_ (.A1(_3160_),
    .A2(_3166_),
    .B1(_3167_),
    .Y(_3168_));
 sky130_fd_sc_hd__o21a_1 _7736_ (.A1(net16),
    .A2(_2064_),
    .B1(_1963_),
    .X(_3169_));
 sky130_fd_sc_hd__and2_1 _7737_ (.A(_3152_),
    .B(_3169_),
    .X(_3170_));
 sky130_fd_sc_hd__nor2_1 _7738_ (.A(_3152_),
    .B(_3169_),
    .Y(_3171_));
 sky130_fd_sc_hd__nor2_1 _7739_ (.A(_3170_),
    .B(_3171_),
    .Y(_3173_));
 sky130_fd_sc_hd__o21a_1 _7740_ (.A1(_3112_),
    .A2(_3153_),
    .B1(_2109_),
    .X(_3174_));
 sky130_fd_sc_hd__or2_1 _7741_ (.A(_3173_),
    .B(_3174_),
    .X(_3175_));
 sky130_fd_sc_hd__a21oi_1 _7742_ (.A1(_3173_),
    .A2(_3174_),
    .B1(_2117_),
    .Y(_3176_));
 sky130_fd_sc_hd__nand2_1 _7743_ (.A(_3175_),
    .B(_3176_),
    .Y(_3177_));
 sky130_fd_sc_hd__or2_1 _7744_ (.A(_3138_),
    .B(_3145_),
    .X(_3178_));
 sky130_fd_sc_hd__nand2_1 _7745_ (.A(net223),
    .B(_3178_),
    .Y(_3179_));
 sky130_fd_sc_hd__o21ai_1 _7746_ (.A1(net31),
    .A2(_3050_),
    .B1(_3085_),
    .Y(_3180_));
 sky130_fd_sc_hd__mux2_2 _7747_ (.A0(_2883_),
    .A1(_3180_),
    .S(net32),
    .X(_3181_));
 sky130_fd_sc_hd__or3_1 _7748_ (.A(_3117_),
    .B(_3142_),
    .C(_3181_),
    .X(_3182_));
 sky130_fd_sc_hd__xnor2_2 _7749_ (.A(_3143_),
    .B(_3181_),
    .Y(_3184_));
 sky130_fd_sc_hd__xor2_1 _7750_ (.A(_3179_),
    .B(_3184_),
    .X(_3185_));
 sky130_fd_sc_hd__o211a_2 _7751_ (.A1(net183),
    .A2(_3185_),
    .B1(_3177_),
    .C1(_3168_),
    .X(_3186_));
 sky130_fd_sc_hd__a22o_1 _7752_ (.A1(\out_reg[5] ),
    .A2(_0786_),
    .B1(net219),
    .B2(\out_reg[6] ),
    .X(_3187_));
 sky130_fd_sc_hd__o21ba_1 _7753_ (.A1(net239),
    .A2(_3186_),
    .B1_N(_3187_),
    .X(_3188_));
 sky130_fd_sc_hd__nor2_1 _7754_ (.A(net237),
    .B(_3188_),
    .Y(_0026_));
 sky130_fd_sc_hd__nor2_8 _7755_ (.A(_1349_),
    .B(_1384_),
    .Y(_3189_));
 sky130_fd_sc_hd__o21ba_1 _7756_ (.A1(net15),
    .A2(_1556_),
    .B1_N(_3189_),
    .X(_3190_));
 sky130_fd_sc_hd__and4b_4 _7757_ (.A_N(_3069_),
    .B(_3164_),
    .C(_3190_),
    .D(_3036_),
    .X(_3191_));
 sky130_fd_sc_hd__nor2_1 _7758_ (.A(_3165_),
    .B(_3190_),
    .Y(_3192_));
 sky130_fd_sc_hd__nor2_2 _7759_ (.A(_3191_),
    .B(_3192_),
    .Y(_3194_));
 sky130_fd_sc_hd__or4bb_4 _7760_ (.A(_3100_),
    .B(_3134_),
    .C_N(_3166_),
    .D_N(_3101_),
    .X(_3195_));
 sky130_fd_sc_hd__a21oi_1 _7761_ (.A1(net224),
    .A2(_3195_),
    .B1(_3194_),
    .Y(_3196_));
 sky130_fd_sc_hd__a31o_1 _7762_ (.A1(net225),
    .A2(_3194_),
    .A3(_3195_),
    .B1(_1562_),
    .X(_3197_));
 sky130_fd_sc_hd__or2_1 _7763_ (.A(_3196_),
    .B(_3197_),
    .X(_3198_));
 sky130_fd_sc_hd__nor2_1 _7764_ (.A(_3178_),
    .B(_3184_),
    .Y(_3199_));
 sky130_fd_sc_hd__or2_1 _7765_ (.A(net221),
    .B(_3199_),
    .X(_3200_));
 sky130_fd_sc_hd__nor2_4 _7766_ (.A(_2816_),
    .B(_2838_),
    .Y(_3201_));
 sky130_fd_sc_hd__a21o_1 _7767_ (.A1(_2838_),
    .A2(_2972_),
    .B1(_3201_),
    .X(_3202_));
 sky130_fd_sc_hd__or2_1 _7768_ (.A(_3182_),
    .B(_3202_),
    .X(_3203_));
 sky130_fd_sc_hd__nand2_1 _7769_ (.A(_3182_),
    .B(_3202_),
    .Y(_3205_));
 sky130_fd_sc_hd__nand2_1 _7770_ (.A(_3203_),
    .B(_3205_),
    .Y(_3206_));
 sky130_fd_sc_hd__a21oi_1 _7771_ (.A1(_3200_),
    .A2(_3206_),
    .B1(net183),
    .Y(_3207_));
 sky130_fd_sc_hd__o21ai_1 _7772_ (.A1(_3200_),
    .A2(_3206_),
    .B1(_3207_),
    .Y(_3208_));
 sky130_fd_sc_hd__and2_2 _7773_ (.A(_1930_),
    .B(net16),
    .X(_3209_));
 sky130_fd_sc_hd__a21oi_1 _7774_ (.A1(_1965_),
    .A2(_2105_),
    .B1(_3209_),
    .Y(_3210_));
 sky130_fd_sc_hd__and2_1 _7775_ (.A(_3170_),
    .B(_3210_),
    .X(_3211_));
 sky130_fd_sc_hd__nor2_1 _7776_ (.A(_3170_),
    .B(_3210_),
    .Y(_3212_));
 sky130_fd_sc_hd__nor2_1 _7777_ (.A(_3211_),
    .B(_3212_),
    .Y(_3213_));
 sky130_fd_sc_hd__a21oi_1 _7778_ (.A1(_2109_),
    .A2(_3175_),
    .B1(_3213_),
    .Y(_3214_));
 sky130_fd_sc_hd__a311o_1 _7779_ (.A1(_2109_),
    .A2(_3175_),
    .A3(_3213_),
    .B1(_3214_),
    .C1(_2117_),
    .X(_3216_));
 sky130_fd_sc_hd__a31o_2 _7780_ (.A1(_3198_),
    .A2(_3208_),
    .A3(_3216_),
    .B1(net241),
    .X(_3217_));
 sky130_fd_sc_hd__a22oi_1 _7781_ (.A1(\out_reg[6] ),
    .A2(_0786_),
    .B1(net220),
    .B2(\out_reg[7] ),
    .Y(_3218_));
 sky130_fd_sc_hd__a21oi_1 _7782_ (.A1(_3217_),
    .A2(_3218_),
    .B1(net236),
    .Y(_0027_));
 sky130_fd_sc_hd__o21a_1 _7783_ (.A1(_3194_),
    .A2(_3195_),
    .B1(net225),
    .X(_3219_));
 sky130_fd_sc_hd__or2_4 _7784_ (.A(net14),
    .B(_1469_),
    .X(_3220_));
 sky130_fd_sc_hd__o21bai_2 _7785_ (.A1(_3191_),
    .A2(_3220_),
    .B1_N(_3189_),
    .Y(_3221_));
 sky130_fd_sc_hd__a21oi_4 _7786_ (.A1(_3191_),
    .A2(_3220_),
    .B1(_3221_),
    .Y(_3222_));
 sky130_fd_sc_hd__xor2_1 _7787_ (.A(_3219_),
    .B(_3222_),
    .X(_3223_));
 sky130_fd_sc_hd__or2_1 _7788_ (.A(net16),
    .B(_2090_),
    .X(_3224_));
 sky130_fd_sc_hd__and3_2 _7789_ (.A(_3170_),
    .B(_3210_),
    .C(_3224_),
    .X(_3226_));
 sky130_fd_sc_hd__o21bai_1 _7790_ (.A1(_3211_),
    .A2(_3224_),
    .B1_N(_3209_),
    .Y(_3227_));
 sky130_fd_sc_hd__nor2_2 _7791_ (.A(_3226_),
    .B(_3227_),
    .Y(_3228_));
 sky130_fd_sc_hd__o31a_2 _7792_ (.A1(_3173_),
    .A2(_3174_),
    .A3(_3213_),
    .B1(_2109_),
    .X(_3229_));
 sky130_fd_sc_hd__nor2_4 _7793_ (.A(_3228_),
    .B(_3229_),
    .Y(_3230_));
 sky130_fd_sc_hd__a21o_1 _7794_ (.A1(_3228_),
    .A2(_3229_),
    .B1(_2117_),
    .X(_3231_));
 sky130_fd_sc_hd__nand2_1 _7795_ (.A(_3199_),
    .B(_3206_),
    .Y(_3232_));
 sky130_fd_sc_hd__nand2_1 _7796_ (.A(net223),
    .B(_3232_),
    .Y(_3233_));
 sky130_fd_sc_hd__nor2_1 _7797_ (.A(net33),
    .B(_2921_),
    .Y(_3234_));
 sky130_fd_sc_hd__or2_2 _7798_ (.A(_3203_),
    .B(_3234_),
    .X(_3235_));
 sky130_fd_sc_hd__o21ai_1 _7799_ (.A1(_3201_),
    .A2(_3234_),
    .B1(_3203_),
    .Y(_3237_));
 sky130_fd_sc_hd__and2_2 _7800_ (.A(_3235_),
    .B(_3237_),
    .X(_3238_));
 sky130_fd_sc_hd__xor2_2 _7801_ (.A(_3233_),
    .B(_3238_),
    .X(_3239_));
 sky130_fd_sc_hd__o22ai_1 _7802_ (.A1(_3230_),
    .A2(_3231_),
    .B1(_3239_),
    .B2(net183),
    .Y(_3240_));
 sky130_fd_sc_hd__a211o_2 _7803_ (.A1(_1560_),
    .A2(_3223_),
    .B1(_3240_),
    .C1(net241),
    .X(_3241_));
 sky130_fd_sc_hd__a21bo_1 _7804_ (.A1(\out_reg[7] ),
    .A2(net228),
    .B1_N(net239),
    .X(_3242_));
 sky130_fd_sc_hd__a22oi_1 _7805_ (.A1(\out_reg[8] ),
    .A2(net220),
    .B1(_3241_),
    .B2(_3242_),
    .Y(_3243_));
 sky130_fd_sc_hd__nor2_1 _7806_ (.A(net237),
    .B(_3243_),
    .Y(_0028_));
 sky130_fd_sc_hd__o31a_4 _7807_ (.A1(_3194_),
    .A2(_3195_),
    .A3(_3222_),
    .B1(net224),
    .X(_3244_));
 sky130_fd_sc_hd__a211o_4 _7808_ (.A1(_1412_),
    .A2(_1503_),
    .B1(_2994_),
    .C1(net14),
    .X(_3245_));
 sky130_fd_sc_hd__and2b_1 _7809_ (.A_N(_3189_),
    .B(_3245_),
    .X(_3247_));
 sky130_fd_sc_hd__a21oi_2 _7810_ (.A1(_3191_),
    .A2(_3220_),
    .B1(_3247_),
    .Y(_3248_));
 sky130_fd_sc_hd__a31oi_4 _7811_ (.A1(_3191_),
    .A2(_3220_),
    .A3(_3245_),
    .B1(_3248_),
    .Y(_3249_));
 sky130_fd_sc_hd__nand2_1 _7812_ (.A(_3244_),
    .B(_3249_),
    .Y(_3250_));
 sky130_fd_sc_hd__or2_1 _7813_ (.A(_3244_),
    .B(_3249_),
    .X(_3251_));
 sky130_fd_sc_hd__o21a_1 _7814_ (.A1(_3232_),
    .A2(_3238_),
    .B1(net223),
    .X(_3252_));
 sky130_fd_sc_hd__a21oi_4 _7815_ (.A1(_2838_),
    .A2(_3017_),
    .B1(_3201_),
    .Y(_3253_));
 sky130_fd_sc_hd__and2b_1 _7816_ (.A_N(_3235_),
    .B(_3253_),
    .X(_3254_));
 sky130_fd_sc_hd__xnor2_2 _7817_ (.A(_3235_),
    .B(_3253_),
    .Y(_3255_));
 sky130_fd_sc_hd__o21bai_1 _7818_ (.A1(_3252_),
    .A2(_3255_),
    .B1_N(net183),
    .Y(_3256_));
 sky130_fd_sc_hd__a21oi_1 _7819_ (.A1(_3252_),
    .A2(_3255_),
    .B1(_3256_),
    .Y(_3258_));
 sky130_fd_sc_hd__o21ba_1 _7820_ (.A1(net16),
    .A2(_3006_),
    .B1_N(_3209_),
    .X(_3259_));
 sky130_fd_sc_hd__nand2_2 _7821_ (.A(_3226_),
    .B(_3259_),
    .Y(_3260_));
 sky130_fd_sc_hd__or2_1 _7822_ (.A(_3226_),
    .B(_3259_),
    .X(_3261_));
 sky130_fd_sc_hd__nand2_2 _7823_ (.A(_3260_),
    .B(_3261_),
    .Y(_3262_));
 sky130_fd_sc_hd__o21ai_2 _7824_ (.A1(net72),
    .A2(_3230_),
    .B1(_3262_),
    .Y(_3263_));
 sky130_fd_sc_hd__o31a_2 _7825_ (.A1(net72),
    .A2(_3230_),
    .A3(_3262_),
    .B1(_2116_),
    .X(_3264_));
 sky130_fd_sc_hd__a31o_2 _7826_ (.A1(_1560_),
    .A2(_3250_),
    .A3(_3251_),
    .B1(_3258_),
    .X(_3265_));
 sky130_fd_sc_hd__a21oi_4 _7827_ (.A1(_3263_),
    .A2(_3264_),
    .B1(_3265_),
    .Y(_3266_));
 sky130_fd_sc_hd__a22o_1 _7828_ (.A1(\out_reg[8] ),
    .A2(_0786_),
    .B1(net220),
    .B2(\out_reg[9] ),
    .X(_3267_));
 sky130_fd_sc_hd__o21ba_1 _7829_ (.A1(net239),
    .A2(_3266_),
    .B1_N(_3267_),
    .X(_3269_));
 sky130_fd_sc_hd__nor2_1 _7830_ (.A(net237),
    .B(_3269_),
    .Y(_0029_));
 sky130_fd_sc_hd__and2_1 _7831_ (.A(_1384_),
    .B(_3034_),
    .X(_3270_));
 sky130_fd_sc_hd__inv_2 _7832_ (.A(_3270_),
    .Y(_3271_));
 sky130_fd_sc_hd__and4_4 _7833_ (.A(_3191_),
    .B(_3220_),
    .C(_3245_),
    .D(_3271_),
    .X(_3272_));
 sky130_fd_sc_hd__nor2_1 _7834_ (.A(_3189_),
    .B(_3270_),
    .Y(_3273_));
 sky130_fd_sc_hd__a31o_1 _7835_ (.A1(_3191_),
    .A2(_3220_),
    .A3(_3245_),
    .B1(_3273_),
    .X(_3274_));
 sky130_fd_sc_hd__and2b_1 _7836_ (.A_N(_3272_),
    .B(_3274_),
    .X(_3275_));
 sky130_fd_sc_hd__and2_1 _7837_ (.A(_1471_),
    .B(_3249_),
    .X(_3276_));
 sky130_fd_sc_hd__o21ai_1 _7838_ (.A1(_3244_),
    .A2(_3276_),
    .B1(_3275_),
    .Y(_3277_));
 sky130_fd_sc_hd__or3_1 _7839_ (.A(_3244_),
    .B(_3275_),
    .C(_3276_),
    .X(_3279_));
 sky130_fd_sc_hd__a21oi_2 _7840_ (.A1(_1965_),
    .A2(_3041_),
    .B1(_3260_),
    .Y(_3280_));
 sky130_fd_sc_hd__a31o_1 _7841_ (.A1(_1965_),
    .A2(_3041_),
    .A3(_3260_),
    .B1(_3209_),
    .X(_3281_));
 sky130_fd_sc_hd__or2_2 _7842_ (.A(_3280_),
    .B(_3281_),
    .X(_3282_));
 sky130_fd_sc_hd__a21o_1 _7843_ (.A1(_3230_),
    .A2(_3262_),
    .B1(net72),
    .X(_3283_));
 sky130_fd_sc_hd__nand2_1 _7844_ (.A(_3282_),
    .B(_3283_),
    .Y(_3284_));
 sky130_fd_sc_hd__o21a_1 _7845_ (.A1(_3282_),
    .A2(_3283_),
    .B1(_2116_),
    .X(_3285_));
 sky130_fd_sc_hd__o31a_1 _7846_ (.A1(_3232_),
    .A2(_3238_),
    .A3(_3255_),
    .B1(net223),
    .X(_3286_));
 sky130_fd_sc_hd__or2_1 _7847_ (.A(net32),
    .B(_3051_),
    .X(_3287_));
 sky130_fd_sc_hd__nand2_2 _7848_ (.A(_3254_),
    .B(_3287_),
    .Y(_3288_));
 sky130_fd_sc_hd__o221a_1 _7849_ (.A1(_2816_),
    .A2(_2838_),
    .B1(_3254_),
    .B2(_3287_),
    .C1(_3288_),
    .X(_3290_));
 sky130_fd_sc_hd__a21oi_1 _7850_ (.A1(_3286_),
    .A2(_3290_),
    .B1(net182),
    .Y(_3291_));
 sky130_fd_sc_hd__o21a_1 _7851_ (.A1(_3286_),
    .A2(_3290_),
    .B1(_3291_),
    .X(_3292_));
 sky130_fd_sc_hd__a211o_1 _7852_ (.A1(_3284_),
    .A2(_3285_),
    .B1(_3292_),
    .C1(net242),
    .X(_3293_));
 sky130_fd_sc_hd__a31o_2 _7853_ (.A1(_1560_),
    .A2(_3277_),
    .A3(_3279_),
    .B1(_3293_),
    .X(_3294_));
 sky130_fd_sc_hd__a21bo_1 _7854_ (.A1(\out_reg[9] ),
    .A2(net228),
    .B1_N(net240),
    .X(_3295_));
 sky130_fd_sc_hd__a22oi_1 _7855_ (.A1(\out_reg[10] ),
    .A2(net220),
    .B1(_3294_),
    .B2(_3295_),
    .Y(_3296_));
 sky130_fd_sc_hd__nor2_1 _7856_ (.A(net237),
    .B(_3296_),
    .Y(_0030_));
 sky130_fd_sc_hd__nand2_1 _7857_ (.A(\out_reg[11] ),
    .B(net219),
    .Y(_3297_));
 sky130_fd_sc_hd__or2_4 _7858_ (.A(net15),
    .B(_3067_),
    .X(_3298_));
 sky130_fd_sc_hd__xnor2_1 _7859_ (.A(_3272_),
    .B(_3298_),
    .Y(_3300_));
 sky130_fd_sc_hd__nor2_1 _7860_ (.A(_3189_),
    .B(_3300_),
    .Y(_3301_));
 sky130_fd_sc_hd__o21a_1 _7861_ (.A1(_3249_),
    .A2(_3275_),
    .B1(net224),
    .X(_3302_));
 sky130_fd_sc_hd__o21ai_1 _7862_ (.A1(_3244_),
    .A2(_3302_),
    .B1(_3301_),
    .Y(_3303_));
 sky130_fd_sc_hd__o311a_2 _7863_ (.A1(_3244_),
    .A2(_3301_),
    .A3(_3302_),
    .B1(_3303_),
    .C1(_1560_),
    .X(_3304_));
 sky130_fd_sc_hd__a21oi_1 _7864_ (.A1(_1965_),
    .A2(_3078_),
    .B1(_3209_),
    .Y(_3305_));
 sky130_fd_sc_hd__and2_1 _7865_ (.A(_3280_),
    .B(_3305_),
    .X(_3306_));
 sky130_fd_sc_hd__nor2_1 _7866_ (.A(_3280_),
    .B(_3305_),
    .Y(_3307_));
 sky130_fd_sc_hd__or2_1 _7867_ (.A(_3306_),
    .B(_3307_),
    .X(_3308_));
 sky130_fd_sc_hd__a31o_1 _7868_ (.A1(_3230_),
    .A2(_3262_),
    .A3(_3282_),
    .B1(net72),
    .X(_3309_));
 sky130_fd_sc_hd__xor2_1 _7869_ (.A(_3308_),
    .B(_3309_),
    .X(_3311_));
 sky130_fd_sc_hd__o21bai_2 _7870_ (.A1(net32),
    .A2(_3086_),
    .B1_N(_3201_),
    .Y(_3312_));
 sky130_fd_sc_hd__or2_4 _7871_ (.A(_3288_),
    .B(_3312_),
    .X(_3313_));
 sky130_fd_sc_hd__xnor2_1 _7872_ (.A(_3288_),
    .B(_3312_),
    .Y(_3314_));
 sky130_fd_sc_hd__inv_2 _7873_ (.A(_3314_),
    .Y(_3315_));
 sky130_fd_sc_hd__or4_2 _7874_ (.A(_3232_),
    .B(_3238_),
    .C(_3255_),
    .D(_3290_),
    .X(_3316_));
 sky130_fd_sc_hd__a21o_1 _7875_ (.A1(net222),
    .A2(_3316_),
    .B1(_3315_),
    .X(_3317_));
 sky130_fd_sc_hd__a31o_1 _7876_ (.A1(net222),
    .A2(_3315_),
    .A3(_3316_),
    .B1(net182),
    .X(_3318_));
 sky130_fd_sc_hd__and2b_1 _7877_ (.A_N(_3318_),
    .B(_3317_),
    .X(_3319_));
 sky130_fd_sc_hd__a211o_1 _7878_ (.A1(_2116_),
    .A2(_3311_),
    .B1(_3319_),
    .C1(net241),
    .X(_3320_));
 sky130_fd_sc_hd__nand2_1 _7879_ (.A(\out_reg[10] ),
    .B(_0775_),
    .Y(_3322_));
 sky130_fd_sc_hd__a2bb2o_1 _7880_ (.A1_N(_3304_),
    .A2_N(_3320_),
    .B1(_3322_),
    .B2(net240),
    .X(_3323_));
 sky130_fd_sc_hd__a21oi_1 _7881_ (.A1(_3297_),
    .A2(_3323_),
    .B1(net236),
    .Y(_0031_));
 sky130_fd_sc_hd__a21oi_4 _7882_ (.A1(_1384_),
    .A2(_3095_),
    .B1(_3189_),
    .Y(_3324_));
 sky130_fd_sc_hd__and3_1 _7883_ (.A(_3272_),
    .B(_3298_),
    .C(_3324_),
    .X(_3325_));
 sky130_fd_sc_hd__a21oi_2 _7884_ (.A1(_3272_),
    .A2(_3298_),
    .B1(_3324_),
    .Y(_3326_));
 sky130_fd_sc_hd__nor2_2 _7885_ (.A(_3325_),
    .B(_3326_),
    .Y(_3327_));
 sky130_fd_sc_hd__or3_1 _7886_ (.A(_1472_),
    .B(_3189_),
    .C(_3300_),
    .X(_3328_));
 sky130_fd_sc_hd__or3b_2 _7887_ (.A(_3244_),
    .B(_3302_),
    .C_N(_3328_),
    .X(_3329_));
 sky130_fd_sc_hd__xnor2_2 _7888_ (.A(_3327_),
    .B(_3329_),
    .Y(_3330_));
 sky130_fd_sc_hd__nor2_4 _7889_ (.A(net32),
    .B(_3115_),
    .Y(_3332_));
 sky130_fd_sc_hd__nor2_4 _7890_ (.A(_3313_),
    .B(_3332_),
    .Y(_3333_));
 sky130_fd_sc_hd__a221oi_4 _7891_ (.A1(_2817_),
    .A2(net32),
    .B1(_3313_),
    .B2(_3332_),
    .C1(_3333_),
    .Y(_3334_));
 sky130_fd_sc_hd__a21oi_1 _7892_ (.A1(net222),
    .A2(_3317_),
    .B1(_3334_),
    .Y(_3335_));
 sky130_fd_sc_hd__a311o_1 _7893_ (.A1(net222),
    .A2(_3317_),
    .A3(_3334_),
    .B1(_3335_),
    .C1(net182),
    .X(_3336_));
 sky130_fd_sc_hd__or2_1 _7894_ (.A(net16),
    .B(_3104_),
    .X(_3337_));
 sky130_fd_sc_hd__and3_2 _7895_ (.A(_3280_),
    .B(_3305_),
    .C(_3337_),
    .X(_3338_));
 sky130_fd_sc_hd__inv_2 _7896_ (.A(_3338_),
    .Y(_3339_));
 sky130_fd_sc_hd__o21bai_1 _7897_ (.A1(_3306_),
    .A2(_3337_),
    .B1_N(_3209_),
    .Y(_3340_));
 sky130_fd_sc_hd__nor2_1 _7898_ (.A(_3338_),
    .B(_3340_),
    .Y(_3341_));
 sky130_fd_sc_hd__o21ai_1 _7899_ (.A1(net72),
    .A2(_3308_),
    .B1(_3309_),
    .Y(_3343_));
 sky130_fd_sc_hd__or2_1 _7900_ (.A(_3341_),
    .B(_3343_),
    .X(_3344_));
 sky130_fd_sc_hd__a21oi_1 _7901_ (.A1(_3341_),
    .A2(_3343_),
    .B1(_2117_),
    .Y(_3345_));
 sky130_fd_sc_hd__o2bb2a_1 _7902_ (.A1_N(_3344_),
    .A2_N(_3345_),
    .B1(_1562_),
    .B2(_3330_),
    .X(_3346_));
 sky130_fd_sc_hd__a21oi_2 _7903_ (.A1(_3336_),
    .A2(_3346_),
    .B1(net241),
    .Y(_3347_));
 sky130_fd_sc_hd__a22o_1 _7904_ (.A1(\out_reg[11] ),
    .A2(_0786_),
    .B1(net219),
    .B2(\out_reg[12] ),
    .X(_3348_));
 sky130_fd_sc_hd__o21ba_1 _7905_ (.A1(_3347_),
    .A2(_3348_),
    .B1_N(net236),
    .X(_0032_));
 sky130_fd_sc_hd__o2111a_1 _7906_ (.A1(net15),
    .A2(_3128_),
    .B1(_3272_),
    .C1(_3298_),
    .D1(_3324_),
    .X(_3349_));
 sky130_fd_sc_hd__a311o_1 _7907_ (.A1(_3067_),
    .A2(_3272_),
    .A3(_3324_),
    .B1(_3128_),
    .C1(net15),
    .X(_3350_));
 sky130_fd_sc_hd__or3b_4 _7908_ (.A(_3189_),
    .B(_3349_),
    .C_N(_3350_),
    .X(_3351_));
 sky130_fd_sc_hd__or3_1 _7909_ (.A(net221),
    .B(_3325_),
    .C(_3326_),
    .X(_3353_));
 sky130_fd_sc_hd__and4bb_2 _7910_ (.A_N(_3244_),
    .B_N(_3302_),
    .C(_3328_),
    .D(_3353_),
    .X(_3354_));
 sky130_fd_sc_hd__xnor2_1 _7911_ (.A(_3351_),
    .B(_3354_),
    .Y(_3355_));
 sky130_fd_sc_hd__a21o_2 _7912_ (.A1(_2838_),
    .A2(_3141_),
    .B1(_3201_),
    .X(_3356_));
 sky130_fd_sc_hd__or3_1 _7913_ (.A(_3313_),
    .B(_3332_),
    .C(_3356_),
    .X(_3357_));
 sky130_fd_sc_hd__xor2_2 _7914_ (.A(_3333_),
    .B(_3356_),
    .X(_3358_));
 sky130_fd_sc_hd__o21ai_1 _7915_ (.A1(_3317_),
    .A2(_3334_),
    .B1(net222),
    .Y(_3359_));
 sky130_fd_sc_hd__nand2_1 _7916_ (.A(_3358_),
    .B(_3359_),
    .Y(_3360_));
 sky130_fd_sc_hd__nor2_1 _7917_ (.A(_3358_),
    .B(_3359_),
    .Y(_3361_));
 sky130_fd_sc_hd__or3b_1 _7918_ (.A(_3361_),
    .B(net182),
    .C_N(_3360_),
    .X(_3362_));
 sky130_fd_sc_hd__a21o_1 _7919_ (.A1(_1965_),
    .A2(_3148_),
    .B1(_3209_),
    .X(_3364_));
 sky130_fd_sc_hd__or2_1 _7920_ (.A(_3339_),
    .B(_3364_),
    .X(_3365_));
 sky130_fd_sc_hd__xnor2_1 _7921_ (.A(_3338_),
    .B(_3364_),
    .Y(_3366_));
 sky130_fd_sc_hd__a21o_1 _7922_ (.A1(_2109_),
    .A2(_3344_),
    .B1(_3366_),
    .X(_3367_));
 sky130_fd_sc_hd__nand2_1 _7923_ (.A(_2116_),
    .B(_3367_),
    .Y(_3368_));
 sky130_fd_sc_hd__a31o_1 _7924_ (.A1(_2109_),
    .A2(_3344_),
    .A3(_3366_),
    .B1(_3368_),
    .X(_3369_));
 sky130_fd_sc_hd__o211a_1 _7925_ (.A1(_1562_),
    .A2(_3355_),
    .B1(_3362_),
    .C1(_3369_),
    .X(_3370_));
 sky130_fd_sc_hd__a22o_1 _7926_ (.A1(\out_reg[12] ),
    .A2(_0786_),
    .B1(net219),
    .B2(\out_reg[13] ),
    .X(_3371_));
 sky130_fd_sc_hd__o21ba_1 _7927_ (.A1(net240),
    .A2(_3370_),
    .B1_N(_3371_),
    .X(_3372_));
 sky130_fd_sc_hd__nor2_1 _7928_ (.A(net236),
    .B(_3372_),
    .Y(_0033_));
 sky130_fd_sc_hd__or2_1 _7929_ (.A(net221),
    .B(_3351_),
    .X(_3374_));
 sky130_fd_sc_hd__nor2_1 _7930_ (.A(net15),
    .B(_3349_),
    .Y(_3375_));
 sky130_fd_sc_hd__a21o_1 _7931_ (.A1(_3162_),
    .A2(_3375_),
    .B1(_3189_),
    .X(_3376_));
 sky130_fd_sc_hd__a21oi_1 _7932_ (.A1(_3354_),
    .A2(_3374_),
    .B1(_3376_),
    .Y(_3377_));
 sky130_fd_sc_hd__a31o_1 _7933_ (.A1(_3354_),
    .A2(_3374_),
    .A3(_3376_),
    .B1(_1562_),
    .X(_3378_));
 sky130_fd_sc_hd__or2_2 _7934_ (.A(_3377_),
    .B(_3378_),
    .X(_3379_));
 sky130_fd_sc_hd__nand2_1 _7935_ (.A(_2109_),
    .B(_3367_),
    .Y(_3380_));
 sky130_fd_sc_hd__a21oi_1 _7936_ (.A1(_1930_),
    .A2(_3365_),
    .B1(_3380_),
    .Y(_3381_));
 sky130_fd_sc_hd__a311o_1 _7937_ (.A1(_1930_),
    .A2(_3365_),
    .A3(_3380_),
    .B1(_3381_),
    .C1(_2117_),
    .X(_3382_));
 sky130_fd_sc_hd__a31o_1 _7938_ (.A1(_2838_),
    .A2(_3180_),
    .A3(_3357_),
    .B1(_3201_),
    .X(_3383_));
 sky130_fd_sc_hd__nand2_1 _7939_ (.A(net222),
    .B(_3360_),
    .Y(_3385_));
 sky130_fd_sc_hd__xnor2_1 _7940_ (.A(_3383_),
    .B(_3385_),
    .Y(_3386_));
 sky130_fd_sc_hd__o21ba_1 _7941_ (.A1(net182),
    .A2(_3386_),
    .B1_N(net241),
    .X(_3387_));
 sky130_fd_sc_hd__nand2_1 _7942_ (.A(\out_reg[13] ),
    .B(net228),
    .Y(_3388_));
 sky130_fd_sc_hd__a32o_1 _7943_ (.A1(_3379_),
    .A2(_3382_),
    .A3(_3387_),
    .B1(_3388_),
    .B2(net242),
    .X(_3389_));
 sky130_fd_sc_hd__nand2_1 _7944_ (.A(\out_reg[14] ),
    .B(net220),
    .Y(_3390_));
 sky130_fd_sc_hd__a21oi_1 _7945_ (.A1(_3389_),
    .A2(_3390_),
    .B1(net237),
    .Y(_0034_));
 sky130_fd_sc_hd__o21ai_1 _7946_ (.A1(net72),
    .A2(_2115_),
    .B1(_2114_),
    .Y(_3391_));
 sky130_fd_sc_hd__or3_1 _7947_ (.A(\cmd[7] ),
    .B(\cmd[6] ),
    .C(_3391_),
    .X(_3392_));
 sky130_fd_sc_hd__nand2_1 _7948_ (.A(\cmd[7] ),
    .B(\cmd[6] ),
    .Y(_3393_));
 sky130_fd_sc_hd__nand2_1 _7949_ (.A(_0668_),
    .B(net212),
    .Y(_3395_));
 sky130_fd_sc_hd__a22oi_2 _7950_ (.A1(\cmd[6] ),
    .A2(_2113_),
    .B1(_3395_),
    .B2(\cmd[7] ),
    .Y(_3396_));
 sky130_fd_sc_hd__a221o_1 _7951_ (.A1(net234),
    .A2(net201),
    .B1(_1215_),
    .B2(net222),
    .C1(_3396_),
    .X(_3397_));
 sky130_fd_sc_hd__a31o_1 _7952_ (.A1(_3392_),
    .A2(_3393_),
    .A3(_3397_),
    .B1(net242),
    .X(_3398_));
 sky130_fd_sc_hd__o22a_1 _7953_ (.A1(\out_reg[14] ),
    .A2(_0797_),
    .B1(_2985_),
    .B2(\out_reg[15] ),
    .X(_3399_));
 sky130_fd_sc_hd__and3b_1 _7954_ (.A_N(net238),
    .B(_3398_),
    .C(_3399_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _7955_ (.A0(\out_reg[15] ),
    .A1(net5),
    .S(net217),
    .X(_0036_));
 sky130_fd_sc_hd__or4b_2 _7956_ (.A(\counter[3] ),
    .B(_0635_),
    .C(_0701_),
    .D_N(\counter[4] ),
    .X(_3400_));
 sky130_fd_sc_hd__inv_2 _7957_ (.A(_3400_),
    .Y(_3401_));
 sky130_fd_sc_hd__or3b_2 _7958_ (.A(net238),
    .B(_3401_),
    .C_N(net240),
    .X(_3402_));
 sky130_fd_sc_hd__a21oi_1 _7959_ (.A1(\in_reg[1] ),
    .A2(_0712_),
    .B1(mode),
    .Y(_3404_));
 sky130_fd_sc_hd__nor2_1 _7960_ (.A(_3402_),
    .B(_3404_),
    .Y(_0037_));
 sky130_fd_sc_hd__nor2_1 _7961_ (.A(_0712_),
    .B(_3402_),
    .Y(_3405_));
 sky130_fd_sc_hd__o21ai_1 _7962_ (.A1(\counter[0] ),
    .A2(net228),
    .B1(_3405_),
    .Y(_3406_));
 sky130_fd_sc_hd__a21oi_1 _7963_ (.A1(\counter[0] ),
    .A2(net228),
    .B1(_3406_),
    .Y(_0038_));
 sky130_fd_sc_hd__and3_2 _7964_ (.A(\counter[1] ),
    .B(\counter[0] ),
    .C(net228),
    .X(_3407_));
 sky130_fd_sc_hd__a21o_1 _7965_ (.A1(\counter[0] ),
    .A2(net228),
    .B1(\counter[1] ),
    .X(_3408_));
 sky130_fd_sc_hd__and3b_1 _7966_ (.A_N(_3407_),
    .B(_3408_),
    .C(_3405_),
    .X(_0039_));
 sky130_fd_sc_hd__o21ai_1 _7967_ (.A1(\counter[2] ),
    .A2(_3407_),
    .B1(_3405_),
    .Y(_3409_));
 sky130_fd_sc_hd__a21oi_1 _7968_ (.A1(\counter[2] ),
    .A2(_3407_),
    .B1(_3409_),
    .Y(_0040_));
 sky130_fd_sc_hd__a21o_1 _7969_ (.A1(\counter[2] ),
    .A2(_3407_),
    .B1(\counter[3] ),
    .X(_3411_));
 sky130_fd_sc_hd__and3_1 _7970_ (.A(\counter[3] ),
    .B(\counter[2] ),
    .C(_3407_),
    .X(_3412_));
 sky130_fd_sc_hd__and3b_1 _7971_ (.A_N(_3412_),
    .B(_3405_),
    .C(_3411_),
    .X(_0041_));
 sky130_fd_sc_hd__a211o_1 _7972_ (.A1(\counter[4] ),
    .A2(_3412_),
    .B1(_3402_),
    .C1(_0712_),
    .X(_3413_));
 sky130_fd_sc_hd__o21ba_1 _7973_ (.A1(\counter[4] ),
    .A2(_3412_),
    .B1_N(_3413_),
    .X(_0042_));
 sky130_fd_sc_hd__or4b_1 _7974_ (.A(net238),
    .B(\cmd[0] ),
    .C(_3400_),
    .D_N(net240),
    .X(_3414_));
 sky130_fd_sc_hd__mux2_1 _7975_ (.A0(\in_reg[0] ),
    .A1(net235),
    .S(net208),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _7976_ (.A0(\in_reg[1] ),
    .A1(\posit_add.in1[1] ),
    .S(net208),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _7977_ (.A0(\in_reg[2] ),
    .A1(\posit_add.in1[2] ),
    .S(net209),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _7978_ (.A0(\in_reg[3] ),
    .A1(\posit_add.in1[3] ),
    .S(net208),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _7979_ (.A0(\in_reg[4] ),
    .A1(\posit_add.in1[4] ),
    .S(net208),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _7980_ (.A0(\in_reg[5] ),
    .A1(\posit_add.in1[5] ),
    .S(net209),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _7981_ (.A0(\in_reg[6] ),
    .A1(\posit_add.in1[6] ),
    .S(net209),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _7982_ (.A0(\in_reg[7] ),
    .A1(\posit_add.in1[7] ),
    .S(net208),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _7983_ (.A0(\in_reg[8] ),
    .A1(\posit_add.in1[8] ),
    .S(net208),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _7984_ (.A0(\in_reg[9] ),
    .A1(\posit_add.in1[9] ),
    .S(net208),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _7985_ (.A0(\in_reg[10] ),
    .A1(\posit_add.in1[10] ),
    .S(net208),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _7986_ (.A0(\in_reg[11] ),
    .A1(\posit_add.in1[11] ),
    .S(net208),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _7987_ (.A0(\in_reg[12] ),
    .A1(\posit_add.in1[12] ),
    .S(net208),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _7988_ (.A0(\in_reg[13] ),
    .A1(\posit_add.in1[13] ),
    .S(net209),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _7989_ (.A0(\in_reg[14] ),
    .A1(\posit_add.in1[14] ),
    .S(net209),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _7990_ (.A0(\in_reg[15] ),
    .A1(net233),
    .S(net209),
    .X(_0058_));
 sky130_fd_sc_hd__and4b_1 _7991_ (.A_N(net238),
    .B(\cmd[0] ),
    .C(_3401_),
    .D(net240),
    .X(_3417_));
 sky130_fd_sc_hd__mux2_1 _7992_ (.A0(\posit_add.in2[0] ),
    .A1(\in_reg[0] ),
    .S(net206),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _7993_ (.A0(\posit_add.in2[1] ),
    .A1(\in_reg[1] ),
    .S(net206),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _7994_ (.A0(\posit_add.in2[2] ),
    .A1(\in_reg[2] ),
    .S(net206),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _7995_ (.A0(\posit_add.in2[3] ),
    .A1(\in_reg[3] ),
    .S(net206),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _7996_ (.A0(\posit_add.in2[4] ),
    .A1(\in_reg[4] ),
    .S(net207),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _7997_ (.A0(\posit_add.in2[5] ),
    .A1(\in_reg[5] ),
    .S(net207),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _7998_ (.A0(\posit_add.in2[6] ),
    .A1(\in_reg[6] ),
    .S(net206),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _7999_ (.A0(\posit_add.in2[7] ),
    .A1(\in_reg[7] ),
    .S(net206),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _8000_ (.A0(\posit_add.in2[8] ),
    .A1(\in_reg[8] ),
    .S(net206),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _8001_ (.A0(\posit_add.in2[9] ),
    .A1(\in_reg[9] ),
    .S(net206),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _8002_ (.A0(\posit_add.in2[10] ),
    .A1(\in_reg[10] ),
    .S(net206),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _8003_ (.A0(\posit_add.in2[11] ),
    .A1(\in_reg[11] ),
    .S(net206),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _8004_ (.A0(\posit_add.in2[12] ),
    .A1(\in_reg[12] ),
    .S(net207),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _8005_ (.A0(\posit_add.in2[13] ),
    .A1(\in_reg[13] ),
    .S(net207),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _8006_ (.A0(\posit_add.in2[14] ),
    .A1(\in_reg[14] ),
    .S(net207),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _8007_ (.A0(net231),
    .A1(\in_reg[15] ),
    .S(net207),
    .X(_0074_));
 sky130_fd_sc_hd__dfxtp_1 _8008_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0000_),
    .Q(\cmd[0] ));
 sky130_fd_sc_hd__dfxtp_4 _8009_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0001_),
    .Q(\cmd[6] ));
 sky130_fd_sc_hd__dfxtp_4 _8010_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0002_),
    .Q(\cmd[7] ));
 sky130_fd_sc_hd__dfxtp_2 _8011_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0003_),
    .Q(\in_reg[0] ));
 sky130_fd_sc_hd__dfxtp_2 _8012_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0004_),
    .Q(\in_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8013_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0005_),
    .Q(\in_reg[2] ));
 sky130_fd_sc_hd__dfxtp_2 _8014_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0006_),
    .Q(\in_reg[3] ));
 sky130_fd_sc_hd__dfxtp_2 _8015_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0007_),
    .Q(\in_reg[4] ));
 sky130_fd_sc_hd__dfxtp_2 _8016_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0008_),
    .Q(\in_reg[5] ));
 sky130_fd_sc_hd__dfxtp_2 _8017_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0009_),
    .Q(\in_reg[6] ));
 sky130_fd_sc_hd__dfxtp_2 _8018_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0010_),
    .Q(\in_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8019_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0011_),
    .Q(\in_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8020_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0012_),
    .Q(\in_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8021_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0013_),
    .Q(\in_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8022_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0014_),
    .Q(\in_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8023_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0015_),
    .Q(\in_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8024_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0016_),
    .Q(\in_reg[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8025_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0017_),
    .Q(\in_reg[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8026_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0018_),
    .Q(\in_reg[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8027_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0019_),
    .Q(last_SCLK));
 sky130_fd_sc_hd__dfxtp_1 _8028_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0020_),
    .Q(\out_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8029_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0021_),
    .Q(\out_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8030_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0022_),
    .Q(\out_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8031_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0023_),
    .Q(\out_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8032_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0024_),
    .Q(\out_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8033_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0025_),
    .Q(\out_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8034_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0026_),
    .Q(\out_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8035_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0027_),
    .Q(\out_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8036_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0028_),
    .Q(\out_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8037_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0029_),
    .Q(\out_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8038_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0030_),
    .Q(\out_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8039_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0031_),
    .Q(\out_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8040_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0032_),
    .Q(\out_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8041_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0033_),
    .Q(\out_reg[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8042_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0034_),
    .Q(\out_reg[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8043_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0035_),
    .Q(\out_reg[15] ));
 sky130_fd_sc_hd__dfxtp_4 _8044_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0036_),
    .Q(net5));
 sky130_fd_sc_hd__dfxtp_2 _8045_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0037_),
    .Q(mode));
 sky130_fd_sc_hd__dfxtp_1 _8046_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0038_),
    .Q(\counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8047_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0039_),
    .Q(\counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8048_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0040_),
    .Q(\counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8049_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0041_),
    .Q(\counter[3] ));
 sky130_fd_sc_hd__dfxtp_2 _8050_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0042_),
    .Q(\counter[4] ));
 sky130_fd_sc_hd__dfxtp_4 _8051_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0043_),
    .Q(\posit_add.in1[0] ));
 sky130_fd_sc_hd__dfxtp_4 _8052_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0044_),
    .Q(\posit_add.in1[1] ));
 sky130_fd_sc_hd__dfxtp_4 _8053_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0045_),
    .Q(\posit_add.in1[2] ));
 sky130_fd_sc_hd__dfxtp_4 _8054_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0046_),
    .Q(\posit_add.in1[3] ));
 sky130_fd_sc_hd__dfxtp_4 _8055_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0047_),
    .Q(\posit_add.in1[4] ));
 sky130_fd_sc_hd__dfxtp_4 _8056_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0048_),
    .Q(\posit_add.in1[5] ));
 sky130_fd_sc_hd__dfxtp_4 _8057_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0049_),
    .Q(\posit_add.in1[6] ));
 sky130_fd_sc_hd__dfxtp_4 _8058_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0050_),
    .Q(\posit_add.in1[7] ));
 sky130_fd_sc_hd__dfxtp_4 _8059_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0051_),
    .Q(\posit_add.in1[8] ));
 sky130_fd_sc_hd__dfxtp_4 _8060_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0052_),
    .Q(\posit_add.in1[9] ));
 sky130_fd_sc_hd__dfxtp_4 _8061_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0053_),
    .Q(\posit_add.in1[10] ));
 sky130_fd_sc_hd__dfxtp_4 _8062_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0054_),
    .Q(\posit_add.in1[11] ));
 sky130_fd_sc_hd__dfxtp_4 _8063_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0055_),
    .Q(\posit_add.in1[12] ));
 sky130_fd_sc_hd__dfxtp_4 _8064_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0056_),
    .Q(\posit_add.in1[13] ));
 sky130_fd_sc_hd__dfxtp_2 _8065_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0057_),
    .Q(\posit_add.in1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8066_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0058_),
    .Q(\posit_add.in1[15] ));
 sky130_fd_sc_hd__dfxtp_4 _8067_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0059_),
    .Q(\posit_add.in2[0] ));
 sky130_fd_sc_hd__dfxtp_4 _8068_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0060_),
    .Q(\posit_add.in2[1] ));
 sky130_fd_sc_hd__dfxtp_4 _8069_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0061_),
    .Q(\posit_add.in2[2] ));
 sky130_fd_sc_hd__dfxtp_4 _8070_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0062_),
    .Q(\posit_add.in2[3] ));
 sky130_fd_sc_hd__dfxtp_4 _8071_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0063_),
    .Q(\posit_add.in2[4] ));
 sky130_fd_sc_hd__dfxtp_4 _8072_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0064_),
    .Q(\posit_add.in2[5] ));
 sky130_fd_sc_hd__dfxtp_4 _8073_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0065_),
    .Q(\posit_add.in2[6] ));
 sky130_fd_sc_hd__dfxtp_2 _8074_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0066_),
    .Q(\posit_add.in2[7] ));
 sky130_fd_sc_hd__dfxtp_4 _8075_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0067_),
    .Q(\posit_add.in2[8] ));
 sky130_fd_sc_hd__dfxtp_4 _8076_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0068_),
    .Q(\posit_add.in2[9] ));
 sky130_fd_sc_hd__dfxtp_4 _8077_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0069_),
    .Q(\posit_add.in2[10] ));
 sky130_fd_sc_hd__dfxtp_4 _8078_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0070_),
    .Q(\posit_add.in2[11] ));
 sky130_fd_sc_hd__dfxtp_4 _8079_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0071_),
    .Q(\posit_add.in2[12] ));
 sky130_fd_sc_hd__dfxtp_4 _8080_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0072_),
    .Q(\posit_add.in2[13] ));
 sky130_fd_sc_hd__dfxtp_4 _8081_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0073_),
    .Q(\posit_add.in2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8082_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0074_),
    .Q(\posit_add.in2[15] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__buf_4 fanout10 (.A(_1390_),
    .X(net10));
 sky130_fd_sc_hd__buf_8 fanout100 (.A(_1587_),
    .X(net100));
 sky130_fd_sc_hd__buf_6 fanout101 (.A(_1232_),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_16 fanout102 (.A(net105),
    .X(net102));
 sky130_fd_sc_hd__buf_4 fanout103 (.A(net105),
    .X(net103));
 sky130_fd_sc_hd__buf_6 fanout104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_16 fanout105 (.A(_0588_),
    .X(net105));
 sky130_fd_sc_hd__buf_8 fanout106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__buf_6 fanout107 (.A(net109),
    .X(net107));
 sky130_fd_sc_hd__buf_6 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_16 fanout109 (.A(_0549_),
    .X(net109));
 sky130_fd_sc_hd__buf_4 fanout11 (.A(_1389_),
    .X(net11));
 sky130_fd_sc_hd__buf_12 fanout110 (.A(_0542_),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_16 fanout111 (.A(_0542_),
    .X(net111));
 sky130_fd_sc_hd__buf_6 fanout112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__buf_8 fanout113 (.A(_0541_),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_16 fanout114 (.A(_3589_),
    .X(net114));
 sky130_fd_sc_hd__buf_8 fanout115 (.A(_3538_),
    .X(net115));
 sky130_fd_sc_hd__buf_6 fanout116 (.A(_3538_),
    .X(net116));
 sky130_fd_sc_hd__buf_8 fanout117 (.A(net119),
    .X(net117));
 sky130_fd_sc_hd__buf_4 fanout118 (.A(net119),
    .X(net118));
 sky130_fd_sc_hd__buf_4 fanout119 (.A(_3522_),
    .X(net119));
 sky130_fd_sc_hd__buf_4 fanout12 (.A(_1389_),
    .X(net12));
 sky130_fd_sc_hd__buf_8 fanout120 (.A(_3505_),
    .X(net120));
 sky130_fd_sc_hd__buf_4 fanout121 (.A(_3505_),
    .X(net121));
 sky130_fd_sc_hd__buf_8 fanout122 (.A(net123),
    .X(net122));
 sky130_fd_sc_hd__buf_12 fanout123 (.A(_3511_),
    .X(net123));
 sky130_fd_sc_hd__buf_8 fanout124 (.A(_3510_),
    .X(net124));
 sky130_fd_sc_hd__buf_6 fanout125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__buf_4 fanout126 (.A(net127),
    .X(net126));
 sky130_fd_sc_hd__buf_8 fanout127 (.A(_3476_),
    .X(net127));
 sky130_fd_sc_hd__buf_8 fanout128 (.A(_3475_),
    .X(net128));
 sky130_fd_sc_hd__buf_4 fanout129 (.A(_1902_),
    .X(net129));
 sky130_fd_sc_hd__buf_4 fanout13 (.A(_1388_),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 fanout130 (.A(_1902_),
    .X(net130));
 sky130_fd_sc_hd__buf_4 fanout131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(_1792_),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_8 fanout133 (.A(_1781_),
    .X(net133));
 sky130_fd_sc_hd__buf_6 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__buf_12 fanout135 (.A(_3509_),
    .X(net135));
 sky130_fd_sc_hd__buf_6 fanout136 (.A(net137),
    .X(net136));
 sky130_fd_sc_hd__buf_8 fanout137 (.A(_3508_),
    .X(net137));
 sky130_fd_sc_hd__buf_4 fanout138 (.A(_3499_),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_16 fanout139 (.A(_3499_),
    .X(net139));
 sky130_fd_sc_hd__buf_12 fanout14 (.A(net15),
    .X(net14));
 sky130_fd_sc_hd__buf_12 fanout140 (.A(_3498_),
    .X(net140));
 sky130_fd_sc_hd__buf_4 fanout141 (.A(net143),
    .X(net141));
 sky130_fd_sc_hd__buf_4 fanout142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__buf_8 fanout143 (.A(net144),
    .X(net143));
 sky130_fd_sc_hd__buf_6 fanout144 (.A(_3495_),
    .X(net144));
 sky130_fd_sc_hd__buf_6 fanout145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__buf_8 fanout146 (.A(_3494_),
    .X(net146));
 sky130_fd_sc_hd__buf_6 fanout147 (.A(net148),
    .X(net147));
 sky130_fd_sc_hd__buf_8 fanout148 (.A(net149),
    .X(net148));
 sky130_fd_sc_hd__buf_6 fanout149 (.A(_3489_),
    .X(net149));
 sky130_fd_sc_hd__buf_6 fanout15 (.A(_1383_),
    .X(net15));
 sky130_fd_sc_hd__buf_6 fanout150 (.A(net152),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_4 fanout151 (.A(net152),
    .X(net151));
 sky130_fd_sc_hd__buf_4 fanout152 (.A(net153),
    .X(net152));
 sky130_fd_sc_hd__buf_4 fanout153 (.A(net154),
    .X(net153));
 sky130_fd_sc_hd__buf_8 fanout154 (.A(_3488_),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_8 fanout155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_8 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__buf_6 fanout157 (.A(_3485_),
    .X(net157));
 sky130_fd_sc_hd__buf_4 fanout158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__buf_6 fanout159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__buf_4 fanout16 (.A(_1964_),
    .X(net16));
 sky130_fd_sc_hd__buf_8 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_16 fanout161 (.A(_3484_),
    .X(net161));
 sky130_fd_sc_hd__buf_8 fanout162 (.A(_3481_),
    .X(net162));
 sky130_fd_sc_hd__buf_4 fanout163 (.A(_3481_),
    .X(net163));
 sky130_fd_sc_hd__buf_6 fanout164 (.A(net166),
    .X(net164));
 sky130_fd_sc_hd__buf_6 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__buf_12 fanout166 (.A(_3480_),
    .X(net166));
 sky130_fd_sc_hd__buf_8 fanout167 (.A(net169),
    .X(net167));
 sky130_fd_sc_hd__buf_4 fanout168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__buf_6 fanout169 (.A(_1726_),
    .X(net169));
 sky130_fd_sc_hd__buf_2 fanout17 (.A(_1964_),
    .X(net17));
 sky130_fd_sc_hd__buf_6 fanout170 (.A(net171),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_16 fanout171 (.A(_1462_),
    .X(net171));
 sky130_fd_sc_hd__buf_12 fanout172 (.A(_1451_),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 fanout173 (.A(_1451_),
    .X(net173));
 sky130_fd_sc_hd__buf_12 fanout174 (.A(net176),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_4 fanout175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__buf_8 fanout176 (.A(_3703_),
    .X(net176));
 sky130_fd_sc_hd__buf_8 fanout177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__buf_8 fanout178 (.A(_3497_),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_4 fanout179 (.A(_3497_),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_8 fanout18 (.A(net19),
    .X(net18));
 sky130_fd_sc_hd__buf_8 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__buf_6 fanout181 (.A(_3496_),
    .X(net181));
 sky130_fd_sc_hd__buf_4 fanout182 (.A(_2979_),
    .X(net182));
 sky130_fd_sc_hd__buf_2 fanout183 (.A(_2979_),
    .X(net183));
 sky130_fd_sc_hd__buf_6 fanout184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__buf_4 fanout185 (.A(_3215_),
    .X(net185));
 sky130_fd_sc_hd__buf_12 fanout186 (.A(net187),
    .X(net186));
 sky130_fd_sc_hd__buf_6 fanout187 (.A(_3204_),
    .X(net187));
 sky130_fd_sc_hd__buf_4 fanout188 (.A(net189),
    .X(net188));
 sky130_fd_sc_hd__buf_6 fanout189 (.A(_3140_),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_4 fanout19 (.A(_1958_),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_16 fanout190 (.A(_3129_),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_8 fanout191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__buf_6 fanout192 (.A(_2990_),
    .X(net192));
 sky130_fd_sc_hd__buf_6 fanout193 (.A(_2980_),
    .X(net193));
 sky130_fd_sc_hd__buf_8 fanout194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__buf_2 fanout195 (.A(_2859_),
    .X(net195));
 sky130_fd_sc_hd__buf_6 fanout196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__buf_4 fanout197 (.A(net198),
    .X(net197));
 sky130_fd_sc_hd__buf_2 fanout198 (.A(_2848_),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_16 fanout199 (.A(_0333_),
    .X(net199));
 sky130_fd_sc_hd__buf_4 fanout20 (.A(net21),
    .X(net20));
 sky130_fd_sc_hd__buf_8 fanout200 (.A(net202),
    .X(net200));
 sky130_fd_sc_hd__buf_12 fanout201 (.A(net202),
    .X(net201));
 sky130_fd_sc_hd__buf_12 fanout202 (.A(_0332_),
    .X(net202));
 sky130_fd_sc_hd__buf_12 fanout203 (.A(net205),
    .X(net203));
 sky130_fd_sc_hd__buf_12 fanout204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__buf_6 fanout205 (.A(_1077_),
    .X(net205));
 sky130_fd_sc_hd__buf_6 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__buf_4 fanout207 (.A(_3417_),
    .X(net207));
 sky130_fd_sc_hd__buf_6 fanout208 (.A(net209),
    .X(net208));
 sky130_fd_sc_hd__buf_4 fanout209 (.A(_3414_),
    .X(net209));
 sky130_fd_sc_hd__buf_2 fanout21 (.A(net22),
    .X(net21));
 sky130_fd_sc_hd__buf_8 fanout210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__buf_12 fanout211 (.A(_3507_),
    .X(net211));
 sky130_fd_sc_hd__buf_12 fanout212 (.A(_3507_),
    .X(net212));
 sky130_fd_sc_hd__buf_4 fanout213 (.A(_3507_),
    .X(net213));
 sky130_fd_sc_hd__buf_6 fanout214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__buf_12 fanout215 (.A(net216),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_16 fanout216 (.A(_2210_),
    .X(net216));
 sky130_fd_sc_hd__buf_6 fanout217 (.A(_0808_),
    .X(net217));
 sky130_fd_sc_hd__buf_4 fanout218 (.A(_0808_),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_4 fanout219 (.A(_2984_),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_4 fanout22 (.A(_1937_),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout220 (.A(_2984_),
    .X(net220));
 sky130_fd_sc_hd__buf_4 fanout221 (.A(_1472_),
    .X(net221));
 sky130_fd_sc_hd__buf_4 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__buf_4 fanout223 (.A(_1471_),
    .X(net223));
 sky130_fd_sc_hd__buf_8 fanout224 (.A(net225),
    .X(net224));
 sky130_fd_sc_hd__buf_4 fanout225 (.A(net226),
    .X(net225));
 sky130_fd_sc_hd__buf_8 fanout226 (.A(_1471_),
    .X(net226));
 sky130_fd_sc_hd__buf_6 fanout227 (.A(_2122_),
    .X(net227));
 sky130_fd_sc_hd__buf_4 fanout228 (.A(_0775_),
    .X(net228));
 sky130_fd_sc_hd__buf_8 fanout229 (.A(net230),
    .X(net229));
 sky130_fd_sc_hd__buf_4 fanout23 (.A(net24),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 fanout230 (.A(net231),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_16 fanout231 (.A(\posit_add.in2[15] ),
    .X(net231));
 sky130_fd_sc_hd__buf_6 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__buf_6 fanout233 (.A(net234),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_16 fanout234 (.A(\posit_add.in1[15] ),
    .X(net234));
 sky130_fd_sc_hd__buf_6 fanout235 (.A(\posit_add.in1[0] ),
    .X(net235));
 sky130_fd_sc_hd__buf_4 fanout236 (.A(net238),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_2 fanout237 (.A(net238),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_4 fanout238 (.A(net4),
    .X(net238));
 sky130_fd_sc_hd__buf_4 fanout239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__buf_4 fanout24 (.A(_1951_),
    .X(net24));
 sky130_fd_sc_hd__buf_4 fanout240 (.A(net242),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_8 fanout241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__buf_4 fanout242 (.A(net1),
    .X(net242));
 sky130_fd_sc_hd__buf_4 fanout25 (.A(net26),
    .X(net25));
 sky130_fd_sc_hd__buf_2 fanout26 (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__buf_4 fanout27 (.A(_2847_),
    .X(net27));
 sky130_fd_sc_hd__buf_4 fanout28 (.A(net29),
    .X(net28));
 sky130_fd_sc_hd__buf_6 fanout29 (.A(_2846_),
    .X(net29));
 sky130_fd_sc_hd__buf_6 fanout30 (.A(net31),
    .X(net30));
 sky130_fd_sc_hd__buf_6 fanout31 (.A(_2842_),
    .X(net31));
 sky130_fd_sc_hd__buf_6 fanout32 (.A(net33),
    .X(net32));
 sky130_fd_sc_hd__buf_4 fanout33 (.A(_2839_),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_8 fanout34 (.A(net35),
    .X(net34));
 sky130_fd_sc_hd__buf_4 fanout35 (.A(_1912_),
    .X(net35));
 sky130_fd_sc_hd__buf_4 fanout36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 fanout37 (.A(_1897_),
    .X(net37));
 sky130_fd_sc_hd__buf_4 fanout38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__buf_4 fanout39 (.A(_1884_),
    .X(net39));
 sky130_fd_sc_hd__buf_6 fanout40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__buf_4 fanout41 (.A(_2799_),
    .X(net41));
 sky130_fd_sc_hd__buf_8 fanout42 (.A(_0349_),
    .X(net42));
 sky130_fd_sc_hd__buf_12 fanout43 (.A(_0326_),
    .X(net43));
 sky130_fd_sc_hd__buf_4 fanout44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 fanout45 (.A(_1784_),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_16 fanout46 (.A(_0410_),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_16 fanout47 (.A(_0289_),
    .X(net47));
 sky130_fd_sc_hd__buf_8 fanout48 (.A(_0474_),
    .X(net48));
 sky130_fd_sc_hd__buf_8 fanout49 (.A(_0605_),
    .X(net49));
 sky130_fd_sc_hd__buf_4 fanout50 (.A(net52),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 fanout51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__buf_6 fanout52 (.A(_0590_),
    .X(net52));
 sky130_fd_sc_hd__buf_8 fanout53 (.A(_0516_),
    .X(net53));
 sky130_fd_sc_hd__buf_8 fanout54 (.A(_0526_),
    .X(net54));
 sky130_fd_sc_hd__buf_6 fanout55 (.A(_0123_),
    .X(net55));
 sky130_fd_sc_hd__buf_6 fanout56 (.A(_0099_),
    .X(net56));
 sky130_fd_sc_hd__buf_4 fanout57 (.A(_0075_),
    .X(net57));
 sky130_fd_sc_hd__buf_4 fanout58 (.A(_3893_),
    .X(net58));
 sky130_fd_sc_hd__buf_8 fanout59 (.A(_3893_),
    .X(net59));
 sky130_fd_sc_hd__buf_6 fanout6 (.A(net8),
    .X(net6));
 sky130_fd_sc_hd__buf_8 fanout60 (.A(_3997_),
    .X(net60));
 sky130_fd_sc_hd__buf_6 fanout61 (.A(_1657_),
    .X(net61));
 sky130_fd_sc_hd__buf_4 fanout62 (.A(_1653_),
    .X(net62));
 sky130_fd_sc_hd__buf_4 fanout63 (.A(_1647_),
    .X(net63));
 sky130_fd_sc_hd__buf_12 fanout64 (.A(_0296_),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_8 fanout65 (.A(_0296_),
    .X(net65));
 sky130_fd_sc_hd__buf_12 fanout66 (.A(net67),
    .X(net66));
 sky130_fd_sc_hd__buf_12 fanout67 (.A(_0295_),
    .X(net67));
 sky130_fd_sc_hd__buf_6 fanout68 (.A(_3646_),
    .X(net68));
 sky130_fd_sc_hd__buf_6 fanout69 (.A(net70),
    .X(net69));
 sky130_fd_sc_hd__buf_2 fanout7 (.A(net8),
    .X(net7));
 sky130_fd_sc_hd__buf_12 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__buf_6 fanout71 (.A(_3463_),
    .X(net71));
 sky130_fd_sc_hd__buf_4 fanout72 (.A(_2108_),
    .X(net72));
 sky130_fd_sc_hd__buf_12 fanout73 (.A(_0548_),
    .X(net73));
 sky130_fd_sc_hd__buf_8 fanout74 (.A(net75),
    .X(net74));
 sky130_fd_sc_hd__buf_12 fanout75 (.A(_0498_),
    .X(net75));
 sky130_fd_sc_hd__buf_8 fanout76 (.A(net77),
    .X(net76));
 sky130_fd_sc_hd__buf_12 fanout77 (.A(_0497_),
    .X(net77));
 sky130_fd_sc_hd__buf_6 fanout78 (.A(_0431_),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_16 fanout79 (.A(_0431_),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_4 fanout8 (.A(_1413_),
    .X(net8));
 sky130_fd_sc_hd__buf_12 fanout80 (.A(_0430_),
    .X(net80));
 sky130_fd_sc_hd__buf_12 fanout81 (.A(net82),
    .X(net81));
 sky130_fd_sc_hd__buf_12 fanout82 (.A(_0373_),
    .X(net82));
 sky130_fd_sc_hd__buf_12 fanout83 (.A(_0372_),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_16 fanout84 (.A(_0363_),
    .X(net84));
 sky130_fd_sc_hd__buf_12 fanout85 (.A(_0363_),
    .X(net85));
 sky130_fd_sc_hd__buf_6 fanout86 (.A(_0363_),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_16 fanout87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_16 fanout88 (.A(_0315_),
    .X(net88));
 sky130_fd_sc_hd__buf_8 fanout89 (.A(net91),
    .X(net89));
 sky130_fd_sc_hd__buf_4 fanout9 (.A(_1390_),
    .X(net9));
 sky130_fd_sc_hd__buf_2 fanout90 (.A(net91),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_8 fanout91 (.A(_0314_),
    .X(net91));
 sky130_fd_sc_hd__buf_6 fanout92 (.A(_3602_),
    .X(net92));
 sky130_fd_sc_hd__buf_8 fanout93 (.A(_3601_),
    .X(net93));
 sky130_fd_sc_hd__buf_4 fanout94 (.A(_3601_),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_8 fanout95 (.A(_3581_),
    .X(net95));
 sky130_fd_sc_hd__buf_4 fanout96 (.A(_3581_),
    .X(net96));
 sky130_fd_sc_hd__buf_8 fanout97 (.A(_1587_),
    .X(net97));
 sky130_fd_sc_hd__buf_6 fanout98 (.A(_1587_),
    .X(net98));
 sky130_fd_sc_hd__buf_6 fanout99 (.A(_1587_),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(io_in[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input2 (.A(io_in[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(io_in[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(rst),
    .X(net4));
 sky130_fd_sc_hd__buf_4 output5 (.A(net5),
    .X(io_out[3]));
 sky130_fd_sc_hd__conb_1 posit_unit_243 (.LO(net243));
 sky130_fd_sc_hd__conb_1 posit_unit_244 (.LO(net244));
 sky130_fd_sc_hd__conb_1 posit_unit_245 (.LO(net245));
 assign io_out[0] = net243;
 assign io_out[1] = net244;
 assign io_out[2] = net245;
endmodule

