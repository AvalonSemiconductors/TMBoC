// This is the unpowered netlist.
module wrapped_6502 (clk,
    io_oeb,
    rst,
    io_in,
    io_out);
 input clk;
 output io_oeb;
 input rst;
 input [9:0] io_in;
 output [26:0] io_out;

 wire net90;
 wire net91;
 wire \MOS6502.ABH[0] ;
 wire \MOS6502.ABH[1] ;
 wire \MOS6502.ABH[2] ;
 wire \MOS6502.ABH[3] ;
 wire \MOS6502.ABH[4] ;
 wire \MOS6502.ABH[5] ;
 wire \MOS6502.ABH[6] ;
 wire \MOS6502.ABH[7] ;
 wire \MOS6502.ABL[0] ;
 wire \MOS6502.ABL[1] ;
 wire \MOS6502.ABL[2] ;
 wire \MOS6502.ABL[3] ;
 wire \MOS6502.ABL[4] ;
 wire \MOS6502.ABL[5] ;
 wire \MOS6502.ABL[6] ;
 wire \MOS6502.ABL[7] ;
 wire \MOS6502.ADD[0] ;
 wire \MOS6502.ADD[1] ;
 wire \MOS6502.ADD[2] ;
 wire \MOS6502.ADD[3] ;
 wire \MOS6502.ADD[4] ;
 wire \MOS6502.ADD[5] ;
 wire \MOS6502.ADD[6] ;
 wire \MOS6502.ADD[7] ;
 wire \MOS6502.AI[7] ;
 wire \MOS6502.ALU.AI7 ;
 wire \MOS6502.ALU.BI7 ;
 wire \MOS6502.ALU.CO ;
 wire \MOS6502.ALU.HC ;
 wire \MOS6502.ALU.temp[0] ;
 wire \MOS6502.ALU.temp[1] ;
 wire \MOS6502.ALU.temp[2] ;
 wire \MOS6502.ALU.temp[3] ;
 wire \MOS6502.ALU.temp[4] ;
 wire \MOS6502.ALU.temp[5] ;
 wire \MOS6502.ALU.temp[6] ;
 wire \MOS6502.ALU.temp[7] ;
 wire \MOS6502.ALU.temp_BI[7] ;
 wire \MOS6502.ALU.temp_HC ;
 wire \MOS6502.AXYS[0][0] ;
 wire \MOS6502.AXYS[0][1] ;
 wire \MOS6502.AXYS[0][2] ;
 wire \MOS6502.AXYS[0][3] ;
 wire \MOS6502.AXYS[0][4] ;
 wire \MOS6502.AXYS[0][5] ;
 wire \MOS6502.AXYS[0][6] ;
 wire \MOS6502.AXYS[0][7] ;
 wire \MOS6502.AXYS[1][0] ;
 wire \MOS6502.AXYS[1][1] ;
 wire \MOS6502.AXYS[1][2] ;
 wire \MOS6502.AXYS[1][3] ;
 wire \MOS6502.AXYS[1][4] ;
 wire \MOS6502.AXYS[1][5] ;
 wire \MOS6502.AXYS[1][6] ;
 wire \MOS6502.AXYS[1][7] ;
 wire \MOS6502.AXYS[2][0] ;
 wire \MOS6502.AXYS[2][1] ;
 wire \MOS6502.AXYS[2][2] ;
 wire \MOS6502.AXYS[2][3] ;
 wire \MOS6502.AXYS[2][4] ;
 wire \MOS6502.AXYS[2][5] ;
 wire \MOS6502.AXYS[2][6] ;
 wire \MOS6502.AXYS[2][7] ;
 wire \MOS6502.AXYS[3][0] ;
 wire \MOS6502.AXYS[3][1] ;
 wire \MOS6502.AXYS[3][2] ;
 wire \MOS6502.AXYS[3][3] ;
 wire \MOS6502.AXYS[3][4] ;
 wire \MOS6502.AXYS[3][5] ;
 wire \MOS6502.AXYS[3][6] ;
 wire \MOS6502.AXYS[3][7] ;
 wire \MOS6502.C ;
 wire \MOS6502.D ;
 wire \MOS6502.I ;
 wire \MOS6502.IRHOLD[0] ;
 wire \MOS6502.IRHOLD[1] ;
 wire \MOS6502.IRHOLD[2] ;
 wire \MOS6502.IRHOLD[3] ;
 wire \MOS6502.IRHOLD[4] ;
 wire \MOS6502.IRHOLD[5] ;
 wire \MOS6502.IRHOLD[6] ;
 wire \MOS6502.IRHOLD[7] ;
 wire \MOS6502.IRHOLD_valid ;
 wire \MOS6502.IR[5] ;
 wire \MOS6502.IR[6] ;
 wire \MOS6502.IR[7] ;
 wire \MOS6502.N ;
 wire \MOS6502.NMI_1 ;
 wire \MOS6502.NMI_edge ;
 wire \MOS6502.PC[0] ;
 wire \MOS6502.PC[10] ;
 wire \MOS6502.PC[11] ;
 wire \MOS6502.PC[12] ;
 wire \MOS6502.PC[13] ;
 wire \MOS6502.PC[14] ;
 wire \MOS6502.PC[15] ;
 wire \MOS6502.PC[1] ;
 wire \MOS6502.PC[2] ;
 wire \MOS6502.PC[3] ;
 wire \MOS6502.PC[4] ;
 wire \MOS6502.PC[5] ;
 wire \MOS6502.PC[6] ;
 wire \MOS6502.PC[7] ;
 wire \MOS6502.PC[8] ;
 wire \MOS6502.PC[9] ;
 wire \MOS6502.V ;
 wire \MOS6502.Z ;
 wire \MOS6502.adc_bcd ;
 wire \MOS6502.adc_sbc ;
 wire \MOS6502.adj_bcd ;
 wire \MOS6502.backwards ;
 wire \MOS6502.bit_ins ;
 wire \MOS6502.clc ;
 wire \MOS6502.cld ;
 wire \MOS6502.cli ;
 wire \MOS6502.clv ;
 wire \MOS6502.compare ;
 wire \MOS6502.cond_code[0] ;
 wire \MOS6502.cond_code[1] ;
 wire \MOS6502.cond_code[2] ;
 wire \MOS6502.dst_reg[0] ;
 wire \MOS6502.dst_reg[1] ;
 wire \MOS6502.inc ;
 wire \MOS6502.index_y ;
 wire \MOS6502.load_only ;
 wire \MOS6502.load_reg ;
 wire \MOS6502.op[0] ;
 wire \MOS6502.op[1] ;
 wire \MOS6502.op[2] ;
 wire \MOS6502.op[3] ;
 wire \MOS6502.php ;
 wire \MOS6502.plp ;
 wire \MOS6502.res ;
 wire \MOS6502.rotate ;
 wire \MOS6502.sec ;
 wire \MOS6502.sed ;
 wire \MOS6502.sei ;
 wire \MOS6502.shift ;
 wire \MOS6502.shift_right ;
 wire \MOS6502.src_reg[0] ;
 wire \MOS6502.src_reg[1] ;
 wire \MOS6502.state[0] ;
 wire \MOS6502.state[1] ;
 wire \MOS6502.state[2] ;
 wire \MOS6502.state[3] ;
 wire \MOS6502.state[4] ;
 wire \MOS6502.state[5] ;
 wire \MOS6502.store ;
 wire \MOS6502.write_back ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0318_));
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__inv_2 _0828_ (.A(\MOS6502.NMI_edge ),
    .Y(_0221_));
 sky130_fd_sc_hd__inv_2 _0829_ (.A(\MOS6502.I ),
    .Y(_0222_));
 sky130_fd_sc_hd__clkinv_2 _0830_ (.A(net83),
    .Y(_0223_));
 sky130_fd_sc_hd__inv_2 _0831_ (.A(\MOS6502.cld ),
    .Y(_0224_));
 sky130_fd_sc_hd__inv_2 _0832_ (.A(\MOS6502.cli ),
    .Y(_0225_));
 sky130_fd_sc_hd__inv_2 _0833_ (.A(\MOS6502.load_only ),
    .Y(_0226_));
 sky130_fd_sc_hd__inv_2 _0834_ (.A(\MOS6502.shift ),
    .Y(_0227_));
 sky130_fd_sc_hd__inv_2 _0835_ (.A(\MOS6502.rotate ),
    .Y(_0228_));
 sky130_fd_sc_hd__inv_2 _0836_ (.A(net11),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _0837_ (.A(\MOS6502.clc ),
    .Y(_0229_));
 sky130_fd_sc_hd__a21oi_2 _0838_ (.A1(_0222_),
    .A2(net9),
    .B1(\MOS6502.NMI_edge ),
    .Y(_0230_));
 sky130_fd_sc_hd__mux2_8 _0839_ (.A0(net8),
    .A1(\MOS6502.IRHOLD[7] ),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0231_));
 sky130_fd_sc_hd__nand2_8 _0840_ (.A(net70),
    .B(_0231_),
    .Y(_0232_));
 sky130_fd_sc_hd__clkinv_4 _0841_ (.A(_0232_),
    .Y(\MOS6502.IR[7] ));
 sky130_fd_sc_hd__mux2_2 _0842_ (.A0(net6),
    .A1(\MOS6502.IRHOLD[5] ),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0233_));
 sky130_fd_sc_hd__nand2_2 _0843_ (.A(net70),
    .B(_0233_),
    .Y(_0234_));
 sky130_fd_sc_hd__clkinv_4 _0844_ (.A(net52),
    .Y(\MOS6502.IR[5] ));
 sky130_fd_sc_hd__mux2_4 _0845_ (.A0(net7),
    .A1(\MOS6502.IRHOLD[6] ),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0235_));
 sky130_fd_sc_hd__nand2_8 _0846_ (.A(net71),
    .B(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__inv_2 _0847_ (.A(_0236_),
    .Y(\MOS6502.IR[6] ));
 sky130_fd_sc_hd__nand2b_1 _0848_ (.A_N(\MOS6502.state[5] ),
    .B(net80),
    .Y(_0237_));
 sky130_fd_sc_hd__nand2_2 _0849_ (.A(net86),
    .B(net88),
    .Y(_0238_));
 sky130_fd_sc_hd__and4b_1 _0850_ (.A_N(net85),
    .B(net83),
    .C(net86),
    .D(net89),
    .X(_0239_));
 sky130_fd_sc_hd__or3_4 _0851_ (.A(net84),
    .B(_0223_),
    .C(_0238_),
    .X(_0240_));
 sky130_fd_sc_hd__nor2_1 _0852_ (.A(net80),
    .B(\MOS6502.state[5] ),
    .Y(_0241_));
 sky130_fd_sc_hd__or2_4 _0853_ (.A(net80),
    .B(\MOS6502.state[5] ),
    .X(_0242_));
 sky130_fd_sc_hd__nand2b_2 _0854_ (.A_N(net87),
    .B(net89),
    .Y(_0243_));
 sky130_fd_sc_hd__or3_4 _0855_ (.A(net84),
    .B(_0223_),
    .C(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__or2_4 _0856_ (.A(net75),
    .B(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__o21ai_2 _0857_ (.A1(net77),
    .A2(_0240_),
    .B1(_0245_),
    .Y(_0246_));
 sky130_fd_sc_hd__or4bb_4 _0858_ (.A(net88),
    .B(net84),
    .C_N(net82),
    .D_N(net87),
    .X(_0247_));
 sky130_fd_sc_hd__nor2_2 _0859_ (.A(_0242_),
    .B(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__or2_1 _0860_ (.A(net75),
    .B(_0247_),
    .X(_0249_));
 sky130_fd_sc_hd__nor2_1 _0861_ (.A(net78),
    .B(_0247_),
    .Y(_0250_));
 sky130_fd_sc_hd__nand2b_2 _0862_ (.A_N(net80),
    .B(\MOS6502.state[5] ),
    .Y(_0251_));
 sky130_fd_sc_hd__or4b_4 _0863_ (.A(net88),
    .B(net84),
    .C(net82),
    .D_N(net86),
    .X(_0252_));
 sky130_fd_sc_hd__nor2_8 _0864_ (.A(net74),
    .B(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__or2_4 _0865_ (.A(net74),
    .B(_0252_),
    .X(_0254_));
 sky130_fd_sc_hd__nor2_1 _0866_ (.A(net86),
    .B(net89),
    .Y(_0255_));
 sky130_fd_sc_hd__or4b_4 _0867_ (.A(net87),
    .B(net89),
    .C(net85),
    .D_N(net83),
    .X(_0256_));
 sky130_fd_sc_hd__or3b_4 _0868_ (.A(_0223_),
    .B(net76),
    .C_N(_0255_),
    .X(_0257_));
 sky130_fd_sc_hd__nor2_2 _0869_ (.A(net76),
    .B(_0256_),
    .Y(_0258_));
 sky130_fd_sc_hd__or2_2 _0870_ (.A(net67),
    .B(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__or4_4 _0871_ (.A(net48),
    .B(net69),
    .C(_0253_),
    .D(net51),
    .X(_0260_));
 sky130_fd_sc_hd__and2_1 _0872_ (.A(net85),
    .B(net83),
    .X(_0261_));
 sky130_fd_sc_hd__nand2_4 _0873_ (.A(\MOS6502.state[2] ),
    .B(net82),
    .Y(_0262_));
 sky130_fd_sc_hd__or3_1 _0874_ (.A(net88),
    .B(net74),
    .C(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__nand4b_4 _0875_ (.A_N(net89),
    .B(net85),
    .C(net83),
    .D(net86),
    .Y(_0264_));
 sky130_fd_sc_hd__nor2_2 _0876_ (.A(net73),
    .B(_0264_),
    .Y(_0265_));
 sky130_fd_sc_hd__nor2_4 _0877_ (.A(_0260_),
    .B(net65),
    .Y(_0266_));
 sky130_fd_sc_hd__or2_4 _0878_ (.A(_0260_),
    .B(net65),
    .X(_0267_));
 sky130_fd_sc_hd__or4b_4 _0879_ (.A(net86),
    .B(net89),
    .C(net83),
    .D_N(net85),
    .X(_0268_));
 sky130_fd_sc_hd__nor2_2 _0880_ (.A(net75),
    .B(_0268_),
    .Y(_0269_));
 sky130_fd_sc_hd__or3_4 _0881_ (.A(\MOS6502.state[2] ),
    .B(net82),
    .C(_0243_),
    .X(_0270_));
 sky130_fd_sc_hd__nor2_4 _0882_ (.A(net75),
    .B(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__and2_1 _0883_ (.A(net80),
    .B(\MOS6502.state[5] ),
    .X(_0272_));
 sky130_fd_sc_hd__nand2_2 _0884_ (.A(net81),
    .B(\MOS6502.state[5] ),
    .Y(_0273_));
 sky130_fd_sc_hd__nor2_1 _0885_ (.A(_0270_),
    .B(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__nor3_1 _0886_ (.A(_0238_),
    .B(net73),
    .C(_0262_),
    .Y(_0275_));
 sky130_fd_sc_hd__or4_4 _0887_ (.A(_0269_),
    .B(_0271_),
    .C(_0274_),
    .D(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__inv_2 _0888_ (.A(_0276_),
    .Y(_0277_));
 sky130_fd_sc_hd__or2_2 _0889_ (.A(net82),
    .B(_0243_),
    .X(_0278_));
 sky130_fd_sc_hd__nor2_1 _0890_ (.A(net78),
    .B(_0278_),
    .Y(_0279_));
 sky130_fd_sc_hd__o21a_1 _0891_ (.A1(_0276_),
    .A2(_0279_),
    .B1(\MOS6502.store ),
    .X(_0280_));
 sky130_fd_sc_hd__nor2_2 _0892_ (.A(_0267_),
    .B(_0280_),
    .Y(net12));
 sky130_fd_sc_hd__inv_2 _0893_ (.A(net12),
    .Y(net31));
 sky130_fd_sc_hd__or2_4 _0894_ (.A(_0243_),
    .B(_0262_),
    .X(_0281_));
 sky130_fd_sc_hd__nor2_2 _0895_ (.A(net76),
    .B(_0281_),
    .Y(_0282_));
 sky130_fd_sc_hd__or2_1 _0896_ (.A(net75),
    .B(_0281_),
    .X(_0283_));
 sky130_fd_sc_hd__or4bb_4 _0897_ (.A(net85),
    .B(net83),
    .C_N(net86),
    .D_N(net89),
    .X(_0284_));
 sky130_fd_sc_hd__nor2_2 _0898_ (.A(net73),
    .B(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__nor2_2 _0899_ (.A(net73),
    .B(_0268_),
    .Y(_0286_));
 sky130_fd_sc_hd__or2_4 _0900_ (.A(_0285_),
    .B(_0286_),
    .X(_0287_));
 sky130_fd_sc_hd__or2_4 _0901_ (.A(_0282_),
    .B(_0287_),
    .X(_0288_));
 sky130_fd_sc_hd__and2_2 _0902_ (.A(\MOS6502.shift_right ),
    .B(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__nand2_2 _0903_ (.A(\MOS6502.shift_right ),
    .B(_0288_),
    .Y(_0290_));
 sky130_fd_sc_hd__or2_1 _0904_ (.A(net73),
    .B(_0278_),
    .X(_0291_));
 sky130_fd_sc_hd__or4bb_4 _0905_ (.A(net87),
    .B(net82),
    .C_N(net84),
    .D_N(net88),
    .X(_0292_));
 sky130_fd_sc_hd__nor2_1 _0906_ (.A(net73),
    .B(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__a21oi_4 _0907_ (.A1(_0247_),
    .A2(_0292_),
    .B1(net74),
    .Y(_0294_));
 sky130_fd_sc_hd__nor2_2 _0908_ (.A(net67),
    .B(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__nor3_2 _0909_ (.A(net89),
    .B(net77),
    .C(_0262_),
    .Y(_0296_));
 sky130_fd_sc_hd__and2b_4 _0910_ (.A_N(net86),
    .B(_0296_),
    .X(_0297_));
 sky130_fd_sc_hd__nor4_2 _0911_ (.A(_0253_),
    .B(_0258_),
    .C(_0286_),
    .D(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__or2_1 _0912_ (.A(net77),
    .B(_0264_),
    .X(_0299_));
 sky130_fd_sc_hd__o21a_2 _0913_ (.A1(net85),
    .A2(_0291_),
    .B1(_0299_),
    .X(_0300_));
 sky130_fd_sc_hd__nor2_1 _0914_ (.A(net80),
    .B(_0252_),
    .Y(_0301_));
 sky130_fd_sc_hd__nor2_1 _0915_ (.A(net77),
    .B(_0284_),
    .Y(_0302_));
 sky130_fd_sc_hd__o22ai_4 _0916_ (.A1(net76),
    .A2(_0264_),
    .B1(_0284_),
    .B2(net78),
    .Y(_0303_));
 sky130_fd_sc_hd__or4_4 _0917_ (.A(net87),
    .B(net88),
    .C(net84),
    .D(net82),
    .X(_0304_));
 sky130_fd_sc_hd__inv_2 _0918_ (.A(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__nor2_4 _0919_ (.A(_0273_),
    .B(_0304_),
    .Y(_0306_));
 sky130_fd_sc_hd__or2_2 _0920_ (.A(_0303_),
    .B(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__o221a_1 _0921_ (.A1(net80),
    .A2(_0252_),
    .B1(_0283_),
    .B2(\MOS6502.load_only ),
    .C1(_0300_),
    .X(_0308_));
 sky130_fd_sc_hd__nor2_1 _0922_ (.A(_0258_),
    .B(_0307_),
    .Y(_0309_));
 sky130_fd_sc_hd__and4_4 _0923_ (.A(_0295_),
    .B(_0298_),
    .C(_0308_),
    .D(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__inv_2 _0924_ (.A(_0310_),
    .Y(_0311_));
 sky130_fd_sc_hd__nor2_4 _0925_ (.A(net76),
    .B(_0252_),
    .Y(_0312_));
 sky130_fd_sc_hd__and3_2 _0926_ (.A(_0241_),
    .B(_0255_),
    .C(_0261_),
    .X(_0313_));
 sky130_fd_sc_hd__or4_1 _0927_ (.A(net86),
    .B(net88),
    .C(net75),
    .D(_0262_),
    .X(_0314_));
 sky130_fd_sc_hd__nor4_4 _0928_ (.A(_0303_),
    .B(_0306_),
    .C(_0312_),
    .D(net64),
    .Y(_0315_));
 sky130_fd_sc_hd__o22ai_1 _0929_ (.A1(net80),
    .A2(_0256_),
    .B1(_0264_),
    .B2(net78),
    .Y(_0316_));
 sky130_fd_sc_hd__or3_4 _0930_ (.A(net78),
    .B(_0238_),
    .C(_0262_),
    .X(_0317_));
 sky130_fd_sc_hd__nor2_4 _0931_ (.A(_0240_),
    .B(net76),
    .Y(_0318_));
 sky130_fd_sc_hd__and2_2 _0932_ (.A(net77),
    .B(net74),
    .X(_0319_));
 sky130_fd_sc_hd__xor2_2 _0933_ (.A(net81),
    .B(\MOS6502.state[5] ),
    .X(_0320_));
 sky130_fd_sc_hd__a32o_1 _0934_ (.A1(_0255_),
    .A2(_0261_),
    .A3(_0320_),
    .B1(_0241_),
    .B2(_0239_),
    .X(_0321_));
 sky130_fd_sc_hd__and4bb_2 _0935_ (.A_N(_0316_),
    .B_N(_0321_),
    .C(_0317_),
    .D(_0254_),
    .X(_0322_));
 sky130_fd_sc_hd__nand4b_4 _0936_ (.A_N(\MOS6502.src_reg[0] ),
    .B(_0295_),
    .C(_0315_),
    .D(_0322_),
    .Y(_0323_));
 sky130_fd_sc_hd__o31a_1 _0937_ (.A1(_0303_),
    .A2(_0306_),
    .A3(_0312_),
    .B1(\MOS6502.index_y ),
    .X(_0324_));
 sky130_fd_sc_hd__a211o_4 _0938_ (.A1(\MOS6502.dst_reg[0] ),
    .A2(net63),
    .B1(_0315_),
    .C1(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__and2_4 _0939_ (.A(_0323_),
    .B(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__nand2_8 _0940_ (.A(_0323_),
    .B(_0325_),
    .Y(_0327_));
 sky130_fd_sc_hd__and4_1 _0941_ (.A(\MOS6502.src_reg[1] ),
    .B(_0295_),
    .C(_0315_),
    .D(_0322_),
    .X(_0328_));
 sky130_fd_sc_hd__a2111o_4 _0942_ (.A1(\MOS6502.dst_reg[1] ),
    .A2(net64),
    .B1(_0328_),
    .C1(_0307_),
    .D1(_0312_),
    .X(_0329_));
 sky130_fd_sc_hd__or2_1 _0943_ (.A(\MOS6502.AXYS[2][6] ),
    .B(_0326_),
    .X(_0330_));
 sky130_fd_sc_hd__o211a_1 _0944_ (.A1(\MOS6502.AXYS[3][6] ),
    .A2(net45),
    .B1(net44),
    .C1(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__nor2_8 _0945_ (.A(_0326_),
    .B(net44),
    .Y(_0332_));
 sky130_fd_sc_hd__nor2_8 _0946_ (.A(_0327_),
    .B(net44),
    .Y(_0333_));
 sky130_fd_sc_hd__a221oi_4 _0947_ (.A1(\MOS6502.AXYS[0][6] ),
    .A2(_0332_),
    .B1(_0333_),
    .B2(\MOS6502.AXYS[1][6] ),
    .C1(_0331_),
    .Y(_0334_));
 sky130_fd_sc_hd__nor2_1 _0948_ (.A(_0310_),
    .B(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__nor2_8 _0949_ (.A(net75),
    .B(_0292_),
    .Y(_0336_));
 sky130_fd_sc_hd__or2_4 _0950_ (.A(_0285_),
    .B(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__or4bb_4 _0951_ (.A(net88),
    .B(net82),
    .C_N(net84),
    .D_N(net87),
    .X(_0338_));
 sky130_fd_sc_hd__nor2_1 _0952_ (.A(net75),
    .B(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__or3_4 _0953_ (.A(_0238_),
    .B(_0242_),
    .C(_0262_),
    .X(_0340_));
 sky130_fd_sc_hd__or3b_4 _0954_ (.A(net82),
    .B(_0238_),
    .C_N(net84),
    .X(_0341_));
 sky130_fd_sc_hd__a31o_1 _0955_ (.A1(_0240_),
    .A2(_0338_),
    .A3(_0341_),
    .B1(net74),
    .X(_0342_));
 sky130_fd_sc_hd__and2_1 _0956_ (.A(_0340_),
    .B(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__or3b_4 _0957_ (.A(_0246_),
    .B(net69),
    .C_N(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__a221o_2 _0958_ (.A1(\MOS6502.ABH[6] ),
    .A2(net53),
    .B1(_0344_),
    .B2(\MOS6502.ADD[6] ),
    .C1(_0335_),
    .X(_0345_));
 sky130_fd_sc_hd__a21oi_4 _0959_ (.A1(net7),
    .A2(_0337_),
    .B1(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__nor2_1 _0960_ (.A(net46),
    .B(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__or2_1 _0961_ (.A(\MOS6502.AXYS[2][5] ),
    .B(_0326_),
    .X(_0348_));
 sky130_fd_sc_hd__o211a_1 _0962_ (.A1(\MOS6502.AXYS[3][5] ),
    .A2(net45),
    .B1(net44),
    .C1(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__a221oi_4 _0963_ (.A1(\MOS6502.AXYS[0][5] ),
    .A2(_0332_),
    .B1(_0333_),
    .B2(\MOS6502.AXYS[1][5] ),
    .C1(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__nor2_1 _0964_ (.A(_0310_),
    .B(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__a221o_2 _0965_ (.A1(\MOS6502.ABH[5] ),
    .A2(net53),
    .B1(_0344_),
    .B2(\MOS6502.ADD[5] ),
    .C1(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__a21oi_4 _0966_ (.A1(net6),
    .A2(_0337_),
    .B1(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hd__nor2_4 _0967_ (.A(net73),
    .B(_0341_),
    .Y(_0354_));
 sky130_fd_sc_hd__or2_4 _0968_ (.A(net73),
    .B(_0341_),
    .X(_0355_));
 sky130_fd_sc_hd__o21ai_1 _0969_ (.A1(net80),
    .A2(_0338_),
    .B1(_0340_),
    .Y(_0356_));
 sky130_fd_sc_hd__nor2_1 _0970_ (.A(_0247_),
    .B(_0272_),
    .Y(_0357_));
 sky130_fd_sc_hd__a21o_1 _0971_ (.A1(_0239_),
    .A2(_0320_),
    .B1(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__or4bb_1 _0972_ (.A(_0356_),
    .B(_0358_),
    .C_N(_0299_),
    .D_N(_0355_),
    .X(_0359_));
 sky130_fd_sc_hd__and4b_1 _0973_ (.A_N(_0337_),
    .B(_0291_),
    .C(_0245_),
    .D(_0298_),
    .X(_0360_));
 sky130_fd_sc_hd__and2b_4 _0974_ (.A_N(_0359_),
    .B(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__a22o_2 _0975_ (.A1(\MOS6502.PC[5] ),
    .A2(_0336_),
    .B1(_0361_),
    .B2(net6),
    .X(_0362_));
 sky130_fd_sc_hd__and2b_1 _0976_ (.A_N(_0353_),
    .B(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__nor3_4 _0977_ (.A(_0271_),
    .B(_0288_),
    .C(net64),
    .Y(_0364_));
 sky130_fd_sc_hd__a21oi_4 _0978_ (.A1(\MOS6502.op[0] ),
    .A2(_0288_),
    .B1(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__a21bo_1 _0979_ (.A1(_0362_),
    .A2(net42),
    .B1_N(_0353_),
    .X(_0366_));
 sky130_fd_sc_hd__a21oi_4 _0980_ (.A1(\MOS6502.op[1] ),
    .A2(_0288_),
    .B1(_0364_),
    .Y(_0367_));
 sky130_fd_sc_hd__a21o_1 _0981_ (.A1(\MOS6502.op[1] ),
    .A2(_0288_),
    .B1(_0364_),
    .X(_0368_));
 sky130_fd_sc_hd__or2_2 _0982_ (.A(net42),
    .B(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__and2_1 _0983_ (.A(net42),
    .B(_0368_),
    .X(_0370_));
 sky130_fd_sc_hd__inv_2 _0984_ (.A(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__nor2_1 _0985_ (.A(_0365_),
    .B(_0367_),
    .Y(_0372_));
 sky130_fd_sc_hd__mux2_1 _0986_ (.A0(_0369_),
    .A1(_0371_),
    .S(_0363_),
    .X(_0373_));
 sky130_fd_sc_hd__a31o_2 _0987_ (.A1(net46),
    .A2(_0366_),
    .A3(_0373_),
    .B1(_0347_),
    .X(_0374_));
 sky130_fd_sc_hd__a221o_4 _0988_ (.A1(\MOS6502.op[2] ),
    .A2(_0288_),
    .B1(net53),
    .B2(\MOS6502.backwards ),
    .C1(_0260_),
    .X(_0375_));
 sky130_fd_sc_hd__inv_2 _0989_ (.A(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__and2_4 _0990_ (.A(\MOS6502.op[3] ),
    .B(_0288_),
    .X(_0377_));
 sky130_fd_sc_hd__inv_2 _0991_ (.A(_0377_),
    .Y(_0378_));
 sky130_fd_sc_hd__nor2_1 _0992_ (.A(_0375_),
    .B(_0377_),
    .Y(_0379_));
 sky130_fd_sc_hd__mux2_1 _0993_ (.A0(_0379_),
    .A1(_0375_),
    .S(_0362_),
    .X(_0380_));
 sky130_fd_sc_hd__nor2_2 _0994_ (.A(_0376_),
    .B(_0378_),
    .Y(_0381_));
 sky130_fd_sc_hd__or2_2 _0995_ (.A(_0380_),
    .B(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__nand2b_4 _0996_ (.A_N(_0382_),
    .B(_0374_),
    .Y(_0383_));
 sky130_fd_sc_hd__or2_1 _0997_ (.A(\MOS6502.AXYS[2][4] ),
    .B(_0326_),
    .X(_0384_));
 sky130_fd_sc_hd__o211a_1 _0998_ (.A1(\MOS6502.AXYS[3][4] ),
    .A2(net45),
    .B1(net44),
    .C1(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__a221oi_4 _0999_ (.A1(\MOS6502.AXYS[0][4] ),
    .A2(_0332_),
    .B1(_0333_),
    .B2(\MOS6502.AXYS[1][4] ),
    .C1(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__a22o_1 _1000_ (.A1(net5),
    .A2(_0337_),
    .B1(net53),
    .B2(\MOS6502.ABH[4] ),
    .X(_0387_));
 sky130_fd_sc_hd__a21oi_1 _1001_ (.A1(\MOS6502.ADD[4] ),
    .A2(_0344_),
    .B1(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__o21a_2 _1002_ (.A1(_0310_),
    .A2(_0386_),
    .B1(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__a22o_2 _1003_ (.A1(\MOS6502.PC[4] ),
    .A2(_0336_),
    .B1(_0361_),
    .B2(net5),
    .X(_0390_));
 sky130_fd_sc_hd__nand2_1 _1004_ (.A(net42),
    .B(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__o21ai_1 _1005_ (.A1(_0389_),
    .A2(_0391_),
    .B1(_0369_),
    .Y(_0392_));
 sky130_fd_sc_hd__or3b_1 _1006_ (.A(_0368_),
    .B(_0389_),
    .C_N(_0390_),
    .X(_0393_));
 sky130_fd_sc_hd__a22o_1 _1007_ (.A1(_0389_),
    .A2(_0391_),
    .B1(_0392_),
    .B2(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _1008_ (.A0(_0353_),
    .A1(_0394_),
    .S(net46),
    .X(_0395_));
 sky130_fd_sc_hd__or2_4 _1009_ (.A(_0379_),
    .B(_0381_),
    .X(_0396_));
 sky130_fd_sc_hd__inv_2 _1010_ (.A(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__mux2_1 _1011_ (.A0(_0396_),
    .A1(_0375_),
    .S(_0390_),
    .X(_0398_));
 sky130_fd_sc_hd__nor2_2 _1012_ (.A(_0395_),
    .B(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__o21a_1 _1013_ (.A1(_0377_),
    .A2(_0398_),
    .B1(_0395_),
    .X(_0400_));
 sky130_fd_sc_hd__or2_2 _1014_ (.A(_0399_),
    .B(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__or2_1 _1015_ (.A(\MOS6502.AXYS[2][3] ),
    .B(_0326_),
    .X(_0402_));
 sky130_fd_sc_hd__o211a_1 _1016_ (.A1(\MOS6502.AXYS[3][3] ),
    .A2(_0327_),
    .B1(_0329_),
    .C1(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__a221oi_4 _1017_ (.A1(\MOS6502.AXYS[0][3] ),
    .A2(_0332_),
    .B1(_0333_),
    .B2(\MOS6502.AXYS[1][3] ),
    .C1(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__a22o_1 _1018_ (.A1(net4),
    .A2(_0337_),
    .B1(net54),
    .B2(\MOS6502.ABH[3] ),
    .X(_0405_));
 sky130_fd_sc_hd__a21oi_1 _1019_ (.A1(\MOS6502.ADD[3] ),
    .A2(_0344_),
    .B1(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__o21a_2 _1020_ (.A1(_0310_),
    .A2(_0404_),
    .B1(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__a22o_2 _1021_ (.A1(\MOS6502.PC[3] ),
    .A2(_0336_),
    .B1(_0361_),
    .B2(net4),
    .X(_0408_));
 sky130_fd_sc_hd__nand2_1 _1022_ (.A(_0365_),
    .B(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__o21ai_1 _1023_ (.A1(_0407_),
    .A2(_0409_),
    .B1(_0369_),
    .Y(_0410_));
 sky130_fd_sc_hd__nand2_1 _1024_ (.A(_0367_),
    .B(_0408_),
    .Y(_0411_));
 sky130_fd_sc_hd__o21a_1 _1025_ (.A1(_0407_),
    .A2(_0411_),
    .B1(_0410_),
    .X(_0412_));
 sky130_fd_sc_hd__a21o_1 _1026_ (.A1(_0407_),
    .A2(_0409_),
    .B1(_0289_),
    .X(_0413_));
 sky130_fd_sc_hd__o22a_1 _1027_ (.A1(net46),
    .A2(_0389_),
    .B1(_0412_),
    .B2(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_2 _1028_ (.A0(_0396_),
    .A1(_0375_),
    .S(_0408_),
    .X(_0415_));
 sky130_fd_sc_hd__inv_2 _1029_ (.A(_0415_),
    .Y(_0416_));
 sky130_fd_sc_hd__or2_1 _1030_ (.A(_0377_),
    .B(_0415_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_4 _1031_ (.A0(_0416_),
    .A1(_0417_),
    .S(_0414_),
    .X(_0418_));
 sky130_fd_sc_hd__and3_1 _1032_ (.A(\MOS6502.AXYS[1][2] ),
    .B(_0323_),
    .C(_0325_),
    .X(_0419_));
 sky130_fd_sc_hd__a21oi_1 _1033_ (.A1(\MOS6502.AXYS[0][2] ),
    .A2(net45),
    .B1(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__a21o_1 _1034_ (.A1(_0323_),
    .A2(_0325_),
    .B1(\MOS6502.AXYS[2][2] ),
    .X(_0421_));
 sky130_fd_sc_hd__o21ai_1 _1035_ (.A1(\MOS6502.AXYS[3][2] ),
    .A2(net45),
    .B1(_0421_),
    .Y(_0422_));
 sky130_fd_sc_hd__mux2_2 _1036_ (.A0(_0420_),
    .A1(_0422_),
    .S(net44),
    .X(_0423_));
 sky130_fd_sc_hd__a22o_1 _1037_ (.A1(net3),
    .A2(_0337_),
    .B1(net53),
    .B2(\MOS6502.ABH[2] ),
    .X(_0424_));
 sky130_fd_sc_hd__a21oi_1 _1038_ (.A1(\MOS6502.ADD[2] ),
    .A2(_0344_),
    .B1(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hd__o21a_2 _1039_ (.A1(_0310_),
    .A2(_0423_),
    .B1(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__a22o_2 _1040_ (.A1(\MOS6502.PC[2] ),
    .A2(_0336_),
    .B1(_0361_),
    .B2(net3),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_1 _1041_ (.A(_0365_),
    .B(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__o21a_1 _1042_ (.A1(_0426_),
    .A2(_0428_),
    .B1(_0369_),
    .X(_0429_));
 sky130_fd_sc_hd__nor2_1 _1043_ (.A(_0368_),
    .B(_0426_),
    .Y(_0430_));
 sky130_fd_sc_hd__a21oi_1 _1044_ (.A1(_0427_),
    .A2(_0430_),
    .B1(_0429_),
    .Y(_0431_));
 sky130_fd_sc_hd__a21o_1 _1045_ (.A1(_0426_),
    .A2(_0428_),
    .B1(_0289_),
    .X(_0432_));
 sky130_fd_sc_hd__o22a_1 _1046_ (.A1(net46),
    .A2(_0407_),
    .B1(_0431_),
    .B2(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _1047_ (.A0(_0396_),
    .A1(_0375_),
    .S(_0427_),
    .X(_0434_));
 sky130_fd_sc_hd__or2_4 _1048_ (.A(_0433_),
    .B(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__nor2_1 _1049_ (.A(net46),
    .B(_0426_),
    .Y(_0436_));
 sky130_fd_sc_hd__mux2_1 _1050_ (.A0(\MOS6502.AXYS[1][1] ),
    .A1(\MOS6502.AXYS[0][1] ),
    .S(_0327_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _1051_ (.A0(\MOS6502.AXYS[3][1] ),
    .A1(\MOS6502.AXYS[2][1] ),
    .S(net45),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_4 _1052_ (.A0(_0437_),
    .A1(_0438_),
    .S(_0329_),
    .X(_0439_));
 sky130_fd_sc_hd__a22o_1 _1053_ (.A1(net2),
    .A2(_0337_),
    .B1(net54),
    .B2(\MOS6502.ABH[1] ),
    .X(_0440_));
 sky130_fd_sc_hd__a21o_1 _1054_ (.A1(\MOS6502.ADD[1] ),
    .A2(_0344_),
    .B1(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__a21oi_2 _1055_ (.A1(_0311_),
    .A2(_0439_),
    .B1(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__a22o_2 _1056_ (.A1(\MOS6502.PC[1] ),
    .A2(_0336_),
    .B1(_0361_),
    .B2(net2),
    .X(_0443_));
 sky130_fd_sc_hd__and2b_1 _1057_ (.A_N(_0442_),
    .B(_0443_),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _1058_ (.A0(net42),
    .A1(_0367_),
    .S(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__a21bo_1 _1059_ (.A1(net42),
    .A2(_0443_),
    .B1_N(_0442_),
    .X(_0446_));
 sky130_fd_sc_hd__o211a_1 _1060_ (.A1(_0372_),
    .A2(_0445_),
    .B1(_0446_),
    .C1(net46),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _1061_ (.A0(_0397_),
    .A1(_0376_),
    .S(_0443_),
    .X(_0448_));
 sky130_fd_sc_hd__o21a_1 _1062_ (.A1(_0436_),
    .A2(_0447_),
    .B1(_0448_),
    .X(_0449_));
 sky130_fd_sc_hd__or2_2 _1063_ (.A(net46),
    .B(_0442_),
    .X(_0450_));
 sky130_fd_sc_hd__a22oi_4 _1064_ (.A1(\MOS6502.PC[0] ),
    .A2(_0336_),
    .B1(_0361_),
    .B2(net1),
    .Y(_0451_));
 sky130_fd_sc_hd__and3_1 _1065_ (.A(\MOS6502.AXYS[1][0] ),
    .B(_0323_),
    .C(_0325_),
    .X(_0452_));
 sky130_fd_sc_hd__a21oi_1 _1066_ (.A1(\MOS6502.AXYS[0][0] ),
    .A2(net45),
    .B1(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__a21o_1 _1067_ (.A1(_0323_),
    .A2(_0325_),
    .B1(\MOS6502.AXYS[2][0] ),
    .X(_0454_));
 sky130_fd_sc_hd__o21ai_1 _1068_ (.A1(\MOS6502.AXYS[3][0] ),
    .A2(net45),
    .B1(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__mux2_2 _1069_ (.A0(_0453_),
    .A1(_0455_),
    .S(net44),
    .X(_0456_));
 sky130_fd_sc_hd__a22o_1 _1070_ (.A1(net1),
    .A2(_0337_),
    .B1(net54),
    .B2(\MOS6502.ABH[0] ),
    .X(_0457_));
 sky130_fd_sc_hd__a21oi_1 _1071_ (.A1(\MOS6502.ADD[0] ),
    .A2(_0344_),
    .B1(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__o21a_4 _1072_ (.A1(_0310_),
    .A2(_0456_),
    .B1(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__o21ai_1 _1073_ (.A1(_0451_),
    .A2(_0459_),
    .B1(net42),
    .Y(_0460_));
 sky130_fd_sc_hd__a211o_1 _1074_ (.A1(_0367_),
    .A2(_0451_),
    .B1(_0459_),
    .C1(_0370_),
    .X(_0461_));
 sky130_fd_sc_hd__a221o_4 _1075_ (.A1(_0451_),
    .A2(_0459_),
    .B1(_0460_),
    .B2(_0461_),
    .C1(_0289_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_2 _1076_ (.A0(_0375_),
    .A1(_0396_),
    .S(_0451_),
    .X(_0463_));
 sky130_fd_sc_hd__a21oi_2 _1077_ (.A1(_0450_),
    .A2(_0462_),
    .B1(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__o211ai_4 _1078_ (.A1(_0377_),
    .A2(_0463_),
    .B1(_0462_),
    .C1(_0450_),
    .Y(_0465_));
 sky130_fd_sc_hd__and2b_1 _1079_ (.A_N(_0464_),
    .B(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__a32o_1 _1080_ (.A1(_0226_),
    .A2(_0227_),
    .A3(_0282_),
    .B1(_0288_),
    .B2(\MOS6502.rotate ),
    .X(_0467_));
 sky130_fd_sc_hd__nand2_1 _1081_ (.A(\MOS6502.C ),
    .B(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__a32o_1 _1082_ (.A1(_0227_),
    .A2(\MOS6502.inc ),
    .A3(_0287_),
    .B1(_0282_),
    .B2(\MOS6502.compare ),
    .X(_0469_));
 sky130_fd_sc_hd__nor2_1 _1083_ (.A(net76),
    .B(_0284_),
    .Y(_0470_));
 sky130_fd_sc_hd__nor2_1 _1084_ (.A(net77),
    .B(_0268_),
    .Y(_0471_));
 sky130_fd_sc_hd__or2_4 _1085_ (.A(_0470_),
    .B(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__o21a_1 _1086_ (.A1(net53),
    .A2(_0472_),
    .B1(\MOS6502.ALU.CO ),
    .X(_0473_));
 sky130_fd_sc_hd__a21oi_2 _1087_ (.A1(_0252_),
    .A2(_0264_),
    .B1(net78),
    .Y(_0474_));
 sky130_fd_sc_hd__or4b_1 _1088_ (.A(_0294_),
    .B(_0473_),
    .C(_0474_),
    .D_N(_0343_),
    .X(_0475_));
 sky130_fd_sc_hd__a21oi_1 _1089_ (.A1(_0228_),
    .A2(_0469_),
    .B1(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__nand2_2 _1090_ (.A(_0468_),
    .B(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__nor2_1 _1091_ (.A(_0289_),
    .B(_0381_),
    .Y(_0478_));
 sky130_fd_sc_hd__nand2_1 _1092_ (.A(_0477_),
    .B(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__a31o_4 _1093_ (.A1(_0465_),
    .A2(_0477_),
    .A3(_0478_),
    .B1(_0464_),
    .X(_0480_));
 sky130_fd_sc_hd__a211o_2 _1094_ (.A1(_0378_),
    .A2(_0448_),
    .B1(_0447_),
    .C1(_0436_),
    .X(_0481_));
 sky130_fd_sc_hd__nand2b_2 _1095_ (.A_N(_0449_),
    .B(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__a21oi_4 _1096_ (.A1(_0480_),
    .A2(_0481_),
    .B1(_0449_),
    .Y(_0483_));
 sky130_fd_sc_hd__o21ai_2 _1097_ (.A1(_0377_),
    .A2(_0434_),
    .B1(_0433_),
    .Y(_0484_));
 sky130_fd_sc_hd__nand2_4 _1098_ (.A(_0435_),
    .B(_0484_),
    .Y(_0485_));
 sky130_fd_sc_hd__o21a_1 _1099_ (.A1(_0483_),
    .A2(_0485_),
    .B1(_0435_),
    .X(_0486_));
 sky130_fd_sc_hd__nor2_1 _1100_ (.A(_0418_),
    .B(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__o22a_2 _1101_ (.A1(_0414_),
    .A2(_0415_),
    .B1(_0418_),
    .B2(_0486_),
    .X(_0488_));
 sky130_fd_sc_hd__xor2_4 _1102_ (.A(_0483_),
    .B(_0485_),
    .X(\MOS6502.ALU.temp[2] ));
 sky130_fd_sc_hd__xnor2_4 _1103_ (.A(_0480_),
    .B(_0482_),
    .Y(\MOS6502.ALU.temp[1] ));
 sky130_fd_sc_hd__o211ai_4 _1104_ (.A1(_0483_),
    .A2(_0485_),
    .B1(_0418_),
    .C1(_0435_),
    .Y(_0489_));
 sky130_fd_sc_hd__and2_2 _1105_ (.A(\MOS6502.adc_bcd ),
    .B(_0282_),
    .X(_0490_));
 sky130_fd_sc_hd__o211ai_4 _1106_ (.A1(\MOS6502.ALU.temp[2] ),
    .A2(\MOS6502.ALU.temp[1] ),
    .B1(_0489_),
    .C1(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__nand2_1 _1107_ (.A(_0488_),
    .B(_0491_),
    .Y(\MOS6502.ALU.temp_HC ));
 sky130_fd_sc_hd__a21oi_4 _1108_ (.A1(_0488_),
    .A2(_0491_),
    .B1(_0401_),
    .Y(_0492_));
 sky130_fd_sc_hd__o21bai_4 _1109_ (.A1(_0377_),
    .A2(_0382_),
    .B1_N(_0374_),
    .Y(_0493_));
 sky130_fd_sc_hd__o211ai_4 _1110_ (.A1(_0399_),
    .A2(_0492_),
    .B1(_0493_),
    .C1(_0383_),
    .Y(_0494_));
 sky130_fd_sc_hd__or2_1 _1111_ (.A(\MOS6502.AXYS[2][7] ),
    .B(_0326_),
    .X(_0495_));
 sky130_fd_sc_hd__o211a_1 _1112_ (.A1(\MOS6502.AXYS[3][7] ),
    .A2(_0327_),
    .B1(_0329_),
    .C1(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__a221oi_4 _1113_ (.A1(\MOS6502.AXYS[0][7] ),
    .A2(_0332_),
    .B1(_0333_),
    .B2(\MOS6502.AXYS[1][7] ),
    .C1(_0496_),
    .Y(_0497_));
 sky130_fd_sc_hd__nor2_1 _1114_ (.A(_0310_),
    .B(_0497_),
    .Y(_0498_));
 sky130_fd_sc_hd__a22o_2 _1115_ (.A1(net8),
    .A2(_0337_),
    .B1(net54),
    .B2(\MOS6502.ABH[7] ),
    .X(_0499_));
 sky130_fd_sc_hd__a211o_4 _1116_ (.A1(\MOS6502.ADD[7] ),
    .A2(_0344_),
    .B1(_0498_),
    .C1(_0499_),
    .X(\MOS6502.AI[7] ));
 sky130_fd_sc_hd__a22o_2 _1117_ (.A1(\MOS6502.PC[6] ),
    .A2(_0336_),
    .B1(_0361_),
    .B2(net7),
    .X(_0500_));
 sky130_fd_sc_hd__and2b_1 _1118_ (.A_N(_0346_),
    .B(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _1119_ (.A0(net42),
    .A1(_0367_),
    .S(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__a21bo_1 _1120_ (.A1(net42),
    .A2(_0500_),
    .B1_N(_0346_),
    .X(_0503_));
 sky130_fd_sc_hd__o211a_1 _1121_ (.A1(_0372_),
    .A2(_0502_),
    .B1(_0503_),
    .C1(_0290_),
    .X(_0504_));
 sky130_fd_sc_hd__a21oi_1 _1122_ (.A1(_0289_),
    .A2(\MOS6502.AI[7] ),
    .B1(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__mux2_1 _1123_ (.A0(_0379_),
    .A1(_0375_),
    .S(_0500_),
    .X(_0506_));
 sky130_fd_sc_hd__or3_2 _1124_ (.A(_0381_),
    .B(_0505_),
    .C(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__or2_1 _1125_ (.A(_0377_),
    .B(_0506_),
    .X(_0508_));
 sky130_fd_sc_hd__a21bo_1 _1126_ (.A1(_0505_),
    .A2(_0508_),
    .B1_N(_0507_),
    .X(_0509_));
 sky130_fd_sc_hd__a21o_1 _1127_ (.A1(_0383_),
    .A2(_0494_),
    .B1(_0509_),
    .X(_0510_));
 sky130_fd_sc_hd__nand3_1 _1128_ (.A(_0383_),
    .B(_0494_),
    .C(_0509_),
    .Y(_0511_));
 sky130_fd_sc_hd__and2_1 _1129_ (.A(_0510_),
    .B(_0511_),
    .X(\MOS6502.ALU.temp[6] ));
 sky130_fd_sc_hd__a22o_2 _1130_ (.A1(\MOS6502.PC[7] ),
    .A2(_0336_),
    .B1(_0361_),
    .B2(net8),
    .X(_0512_));
 sky130_fd_sc_hd__a21oi_1 _1131_ (.A1(net42),
    .A2(_0512_),
    .B1(\MOS6502.AI[7] ),
    .Y(_0513_));
 sky130_fd_sc_hd__o21ai_1 _1132_ (.A1(_0369_),
    .A2(_0512_),
    .B1(_0290_),
    .Y(_0514_));
 sky130_fd_sc_hd__a31o_1 _1133_ (.A1(_0370_),
    .A2(\MOS6502.AI[7] ),
    .A3(_0512_),
    .B1(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__o2bb2a_1 _1134_ (.A1_N(_0289_),
    .A2_N(_0477_),
    .B1(_0513_),
    .B2(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _1135_ (.A0(_0396_),
    .A1(_0375_),
    .S(_0512_),
    .X(_0517_));
 sky130_fd_sc_hd__a21oi_1 _1136_ (.A1(_0377_),
    .A2(_0516_),
    .B1(_0517_),
    .Y(\MOS6502.ALU.temp_BI[7] ));
 sky130_fd_sc_hd__or2_1 _1137_ (.A(_0516_),
    .B(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__o21ai_1 _1138_ (.A1(_0377_),
    .A2(_0517_),
    .B1(_0516_),
    .Y(_0519_));
 sky130_fd_sc_hd__nand2_1 _1139_ (.A(_0518_),
    .B(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__a21o_1 _1140_ (.A1(_0507_),
    .A2(_0510_),
    .B1(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__nand3_1 _1141_ (.A(_0507_),
    .B(_0510_),
    .C(_0520_),
    .Y(_0522_));
 sky130_fd_sc_hd__and2_1 _1142_ (.A(_0521_),
    .B(_0522_),
    .X(\MOS6502.ALU.temp[7] ));
 sky130_fd_sc_hd__a211o_1 _1143_ (.A1(_0383_),
    .A2(_0493_),
    .B1(_0492_),
    .C1(_0399_),
    .X(_0523_));
 sky130_fd_sc_hd__and2_1 _1144_ (.A(_0494_),
    .B(_0523_),
    .X(\MOS6502.ALU.temp[5] ));
 sky130_fd_sc_hd__a211o_1 _1145_ (.A1(_0518_),
    .A2(_0521_),
    .B1(net46),
    .C1(_0459_),
    .X(_0524_));
 sky130_fd_sc_hd__o211ai_1 _1146_ (.A1(net46),
    .A2(_0459_),
    .B1(_0518_),
    .C1(_0521_),
    .Y(_0525_));
 sky130_fd_sc_hd__o2111a_1 _1147_ (.A1(\MOS6502.ALU.temp[6] ),
    .A2(\MOS6502.ALU.temp[5] ),
    .B1(_0521_),
    .C1(_0490_),
    .D1(_0522_),
    .X(_0526_));
 sky130_fd_sc_hd__a21o_1 _1148_ (.A1(_0524_),
    .A2(_0525_),
    .B1(_0526_),
    .X(_0001_));
 sky130_fd_sc_hd__and2_1 _1149_ (.A(\MOS6502.D ),
    .B(\MOS6502.adc_sbc ),
    .X(_0000_));
 sky130_fd_sc_hd__xnor2_1 _1150_ (.A(_0466_),
    .B(_0479_),
    .Y(\MOS6502.ALU.temp[0] ));
 sky130_fd_sc_hd__nor2_1 _1151_ (.A(_0281_),
    .B(_0319_),
    .Y(_0527_));
 sky130_fd_sc_hd__or2_1 _1152_ (.A(_0281_),
    .B(_0319_),
    .X(_0528_));
 sky130_fd_sc_hd__nor2_2 _1153_ (.A(_0244_),
    .B(_0319_),
    .Y(_0529_));
 sky130_fd_sc_hd__nor2_4 _1154_ (.A(\MOS6502.state[5] ),
    .B(_0341_),
    .Y(_0530_));
 sky130_fd_sc_hd__a211o_4 _1155_ (.A1(net81),
    .A2(_0530_),
    .B1(_0529_),
    .C1(_0527_),
    .X(_0531_));
 sky130_fd_sc_hd__or2_2 _1156_ (.A(net54),
    .B(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__nand2_8 _1157_ (.A(net71),
    .B(net64),
    .Y(_0533_));
 sky130_fd_sc_hd__o31ai_4 _1158_ (.A1(net69),
    .A2(net64),
    .A3(net43),
    .B1(_0533_),
    .Y(_0534_));
 sky130_fd_sc_hd__nor2_8 _1159_ (.A(net71),
    .B(net60),
    .Y(_0535_));
 sky130_fd_sc_hd__a22o_1 _1160_ (.A1(\MOS6502.ADD[0] ),
    .A2(net43),
    .B1(_0535_),
    .B2(\MOS6502.ABL[0] ),
    .X(_0536_));
 sky130_fd_sc_hd__a21oi_2 _1161_ (.A1(\MOS6502.PC[0] ),
    .A2(_0534_),
    .B1(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__or3_1 _1162_ (.A(net88),
    .B(net84),
    .C(net82),
    .X(_0538_));
 sky130_fd_sc_hd__nor2_1 _1163_ (.A(_0529_),
    .B(_0530_),
    .Y(_0539_));
 sky130_fd_sc_hd__xnor2_1 _1164_ (.A(\MOS6502.backwards ),
    .B(\MOS6502.ALU.CO ),
    .Y(_0540_));
 sky130_fd_sc_hd__nand2_1 _1165_ (.A(net53),
    .B(_0540_),
    .Y(_0541_));
 sky130_fd_sc_hd__and3_1 _1166_ (.A(_0240_),
    .B(_0292_),
    .C(_0538_),
    .X(_0542_));
 sky130_fd_sc_hd__o211a_1 _1167_ (.A1(net75),
    .A2(_0542_),
    .B1(_0541_),
    .C1(_0533_),
    .X(_0543_));
 sky130_fd_sc_hd__o211a_1 _1168_ (.A1(net80),
    .A2(_0281_),
    .B1(_0539_),
    .C1(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__or2_1 _1169_ (.A(_0537_),
    .B(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__xor2_1 _1170_ (.A(_0537_),
    .B(_0544_),
    .X(_0002_));
 sky130_fd_sc_hd__a2bb2o_1 _1171_ (.A1_N(\MOS6502.res ),
    .A2_N(_0249_),
    .B1(net43),
    .B2(\MOS6502.ADD[1] ),
    .X(_0546_));
 sky130_fd_sc_hd__nor2_8 _1172_ (.A(_0242_),
    .B(_0341_),
    .Y(_0547_));
 sky130_fd_sc_hd__or4_2 _1173_ (.A(net68),
    .B(net64),
    .C(net43),
    .D(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__a221o_1 _1174_ (.A1(\MOS6502.PC[1] ),
    .A2(_0534_),
    .B1(_0535_),
    .B2(\MOS6502.ABL[1] ),
    .C1(_0546_),
    .X(_0549_));
 sky130_fd_sc_hd__and2b_1 _1175_ (.A_N(_0545_),
    .B(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__and2b_1 _1176_ (.A_N(_0549_),
    .B(_0545_),
    .X(_0551_));
 sky130_fd_sc_hd__nor2_1 _1177_ (.A(_0550_),
    .B(_0551_),
    .Y(_0009_));
 sky130_fd_sc_hd__o21a_2 _1178_ (.A1(_0221_),
    .A2(\MOS6502.res ),
    .B1(net68),
    .X(_0552_));
 sky130_fd_sc_hd__a22o_1 _1179_ (.A1(\MOS6502.ADD[2] ),
    .A2(net43),
    .B1(_0534_),
    .B2(\MOS6502.PC[2] ),
    .X(_0553_));
 sky130_fd_sc_hd__a211oi_4 _1180_ (.A1(\MOS6502.ABL[2] ),
    .A2(_0535_),
    .B1(_0552_),
    .C1(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__or3b_2 _1181_ (.A(_0554_),
    .B(_0545_),
    .C_N(_0549_),
    .X(_0555_));
 sky130_fd_sc_hd__xnor2_1 _1182_ (.A(_0550_),
    .B(_0554_),
    .Y(_0010_));
 sky130_fd_sc_hd__o21ai_4 _1183_ (.A1(net64),
    .A2(net43),
    .B1(_0533_),
    .Y(_0556_));
 sky130_fd_sc_hd__a221o_1 _1184_ (.A1(\MOS6502.ADD[3] ),
    .A2(net43),
    .B1(_0535_),
    .B2(\MOS6502.ABL[3] ),
    .C1(net69),
    .X(_0557_));
 sky130_fd_sc_hd__a21oi_1 _1185_ (.A1(\MOS6502.PC[3] ),
    .A2(_0556_),
    .B1(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__or2_1 _1186_ (.A(_0555_),
    .B(_0558_),
    .X(_0559_));
 sky130_fd_sc_hd__xor2_1 _1187_ (.A(_0555_),
    .B(_0558_),
    .X(_0011_));
 sky130_fd_sc_hd__a221o_1 _1188_ (.A1(\MOS6502.ADD[4] ),
    .A2(net43),
    .B1(_0535_),
    .B2(\MOS6502.ABL[4] ),
    .C1(net69),
    .X(_0560_));
 sky130_fd_sc_hd__a21oi_1 _1189_ (.A1(\MOS6502.PC[4] ),
    .A2(_0556_),
    .B1(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__or2_1 _1190_ (.A(_0559_),
    .B(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__xor2_1 _1191_ (.A(_0559_),
    .B(_0561_),
    .X(_0012_));
 sky130_fd_sc_hd__a221o_1 _1192_ (.A1(\MOS6502.ADD[5] ),
    .A2(net43),
    .B1(_0535_),
    .B2(\MOS6502.ABL[5] ),
    .C1(net69),
    .X(_0563_));
 sky130_fd_sc_hd__a21oi_1 _1193_ (.A1(\MOS6502.PC[5] ),
    .A2(_0556_),
    .B1(_0563_),
    .Y(_0564_));
 sky130_fd_sc_hd__or2_1 _1194_ (.A(_0562_),
    .B(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__xor2_1 _1195_ (.A(_0562_),
    .B(_0564_),
    .X(_0013_));
 sky130_fd_sc_hd__a221o_1 _1196_ (.A1(\MOS6502.ADD[6] ),
    .A2(_0532_),
    .B1(_0535_),
    .B2(\MOS6502.ABL[6] ),
    .C1(net69),
    .X(_0566_));
 sky130_fd_sc_hd__a21oi_1 _1197_ (.A1(\MOS6502.PC[6] ),
    .A2(_0556_),
    .B1(_0566_),
    .Y(_0567_));
 sky130_fd_sc_hd__or2_1 _1198_ (.A(_0565_),
    .B(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__xor2_1 _1199_ (.A(_0565_),
    .B(_0567_),
    .X(_0014_));
 sky130_fd_sc_hd__a221o_1 _1200_ (.A1(\MOS6502.ADD[7] ),
    .A2(net43),
    .B1(_0535_),
    .B2(\MOS6502.ABL[7] ),
    .C1(net69),
    .X(_0569_));
 sky130_fd_sc_hd__a21oi_2 _1201_ (.A1(\MOS6502.PC[7] ),
    .A2(_0556_),
    .B1(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__nor2_2 _1202_ (.A(_0568_),
    .B(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__and2_1 _1203_ (.A(_0568_),
    .B(_0570_),
    .X(_0572_));
 sky130_fd_sc_hd__nor2_1 _1204_ (.A(_0571_),
    .B(_0572_),
    .Y(_0015_));
 sky130_fd_sc_hd__nand2_4 _1205_ (.A(_0533_),
    .B(_0548_),
    .Y(_0573_));
 sky130_fd_sc_hd__or2_4 _1206_ (.A(net54),
    .B(_0535_),
    .X(_0574_));
 sky130_fd_sc_hd__a221o_1 _1207_ (.A1(\MOS6502.ADD[0] ),
    .A2(_0547_),
    .B1(_0574_),
    .B2(\MOS6502.ABH[0] ),
    .C1(net68),
    .X(_0575_));
 sky130_fd_sc_hd__a221o_2 _1208_ (.A1(net1),
    .A2(_0531_),
    .B1(_0573_),
    .B2(\MOS6502.PC[8] ),
    .C1(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__xor2_1 _1209_ (.A(_0571_),
    .B(_0576_),
    .X(_0016_));
 sky130_fd_sc_hd__a221o_1 _1210_ (.A1(\MOS6502.ADD[1] ),
    .A2(_0547_),
    .B1(_0574_),
    .B2(\MOS6502.ABH[1] ),
    .C1(net68),
    .X(_0577_));
 sky130_fd_sc_hd__a221o_1 _1211_ (.A1(net2),
    .A2(_0531_),
    .B1(_0573_),
    .B2(\MOS6502.PC[9] ),
    .C1(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__and3_2 _1212_ (.A(_0571_),
    .B(_0576_),
    .C(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__a21oi_1 _1213_ (.A1(_0571_),
    .A2(_0576_),
    .B1(_0578_),
    .Y(_0580_));
 sky130_fd_sc_hd__nor2_1 _1214_ (.A(_0579_),
    .B(_0580_),
    .Y(_0017_));
 sky130_fd_sc_hd__a221o_1 _1215_ (.A1(\MOS6502.ADD[2] ),
    .A2(_0547_),
    .B1(_0574_),
    .B2(\MOS6502.ABH[2] ),
    .C1(net68),
    .X(_0581_));
 sky130_fd_sc_hd__a221o_2 _1216_ (.A1(net3),
    .A2(_0531_),
    .B1(_0573_),
    .B2(\MOS6502.PC[10] ),
    .C1(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__xor2_1 _1217_ (.A(_0579_),
    .B(_0582_),
    .X(_0003_));
 sky130_fd_sc_hd__a221o_1 _1218_ (.A1(\MOS6502.ADD[3] ),
    .A2(_0547_),
    .B1(_0574_),
    .B2(\MOS6502.ABH[3] ),
    .C1(net68),
    .X(_0583_));
 sky130_fd_sc_hd__a221o_1 _1219_ (.A1(net4),
    .A2(_0531_),
    .B1(_0573_),
    .B2(\MOS6502.PC[11] ),
    .C1(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__and3_2 _1220_ (.A(_0579_),
    .B(_0582_),
    .C(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__a21oi_1 _1221_ (.A1(_0579_),
    .A2(_0582_),
    .B1(_0584_),
    .Y(_0586_));
 sky130_fd_sc_hd__nor2_1 _1222_ (.A(_0585_),
    .B(_0586_),
    .Y(_0004_));
 sky130_fd_sc_hd__a221o_1 _1223_ (.A1(\MOS6502.ADD[4] ),
    .A2(_0547_),
    .B1(_0574_),
    .B2(\MOS6502.ABH[4] ),
    .C1(net68),
    .X(_0587_));
 sky130_fd_sc_hd__a221o_2 _1224_ (.A1(net5),
    .A2(_0531_),
    .B1(_0573_),
    .B2(\MOS6502.PC[12] ),
    .C1(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__xor2_1 _1225_ (.A(_0585_),
    .B(_0588_),
    .X(_0005_));
 sky130_fd_sc_hd__a221o_1 _1226_ (.A1(\MOS6502.ADD[5] ),
    .A2(_0547_),
    .B1(_0574_),
    .B2(\MOS6502.ABH[5] ),
    .C1(net68),
    .X(_0589_));
 sky130_fd_sc_hd__a221o_1 _1227_ (.A1(net6),
    .A2(_0531_),
    .B1(_0573_),
    .B2(\MOS6502.PC[13] ),
    .C1(_0589_),
    .X(_0590_));
 sky130_fd_sc_hd__and3_1 _1228_ (.A(_0585_),
    .B(_0588_),
    .C(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__a21oi_1 _1229_ (.A1(_0585_),
    .A2(_0588_),
    .B1(_0590_),
    .Y(_0592_));
 sky130_fd_sc_hd__nor2_1 _1230_ (.A(_0591_),
    .B(_0592_),
    .Y(_0006_));
 sky130_fd_sc_hd__a221o_1 _1231_ (.A1(\MOS6502.ADD[6] ),
    .A2(_0547_),
    .B1(_0574_),
    .B2(\MOS6502.ABH[6] ),
    .C1(net68),
    .X(_0593_));
 sky130_fd_sc_hd__a221o_1 _1232_ (.A1(net7),
    .A2(_0531_),
    .B1(_0573_),
    .B2(\MOS6502.PC[14] ),
    .C1(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__nand2_1 _1233_ (.A(_0591_),
    .B(_0594_),
    .Y(_0595_));
 sky130_fd_sc_hd__or2_1 _1234_ (.A(_0591_),
    .B(_0594_),
    .X(_0596_));
 sky130_fd_sc_hd__and2_1 _1235_ (.A(_0595_),
    .B(_0596_),
    .X(_0007_));
 sky130_fd_sc_hd__a221o_1 _1236_ (.A1(\MOS6502.ADD[7] ),
    .A2(_0547_),
    .B1(_0574_),
    .B2(\MOS6502.ABH[7] ),
    .C1(net69),
    .X(_0597_));
 sky130_fd_sc_hd__a221o_1 _1237_ (.A1(net8),
    .A2(_0531_),
    .B1(_0573_),
    .B2(\MOS6502.PC[15] ),
    .C1(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__xnor2_1 _1238_ (.A(_0595_),
    .B(_0598_),
    .Y(_0008_));
 sky130_fd_sc_hd__and3_1 _1239_ (.A(_0401_),
    .B(_0488_),
    .C(_0491_),
    .X(_0599_));
 sky130_fd_sc_hd__nor2_1 _1240_ (.A(_0492_),
    .B(_0599_),
    .Y(\MOS6502.ALU.temp[4] ));
 sky130_fd_sc_hd__and2b_1 _1241_ (.A_N(_0487_),
    .B(_0489_),
    .X(\MOS6502.ALU.temp[3] ));
 sky130_fd_sc_hd__mux2_1 _1242_ (.A0(net5),
    .A1(\MOS6502.IRHOLD[4] ),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0600_));
 sky130_fd_sc_hd__and2_4 _1243_ (.A(net70),
    .B(net72),
    .X(_0601_));
 sky130_fd_sc_hd__nand2_1 _1244_ (.A(net70),
    .B(net72),
    .Y(_0602_));
 sky130_fd_sc_hd__mux2_2 _1245_ (.A0(net4),
    .A1(\MOS6502.IRHOLD[3] ),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0603_));
 sky130_fd_sc_hd__nand2_4 _1246_ (.A(net70),
    .B(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hd__mux2_4 _1247_ (.A0(net3),
    .A1(\MOS6502.IRHOLD[2] ),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _1248_ (.A0(net2),
    .A1(\MOS6502.IRHOLD[1] ),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0606_));
 sky130_fd_sc_hd__mux2_1 _1249_ (.A0(net1),
    .A1(\MOS6502.IRHOLD[0] ),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0607_));
 sky130_fd_sc_hd__and2_4 _1250_ (.A(net70),
    .B(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__and2_1 _1251_ (.A(net70),
    .B(_0606_),
    .X(_0609_));
 sky130_fd_sc_hd__nand2_2 _1252_ (.A(net70),
    .B(_0606_),
    .Y(_0610_));
 sky130_fd_sc_hd__and2_4 _1253_ (.A(_0608_),
    .B(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__nand2_4 _1254_ (.A(_0608_),
    .B(_0610_),
    .Y(_0612_));
 sky130_fd_sc_hd__and2_1 _1255_ (.A(net70),
    .B(_0605_),
    .X(_0613_));
 sky130_fd_sc_hd__nand2_8 _1256_ (.A(net70),
    .B(_0605_),
    .Y(_0614_));
 sky130_fd_sc_hd__or2_4 _1257_ (.A(_0604_),
    .B(_0613_),
    .X(_0615_));
 sky130_fd_sc_hd__nand2_2 _1258_ (.A(_0604_),
    .B(_0614_),
    .Y(_0616_));
 sky130_fd_sc_hd__or4_1 _1259_ (.A(_0232_),
    .B(net72),
    .C(_0608_),
    .D(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__o31a_2 _1260_ (.A1(_0601_),
    .A2(_0612_),
    .A3(_0615_),
    .B1(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__or3_1 _1261_ (.A(\MOS6502.ALU.CO ),
    .B(\MOS6502.write_back ),
    .C(\MOS6502.store ),
    .X(_0619_));
 sky130_fd_sc_hd__o32a_1 _1262_ (.A1(\MOS6502.write_back ),
    .A2(net76),
    .A3(_0284_),
    .B1(_0268_),
    .B2(net77),
    .X(_0620_));
 sky130_fd_sc_hd__o211a_1 _1263_ (.A1(net78),
    .A2(_0278_),
    .B1(_0528_),
    .C1(_0263_),
    .X(_0621_));
 sky130_fd_sc_hd__o221a_1 _1264_ (.A1(\MOS6502.write_back ),
    .A2(_0277_),
    .B1(net58),
    .B2(_0618_),
    .C1(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__o31ai_1 _1265_ (.A1(\MOS6502.ALU.CO ),
    .A2(\MOS6502.store ),
    .A3(_0620_),
    .B1(_0622_),
    .Y(_0623_));
 sky130_fd_sc_hd__o21a_1 _1266_ (.A1(\MOS6502.ALU.CO ),
    .A2(\MOS6502.store ),
    .B1(_0471_),
    .X(_0624_));
 sky130_fd_sc_hd__or2_2 _1267_ (.A(_0608_),
    .B(_0609_),
    .X(_0625_));
 sky130_fd_sc_hd__or2_4 _1268_ (.A(_0616_),
    .B(net47),
    .X(_0626_));
 sky130_fd_sc_hd__nand2_2 _1269_ (.A(_0234_),
    .B(net50),
    .Y(_0627_));
 sky130_fd_sc_hd__or2_2 _1270_ (.A(_0231_),
    .B(_0236_),
    .X(_0628_));
 sky130_fd_sc_hd__or3_1 _1271_ (.A(_0626_),
    .B(_0627_),
    .C(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__nor2_1 _1272_ (.A(net58),
    .B(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__or3_1 _1273_ (.A(_0623_),
    .B(_0624_),
    .C(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__nand2_1 _1274_ (.A(_0232_),
    .B(net50),
    .Y(_0632_));
 sky130_fd_sc_hd__nor2_1 _1275_ (.A(\MOS6502.IR[7] ),
    .B(_0627_),
    .Y(_0633_));
 sky130_fd_sc_hd__nor2_1 _1276_ (.A(_0608_),
    .B(_0615_),
    .Y(_0634_));
 sky130_fd_sc_hd__nor2_4 _1277_ (.A(_0615_),
    .B(_0625_),
    .Y(_0635_));
 sky130_fd_sc_hd__nand2_1 _1278_ (.A(net61),
    .B(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__and3_2 _1279_ (.A(net62),
    .B(_0633_),
    .C(_0635_),
    .X(_0637_));
 sky130_fd_sc_hd__or4_2 _1280_ (.A(net59),
    .B(_0601_),
    .C(_0603_),
    .D(_0614_),
    .X(_0638_));
 sky130_fd_sc_hd__o21ai_1 _1281_ (.A1(net76),
    .A2(_0264_),
    .B1(_0638_),
    .Y(_0639_));
 sky130_fd_sc_hd__nor2_1 _1282_ (.A(_0319_),
    .B(_0338_),
    .Y(_0640_));
 sky130_fd_sc_hd__and2b_1 _1283_ (.A_N(_0540_),
    .B(net53),
    .X(_0641_));
 sky130_fd_sc_hd__and2_1 _1284_ (.A(\MOS6502.write_back ),
    .B(_0276_),
    .X(_0642_));
 sky130_fd_sc_hd__or2_1 _1285_ (.A(_0639_),
    .B(_0640_),
    .X(_0643_));
 sky130_fd_sc_hd__or4_1 _1286_ (.A(_0312_),
    .B(_0357_),
    .C(_0474_),
    .D(_0641_),
    .X(_0644_));
 sky130_fd_sc_hd__or3_1 _1287_ (.A(_0642_),
    .B(_0643_),
    .C(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__or3_1 _1288_ (.A(net59),
    .B(net50),
    .C(_0626_),
    .X(_0646_));
 sky130_fd_sc_hd__a2bb2o_1 _1289_ (.A1_N(_0256_),
    .A2_N(_0272_),
    .B1(_0305_),
    .B2(net73),
    .X(_0647_));
 sky130_fd_sc_hd__or4b_1 _1290_ (.A(_0297_),
    .B(_0645_),
    .C(_0647_),
    .D_N(_0646_),
    .X(_0648_));
 sky130_fd_sc_hd__nand2_1 _1291_ (.A(_0633_),
    .B(_0635_),
    .Y(_0649_));
 sky130_fd_sc_hd__or3_1 _1292_ (.A(_0631_),
    .B(_0637_),
    .C(_0648_),
    .X(_0018_));
 sky130_fd_sc_hd__or2_2 _1293_ (.A(_0234_),
    .B(net72),
    .X(_0650_));
 sky130_fd_sc_hd__or4_2 _1294_ (.A(\MOS6502.IR[7] ),
    .B(_0615_),
    .C(net47),
    .D(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__nor2_1 _1295_ (.A(net58),
    .B(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__or4_1 _1296_ (.A(net59),
    .B(_0601_),
    .C(_0612_),
    .D(_0616_),
    .X(_0653_));
 sky130_fd_sc_hd__or3b_1 _1297_ (.A(_0285_),
    .B(_0652_),
    .C_N(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__nor2_1 _1298_ (.A(net77),
    .B(_0244_),
    .Y(_0655_));
 sky130_fd_sc_hd__or2_1 _1299_ (.A(_0608_),
    .B(_0614_),
    .X(_0656_));
 sky130_fd_sc_hd__inv_2 _1300_ (.A(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__or2_2 _1301_ (.A(_0604_),
    .B(_0614_),
    .X(_0658_));
 sky130_fd_sc_hd__or4_1 _1302_ (.A(net47),
    .B(_0627_),
    .C(_0628_),
    .D(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__nor2_1 _1303_ (.A(net58),
    .B(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__or4_1 _1304_ (.A(_0318_),
    .B(_0654_),
    .C(_0655_),
    .D(_0660_),
    .X(_0661_));
 sky130_fd_sc_hd__nand2_2 _1305_ (.A(_0232_),
    .B(_0236_),
    .Y(_0662_));
 sky130_fd_sc_hd__or2_4 _1306_ (.A(_0650_),
    .B(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__or2_2 _1307_ (.A(_0628_),
    .B(_0650_),
    .X(_0664_));
 sky130_fd_sc_hd__or2_1 _1308_ (.A(_0626_),
    .B(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__a211o_1 _1309_ (.A1(_0663_),
    .A2(_0664_),
    .B1(net59),
    .C1(_0626_),
    .X(_0666_));
 sky130_fd_sc_hd__a21o_1 _1310_ (.A1(_0612_),
    .A2(_0614_),
    .B1(_0604_),
    .X(_0667_));
 sky130_fd_sc_hd__mux4_2 _1311_ (.A0(\MOS6502.N ),
    .A1(\MOS6502.V ),
    .A2(\MOS6502.C ),
    .A3(\MOS6502.Z ),
    .S0(\MOS6502.cond_code[1] ),
    .S1(\MOS6502.cond_code[2] ),
    .X(_0668_));
 sky130_fd_sc_hd__xnor2_2 _1312_ (.A(\MOS6502.cond_code[0] ),
    .B(_0668_),
    .Y(_0669_));
 sky130_fd_sc_hd__a21o_1 _1313_ (.A1(_0336_),
    .A2(_0669_),
    .B1(_0293_),
    .X(_0670_));
 sky130_fd_sc_hd__or4_2 _1314_ (.A(net59),
    .B(net50),
    .C(_0612_),
    .D(_0616_),
    .X(_0671_));
 sky130_fd_sc_hd__o211a_1 _1315_ (.A1(net85),
    .A2(_0291_),
    .B1(_0671_),
    .C1(_0245_),
    .X(_0672_));
 sky130_fd_sc_hd__nor3b_1 _1316_ (.A(_0661_),
    .B(_0670_),
    .C_N(_0666_),
    .Y(_0673_));
 sky130_fd_sc_hd__o31a_1 _1317_ (.A1(net58),
    .A2(net50),
    .A3(_0667_),
    .B1(_0672_),
    .X(_0674_));
 sky130_fd_sc_hd__nand3b_1 _1318_ (.A_N(_0645_),
    .B(_0673_),
    .C(_0674_),
    .Y(_0019_));
 sky130_fd_sc_hd__o21ai_1 _1319_ (.A1(_0611_),
    .A2(_0613_),
    .B1(_0604_),
    .Y(_0675_));
 sky130_fd_sc_hd__or3_1 _1320_ (.A(net47),
    .B(_0658_),
    .C(_0664_),
    .X(_0676_));
 sky130_fd_sc_hd__o21a_1 _1321_ (.A1(_0232_),
    .A2(net72),
    .B1(_0663_),
    .X(_0677_));
 sky130_fd_sc_hd__nor2_2 _1322_ (.A(_0608_),
    .B(_0610_),
    .Y(_0678_));
 sky130_fd_sc_hd__or2_2 _1323_ (.A(_0608_),
    .B(_0610_),
    .X(_0679_));
 sky130_fd_sc_hd__a211o_1 _1324_ (.A1(_0612_),
    .A2(_0679_),
    .B1(_0658_),
    .C1(_0601_),
    .X(_0680_));
 sky130_fd_sc_hd__o31a_1 _1325_ (.A1(net47),
    .A2(_0658_),
    .A3(_0677_),
    .B1(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__or2_2 _1326_ (.A(_0615_),
    .B(_0679_),
    .X(_0682_));
 sky130_fd_sc_hd__o31a_1 _1327_ (.A1(\MOS6502.IR[7] ),
    .A2(_0600_),
    .A3(_0609_),
    .B1(_0634_),
    .X(_0683_));
 sky130_fd_sc_hd__and3b_1 _1328_ (.A_N(_0683_),
    .B(_0649_),
    .C(_0629_),
    .X(_0684_));
 sky130_fd_sc_hd__o2111a_1 _1329_ (.A1(_0626_),
    .A2(_0663_),
    .B1(_0676_),
    .C1(_0651_),
    .D1(_0659_),
    .X(_0685_));
 sky130_fd_sc_hd__o21a_1 _1330_ (.A1(_0627_),
    .A2(_0662_),
    .B1(_0664_),
    .X(_0686_));
 sky130_fd_sc_hd__o2111a_1 _1331_ (.A1(net50),
    .A2(_0626_),
    .B1(_0675_),
    .C1(_0618_),
    .D1(net62),
    .X(_0687_));
 sky130_fd_sc_hd__o221a_1 _1332_ (.A1(_0602_),
    .A2(_0667_),
    .B1(_0686_),
    .B2(_0626_),
    .C1(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__and4_1 _1333_ (.A(_0681_),
    .B(_0684_),
    .C(_0685_),
    .D(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__a31o_1 _1334_ (.A1(_0244_),
    .A2(_0268_),
    .A3(_0538_),
    .B1(net74),
    .X(_0690_));
 sky130_fd_sc_hd__o311a_1 _1335_ (.A1(net75),
    .A2(_0292_),
    .A3(_0669_),
    .B1(_0541_),
    .C1(_0283_),
    .X(_0691_));
 sky130_fd_sc_hd__or4bb_2 _1336_ (.A(_0530_),
    .B(_0689_),
    .C_N(_0690_),
    .D_N(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__a211o_1 _1337_ (.A1(_0239_),
    .A2(_0320_),
    .B1(_0692_),
    .C1(_0302_),
    .X(_0693_));
 sky130_fd_sc_hd__a22o_1 _1338_ (.A1(_0470_),
    .A2(_0619_),
    .B1(_0683_),
    .B2(net62),
    .X(_0694_));
 sky130_fd_sc_hd__or4b_1 _1339_ (.A(_0296_),
    .B(_0641_),
    .C(_0643_),
    .D_N(_0646_),
    .X(_0695_));
 sky130_fd_sc_hd__or4_1 _1340_ (.A(_0631_),
    .B(_0670_),
    .C(_0694_),
    .D(_0695_),
    .X(_0696_));
 sky130_fd_sc_hd__or3_1 _1341_ (.A(_0661_),
    .B(_0693_),
    .C(_0696_),
    .X(_0020_));
 sky130_fd_sc_hd__nor2_1 _1342_ (.A(net58),
    .B(_0681_),
    .Y(_0697_));
 sky130_fd_sc_hd__o21ai_1 _1343_ (.A1(net58),
    .A2(_0676_),
    .B1(_0355_),
    .Y(_0698_));
 sky130_fd_sc_hd__or4_2 _1344_ (.A(net59),
    .B(_0602_),
    .C(_0603_),
    .D(_0614_),
    .X(_0699_));
 sky130_fd_sc_hd__nand2_1 _1345_ (.A(_0340_),
    .B(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hd__nand2_1 _1346_ (.A(_0317_),
    .B(_0674_),
    .Y(_0701_));
 sky130_fd_sc_hd__or4_1 _1347_ (.A(_0694_),
    .B(_0698_),
    .C(_0700_),
    .D(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__or4b_1 _1348_ (.A(_0018_),
    .B(_0697_),
    .C(_0702_),
    .D_N(_0673_),
    .X(_0703_));
 sky130_fd_sc_hd__nor2_1 _1349_ (.A(_0693_),
    .B(_0703_),
    .Y(_0704_));
 sky130_fd_sc_hd__o21ai_1 _1350_ (.A1(_0256_),
    .A2(_0272_),
    .B1(_0245_),
    .Y(_0705_));
 sky130_fd_sc_hd__or4_1 _1351_ (.A(_0296_),
    .B(_0358_),
    .C(_0639_),
    .D(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__or4_1 _1352_ (.A(_0623_),
    .B(_0654_),
    .C(_0698_),
    .D(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__or4b_1 _1353_ (.A(_0692_),
    .B(_0704_),
    .C(_0707_),
    .D_N(_0666_),
    .X(_0021_));
 sky130_fd_sc_hd__o211a_1 _1354_ (.A1(net85),
    .A2(_0238_),
    .B1(_0256_),
    .C1(_0338_),
    .X(_0708_));
 sky130_fd_sc_hd__a2bb2o_1 _1355_ (.A1_N(net77),
    .A2_N(_0708_),
    .B1(_0305_),
    .B2(net81),
    .X(_0709_));
 sky130_fd_sc_hd__nor3_4 _1356_ (.A(net67),
    .B(_0297_),
    .C(_0318_),
    .Y(_0710_));
 sky130_fd_sc_hd__nand2_1 _1357_ (.A(_0671_),
    .B(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__or4_1 _1358_ (.A(_0474_),
    .B(_0624_),
    .C(_0655_),
    .D(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__nor2_1 _1359_ (.A(net58),
    .B(_0685_),
    .Y(_0713_));
 sky130_fd_sc_hd__or4_1 _1360_ (.A(_0700_),
    .B(_0709_),
    .C(_0712_),
    .D(_0713_),
    .X(_0022_));
 sky130_fd_sc_hd__a21oi_1 _1361_ (.A1(_0665_),
    .A2(_0684_),
    .B1(net58),
    .Y(_0714_));
 sky130_fd_sc_hd__o41a_2 _1362_ (.A1(net86),
    .A2(net88),
    .A3(_0223_),
    .A4(net74),
    .B1(_0317_),
    .X(_0715_));
 sky130_fd_sc_hd__nand2_1 _1363_ (.A(_0342_),
    .B(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__nand2_1 _1364_ (.A(_0638_),
    .B(_0699_),
    .Y(_0717_));
 sky130_fd_sc_hd__a31o_1 _1365_ (.A1(_0247_),
    .A2(_0278_),
    .A3(_0284_),
    .B1(net73),
    .X(_0718_));
 sky130_fd_sc_hd__or4b_1 _1366_ (.A(_0306_),
    .B(_0642_),
    .C(_0717_),
    .D_N(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__or3_1 _1367_ (.A(_0714_),
    .B(_0716_),
    .C(_0719_),
    .X(_0023_));
 sky130_fd_sc_hd__nor3_4 _1368_ (.A(_0253_),
    .B(net51),
    .C(_0294_),
    .Y(_0720_));
 sky130_fd_sc_hd__or3_4 _1369_ (.A(_0253_),
    .B(net51),
    .C(_0294_),
    .X(_0721_));
 sky130_fd_sc_hd__a211oi_4 _1370_ (.A1(net81),
    .A2(_0530_),
    .B1(_0529_),
    .C1(_0472_),
    .Y(_0722_));
 sky130_fd_sc_hd__o21ai_4 _1371_ (.A1(\MOS6502.state[5] ),
    .A2(_0270_),
    .B1(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__or3_1 _1372_ (.A(net48),
    .B(net68),
    .C(_0716_),
    .X(_0724_));
 sky130_fd_sc_hd__nor2_1 _1373_ (.A(net78),
    .B(_0304_),
    .Y(_0725_));
 sky130_fd_sc_hd__or4b_1 _1374_ (.A(_0274_),
    .B(_0302_),
    .C(net53),
    .D_N(_0340_),
    .X(_0726_));
 sky130_fd_sc_hd__or4_4 _1375_ (.A(_0723_),
    .B(_0724_),
    .C(_0725_),
    .D(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__a211o_4 _1376_ (.A1(net84),
    .A2(_0279_),
    .B1(_0547_),
    .C1(_0269_),
    .X(_0728_));
 sky130_fd_sc_hd__or3_4 _1377_ (.A(net65),
    .B(_0287_),
    .C(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__o21bai_4 _1378_ (.A1(net77),
    .A2(_0252_),
    .B1_N(_0275_),
    .Y(_0730_));
 sky130_fd_sc_hd__a22o_1 _1379_ (.A1(\MOS6502.ADD[0] ),
    .A2(_0727_),
    .B1(net49),
    .B2(net1),
    .X(_0731_));
 sky130_fd_sc_hd__nor4_4 _1380_ (.A(_0721_),
    .B(_0727_),
    .C(_0729_),
    .D(net49),
    .Y(_0732_));
 sky130_fd_sc_hd__or4_4 _1381_ (.A(_0721_),
    .B(_0727_),
    .C(_0729_),
    .D(net49),
    .X(_0733_));
 sky130_fd_sc_hd__a2bb2o_1 _1382_ (.A1_N(_0456_),
    .A2_N(_0720_),
    .B1(net40),
    .B2(\MOS6502.PC[0] ),
    .X(_0734_));
 sky130_fd_sc_hd__a211o_1 _1383_ (.A1(\MOS6502.ABL[0] ),
    .A2(_0729_),
    .B1(_0731_),
    .C1(_0734_),
    .X(net14));
 sky130_fd_sc_hd__a221o_1 _1384_ (.A1(\MOS6502.ABL[1] ),
    .A2(_0729_),
    .B1(net49),
    .B2(net2),
    .C1(net40),
    .X(_0735_));
 sky130_fd_sc_hd__a22o_1 _1385_ (.A1(_0439_),
    .A2(_0721_),
    .B1(_0727_),
    .B2(\MOS6502.ADD[1] ),
    .X(_0736_));
 sky130_fd_sc_hd__o22a_1 _1386_ (.A1(\MOS6502.PC[1] ),
    .A2(_0733_),
    .B1(_0735_),
    .B2(_0736_),
    .X(net15));
 sky130_fd_sc_hd__a221o_1 _1387_ (.A1(\MOS6502.ABL[2] ),
    .A2(_0729_),
    .B1(net49),
    .B2(net3),
    .C1(net40),
    .X(_0737_));
 sky130_fd_sc_hd__a2bb2o_1 _1388_ (.A1_N(_0423_),
    .A2_N(_0720_),
    .B1(_0727_),
    .B2(\MOS6502.ADD[2] ),
    .X(_0738_));
 sky130_fd_sc_hd__o22a_1 _1389_ (.A1(\MOS6502.PC[2] ),
    .A2(_0733_),
    .B1(_0737_),
    .B2(_0738_),
    .X(net16));
 sky130_fd_sc_hd__a221o_1 _1390_ (.A1(\MOS6502.ABL[3] ),
    .A2(_0729_),
    .B1(net49),
    .B2(net4),
    .C1(net40),
    .X(_0739_));
 sky130_fd_sc_hd__a2bb2o_1 _1391_ (.A1_N(_0404_),
    .A2_N(_0720_),
    .B1(_0727_),
    .B2(\MOS6502.ADD[3] ),
    .X(_0740_));
 sky130_fd_sc_hd__o22a_1 _1392_ (.A1(\MOS6502.PC[3] ),
    .A2(_0733_),
    .B1(_0739_),
    .B2(_0740_),
    .X(net17));
 sky130_fd_sc_hd__a221o_1 _1393_ (.A1(\MOS6502.ABL[4] ),
    .A2(_0729_),
    .B1(net49),
    .B2(net5),
    .C1(net40),
    .X(_0741_));
 sky130_fd_sc_hd__a2bb2o_1 _1394_ (.A1_N(_0386_),
    .A2_N(_0720_),
    .B1(_0727_),
    .B2(\MOS6502.ADD[4] ),
    .X(_0742_));
 sky130_fd_sc_hd__o22a_1 _1395_ (.A1(\MOS6502.PC[4] ),
    .A2(_0733_),
    .B1(_0741_),
    .B2(_0742_),
    .X(net18));
 sky130_fd_sc_hd__a221o_1 _1396_ (.A1(\MOS6502.ABL[5] ),
    .A2(_0729_),
    .B1(net49),
    .B2(net6),
    .C1(net40),
    .X(_0743_));
 sky130_fd_sc_hd__a2bb2o_1 _1397_ (.A1_N(_0350_),
    .A2_N(_0720_),
    .B1(_0727_),
    .B2(\MOS6502.ADD[5] ),
    .X(_0744_));
 sky130_fd_sc_hd__o22a_1 _1398_ (.A1(\MOS6502.PC[5] ),
    .A2(_0733_),
    .B1(_0743_),
    .B2(_0744_),
    .X(net19));
 sky130_fd_sc_hd__a221o_1 _1399_ (.A1(\MOS6502.ABL[6] ),
    .A2(_0729_),
    .B1(net49),
    .B2(net7),
    .C1(net40),
    .X(_0745_));
 sky130_fd_sc_hd__a2bb2o_1 _1400_ (.A1_N(_0334_),
    .A2_N(_0720_),
    .B1(_0727_),
    .B2(\MOS6502.ADD[6] ),
    .X(_0746_));
 sky130_fd_sc_hd__o22a_1 _1401_ (.A1(\MOS6502.PC[6] ),
    .A2(_0733_),
    .B1(_0745_),
    .B2(_0746_),
    .X(net20));
 sky130_fd_sc_hd__a221o_1 _1402_ (.A1(\MOS6502.ABL[7] ),
    .A2(_0729_),
    .B1(_0730_),
    .B2(net8),
    .C1(net40),
    .X(_0747_));
 sky130_fd_sc_hd__a2bb2o_1 _1403_ (.A1_N(_0497_),
    .A2_N(_0720_),
    .B1(_0727_),
    .B2(\MOS6502.ADD[7] ),
    .X(_0748_));
 sky130_fd_sc_hd__o22a_1 _1404_ (.A1(\MOS6502.PC[7] ),
    .A2(_0733_),
    .B1(_0747_),
    .B2(_0748_),
    .X(net21));
 sky130_fd_sc_hd__a211o_1 _1405_ (.A1(\MOS6502.ADD[0] ),
    .A2(_0728_),
    .B1(_0724_),
    .C1(_0721_),
    .X(_0749_));
 sky130_fd_sc_hd__or3_4 _1406_ (.A(net65),
    .B(_0287_),
    .C(net53),
    .X(_0750_));
 sky130_fd_sc_hd__a22o_1 _1407_ (.A1(net1),
    .A2(_0723_),
    .B1(_0750_),
    .B2(\MOS6502.ABH[0] ),
    .X(_0751_));
 sky130_fd_sc_hd__a211o_1 _1408_ (.A1(\MOS6502.PC[8] ),
    .A2(net40),
    .B1(_0749_),
    .C1(_0751_),
    .X(net22));
 sky130_fd_sc_hd__a22o_1 _1409_ (.A1(net2),
    .A2(_0723_),
    .B1(_0750_),
    .B2(\MOS6502.ABH[1] ),
    .X(_0752_));
 sky130_fd_sc_hd__a211o_1 _1410_ (.A1(\MOS6502.ADD[1] ),
    .A2(_0728_),
    .B1(net40),
    .C1(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__o21a_1 _1411_ (.A1(\MOS6502.PC[9] ),
    .A2(_0733_),
    .B1(_0753_),
    .X(net23));
 sky130_fd_sc_hd__a22o_1 _1412_ (.A1(net3),
    .A2(_0723_),
    .B1(_0728_),
    .B2(\MOS6502.ADD[2] ),
    .X(_0754_));
 sky130_fd_sc_hd__a221o_1 _1413_ (.A1(\MOS6502.PC[10] ),
    .A2(net41),
    .B1(_0750_),
    .B2(\MOS6502.ABH[2] ),
    .C1(_0754_),
    .X(net25));
 sky130_fd_sc_hd__a22o_1 _1414_ (.A1(net4),
    .A2(_0723_),
    .B1(_0728_),
    .B2(\MOS6502.ADD[3] ),
    .X(_0755_));
 sky130_fd_sc_hd__a221o_1 _1415_ (.A1(\MOS6502.PC[11] ),
    .A2(net41),
    .B1(_0750_),
    .B2(\MOS6502.ABH[3] ),
    .C1(_0755_),
    .X(net26));
 sky130_fd_sc_hd__a22o_1 _1416_ (.A1(net5),
    .A2(_0723_),
    .B1(_0728_),
    .B2(\MOS6502.ADD[4] ),
    .X(_0756_));
 sky130_fd_sc_hd__a221o_1 _1417_ (.A1(\MOS6502.PC[12] ),
    .A2(net41),
    .B1(_0750_),
    .B2(\MOS6502.ABH[4] ),
    .C1(_0756_),
    .X(net27));
 sky130_fd_sc_hd__a22o_1 _1418_ (.A1(net6),
    .A2(_0723_),
    .B1(_0728_),
    .B2(\MOS6502.ADD[5] ),
    .X(_0757_));
 sky130_fd_sc_hd__a221o_1 _1419_ (.A1(\MOS6502.PC[13] ),
    .A2(net41),
    .B1(_0750_),
    .B2(\MOS6502.ABH[5] ),
    .C1(_0757_),
    .X(net28));
 sky130_fd_sc_hd__a22o_1 _1420_ (.A1(net7),
    .A2(_0723_),
    .B1(_0728_),
    .B2(\MOS6502.ADD[6] ),
    .X(_0758_));
 sky130_fd_sc_hd__a221o_1 _1421_ (.A1(\MOS6502.PC[14] ),
    .A2(net41),
    .B1(_0750_),
    .B2(\MOS6502.ABH[6] ),
    .C1(_0758_),
    .X(net29));
 sky130_fd_sc_hd__a22o_1 _1422_ (.A1(net8),
    .A2(_0723_),
    .B1(_0728_),
    .B2(\MOS6502.ADD[7] ),
    .X(_0759_));
 sky130_fd_sc_hd__a221o_1 _1423_ (.A1(\MOS6502.PC[15] ),
    .A2(net41),
    .B1(_0750_),
    .B2(\MOS6502.ABH[7] ),
    .C1(_0759_),
    .X(net30));
 sky130_fd_sc_hd__a21o_2 _1424_ (.A1(\MOS6502.php ),
    .A2(_0253_),
    .B1(net69),
    .X(_0760_));
 sky130_fd_sc_hd__o21bai_4 _1425_ (.A1(\MOS6502.php ),
    .A2(_0254_),
    .B1_N(net65),
    .Y(_0761_));
 sky130_fd_sc_hd__a22o_1 _1426_ (.A1(\MOS6502.PC[8] ),
    .A2(net51),
    .B1(_0760_),
    .B2(\MOS6502.C ),
    .X(_0762_));
 sky130_fd_sc_hd__a22o_1 _1427_ (.A1(\MOS6502.PC[0] ),
    .A2(net48),
    .B1(_0761_),
    .B2(\MOS6502.ADD[0] ),
    .X(_0763_));
 sky130_fd_sc_hd__nand2_1 _1428_ (.A(_0266_),
    .B(_0456_),
    .Y(_0764_));
 sky130_fd_sc_hd__o31a_2 _1429_ (.A1(_0266_),
    .A2(_0762_),
    .A3(_0763_),
    .B1(_0764_),
    .X(net13));
 sky130_fd_sc_hd__a22o_1 _1430_ (.A1(\MOS6502.PC[1] ),
    .A2(net48),
    .B1(_0760_),
    .B2(\MOS6502.Z ),
    .X(_0765_));
 sky130_fd_sc_hd__a221o_1 _1431_ (.A1(\MOS6502.PC[9] ),
    .A2(net51),
    .B1(_0761_),
    .B2(\MOS6502.ADD[1] ),
    .C1(_0266_),
    .X(_0766_));
 sky130_fd_sc_hd__o22a_2 _1432_ (.A1(_0267_),
    .A2(_0439_),
    .B1(_0765_),
    .B2(_0766_),
    .X(net24));
 sky130_fd_sc_hd__a22o_1 _1433_ (.A1(\MOS6502.PC[2] ),
    .A2(net48),
    .B1(_0760_),
    .B2(\MOS6502.I ),
    .X(_0767_));
 sky130_fd_sc_hd__a22o_1 _1434_ (.A1(\MOS6502.PC[10] ),
    .A2(_0259_),
    .B1(_0761_),
    .B2(\MOS6502.ADD[2] ),
    .X(_0768_));
 sky130_fd_sc_hd__nand2_1 _1435_ (.A(_0266_),
    .B(_0423_),
    .Y(_0769_));
 sky130_fd_sc_hd__o31a_2 _1436_ (.A1(_0266_),
    .A2(_0767_),
    .A3(_0768_),
    .B1(_0769_),
    .X(net32));
 sky130_fd_sc_hd__a22o_1 _1437_ (.A1(\MOS6502.PC[3] ),
    .A2(net48),
    .B1(net51),
    .B2(\MOS6502.PC[11] ),
    .X(_0770_));
 sky130_fd_sc_hd__a221o_1 _1438_ (.A1(\MOS6502.D ),
    .A2(_0760_),
    .B1(_0761_),
    .B2(\MOS6502.ADD[3] ),
    .C1(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__o21bai_4 _1439_ (.A1(_0267_),
    .A2(_0404_),
    .B1_N(_0771_),
    .Y(net33));
 sky130_fd_sc_hd__o21a_1 _1440_ (.A1(_0253_),
    .A2(net65),
    .B1(\MOS6502.ADD[4] ),
    .X(_0772_));
 sky130_fd_sc_hd__a221o_1 _1441_ (.A1(\MOS6502.PC[4] ),
    .A2(net48),
    .B1(net51),
    .B2(\MOS6502.PC[12] ),
    .C1(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__a21oi_1 _1442_ (.A1(\MOS6502.php ),
    .A2(_0253_),
    .B1(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__o31a_2 _1443_ (.A1(\MOS6502.NMI_edge ),
    .A2(net9),
    .A3(_0249_),
    .B1(_0774_),
    .X(_0775_));
 sky130_fd_sc_hd__o21ai_2 _1444_ (.A1(_0267_),
    .A2(_0386_),
    .B1(_0775_),
    .Y(net34));
 sky130_fd_sc_hd__nor2_1 _1445_ (.A(_0267_),
    .B(_0350_),
    .Y(_0776_));
 sky130_fd_sc_hd__o21a_1 _1446_ (.A1(_0253_),
    .A2(_0265_),
    .B1(\MOS6502.ADD[5] ),
    .X(_0777_));
 sky130_fd_sc_hd__a221o_1 _1447_ (.A1(\MOS6502.PC[5] ),
    .A2(net48),
    .B1(net51),
    .B2(\MOS6502.PC[13] ),
    .C1(_0760_),
    .X(_0778_));
 sky130_fd_sc_hd__or3_2 _1448_ (.A(_0776_),
    .B(_0777_),
    .C(_0778_),
    .X(net35));
 sky130_fd_sc_hd__a22o_1 _1449_ (.A1(\MOS6502.PC[6] ),
    .A2(net48),
    .B1(_0760_),
    .B2(\MOS6502.V ),
    .X(_0779_));
 sky130_fd_sc_hd__a221o_1 _1450_ (.A1(\MOS6502.PC[14] ),
    .A2(net51),
    .B1(_0761_),
    .B2(\MOS6502.ADD[6] ),
    .C1(_0266_),
    .X(_0780_));
 sky130_fd_sc_hd__o2bb2a_1 _1451_ (.A1_N(_0266_),
    .A2_N(_0334_),
    .B1(_0779_),
    .B2(_0780_),
    .X(net36));
 sky130_fd_sc_hd__a22o_1 _1452_ (.A1(\MOS6502.PC[7] ),
    .A2(net48),
    .B1(net51),
    .B2(\MOS6502.PC[15] ),
    .X(_0781_));
 sky130_fd_sc_hd__a2bb2o_1 _1453_ (.A1_N(_0267_),
    .A2_N(_0497_),
    .B1(_0761_),
    .B2(\MOS6502.ADD[7] ),
    .X(_0782_));
 sky130_fd_sc_hd__a211o_2 _1454_ (.A1(\MOS6502.N ),
    .A2(_0760_),
    .B1(_0781_),
    .C1(_0782_),
    .X(net37));
 sky130_fd_sc_hd__or3b_4 _1455_ (.A(net60),
    .B(net79),
    .C_N(\MOS6502.load_reg ),
    .X(_0783_));
 sky130_fd_sc_hd__nand3_4 _1456_ (.A(_0710_),
    .B(_0715_),
    .C(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__and3_4 _1457_ (.A(net45),
    .B(net44),
    .C(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__mux2_2 _1458_ (.A0(\MOS6502.ADD[0] ),
    .A1(net1),
    .S(net66),
    .X(_0786_));
 sky130_fd_sc_hd__mux2_1 _1459_ (.A0(\MOS6502.AXYS[2][0] ),
    .A1(_0786_),
    .S(_0785_),
    .X(_0030_));
 sky130_fd_sc_hd__and3_1 _1460_ (.A(\MOS6502.adc_bcd ),
    .B(\MOS6502.adj_bcd ),
    .C(\MOS6502.ALU.HC ),
    .X(_0787_));
 sky130_fd_sc_hd__nand2b_2 _1461_ (.A_N(\MOS6502.adc_bcd ),
    .B(\MOS6502.adj_bcd ),
    .Y(_0788_));
 sky130_fd_sc_hd__nor2_2 _1462_ (.A(\MOS6502.ALU.HC ),
    .B(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__or3_1 _1463_ (.A(\MOS6502.ADD[1] ),
    .B(_0787_),
    .C(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__o21a_1 _1464_ (.A1(_0787_),
    .A2(_0789_),
    .B1(\MOS6502.ADD[1] ),
    .X(_0791_));
 sky130_fd_sc_hd__nor2_1 _1465_ (.A(net66),
    .B(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__a22o_2 _1466_ (.A1(net2),
    .A2(net66),
    .B1(_0790_),
    .B2(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__mux2_1 _1467_ (.A0(\MOS6502.AXYS[2][1] ),
    .A1(_0793_),
    .S(_0785_),
    .X(_0031_));
 sky130_fd_sc_hd__or2_1 _1468_ (.A(\MOS6502.ADD[2] ),
    .B(_0787_),
    .X(_0794_));
 sky130_fd_sc_hd__nand2_1 _1469_ (.A(\MOS6502.ADD[2] ),
    .B(_0787_),
    .Y(_0795_));
 sky130_fd_sc_hd__a21oi_1 _1470_ (.A1(_0794_),
    .A2(_0795_),
    .B1(_0791_),
    .Y(_0796_));
 sky130_fd_sc_hd__a31o_1 _1471_ (.A1(_0791_),
    .A2(_0794_),
    .A3(_0795_),
    .B1(net66),
    .X(_0797_));
 sky130_fd_sc_hd__a2bb2o_2 _1472_ (.A1_N(_0796_),
    .A2_N(_0797_),
    .B1(net3),
    .B2(net66),
    .X(_0798_));
 sky130_fd_sc_hd__mux2_1 _1473_ (.A0(\MOS6502.AXYS[2][2] ),
    .A1(_0798_),
    .S(_0785_),
    .X(_0032_));
 sky130_fd_sc_hd__a21bo_1 _1474_ (.A1(_0791_),
    .A2(_0794_),
    .B1_N(_0795_),
    .X(_0799_));
 sky130_fd_sc_hd__xnor2_1 _1475_ (.A(\MOS6502.ADD[3] ),
    .B(_0789_),
    .Y(_0800_));
 sky130_fd_sc_hd__xnor2_1 _1476_ (.A(_0799_),
    .B(_0800_),
    .Y(_0801_));
 sky130_fd_sc_hd__mux2_4 _1477_ (.A0(_0801_),
    .A1(net4),
    .S(net66),
    .X(_0802_));
 sky130_fd_sc_hd__mux2_1 _1478_ (.A0(\MOS6502.AXYS[2][3] ),
    .A1(_0802_),
    .S(_0785_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_2 _1479_ (.A0(\MOS6502.ADD[4] ),
    .A1(net5),
    .S(net66),
    .X(_0803_));
 sky130_fd_sc_hd__mux2_1 _1480_ (.A0(\MOS6502.AXYS[2][4] ),
    .A1(_0803_),
    .S(_0785_),
    .X(_0034_));
 sky130_fd_sc_hd__and3_1 _1481_ (.A(\MOS6502.ALU.CO ),
    .B(\MOS6502.adc_bcd ),
    .C(\MOS6502.adj_bcd ),
    .X(_0804_));
 sky130_fd_sc_hd__nor2_2 _1482_ (.A(\MOS6502.ALU.CO ),
    .B(_0788_),
    .Y(_0805_));
 sky130_fd_sc_hd__o21a_1 _1483_ (.A1(_0804_),
    .A2(_0805_),
    .B1(\MOS6502.ADD[5] ),
    .X(_0806_));
 sky130_fd_sc_hd__or3_1 _1484_ (.A(\MOS6502.ADD[5] ),
    .B(_0804_),
    .C(_0805_),
    .X(_0807_));
 sky130_fd_sc_hd__or3b_1 _1485_ (.A(net67),
    .B(_0806_),
    .C_N(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__a21bo_2 _1486_ (.A1(net6),
    .A2(net66),
    .B1_N(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__mux2_1 _1487_ (.A0(\MOS6502.AXYS[2][5] ),
    .A1(_0809_),
    .S(_0785_),
    .X(_0035_));
 sky130_fd_sc_hd__or2_1 _1488_ (.A(\MOS6502.ADD[6] ),
    .B(_0804_),
    .X(_0810_));
 sky130_fd_sc_hd__nand2_1 _1489_ (.A(\MOS6502.ADD[6] ),
    .B(_0804_),
    .Y(_0811_));
 sky130_fd_sc_hd__a21oi_1 _1490_ (.A1(_0810_),
    .A2(_0811_),
    .B1(_0806_),
    .Y(_0812_));
 sky130_fd_sc_hd__a31o_1 _1491_ (.A1(_0806_),
    .A2(_0810_),
    .A3(_0811_),
    .B1(net66),
    .X(_0813_));
 sky130_fd_sc_hd__a2bb2o_4 _1492_ (.A1_N(_0812_),
    .A2_N(_0813_),
    .B1(net7),
    .B2(net66),
    .X(_0814_));
 sky130_fd_sc_hd__mux2_1 _1493_ (.A0(\MOS6502.AXYS[2][6] ),
    .A1(_0814_),
    .S(_0785_),
    .X(_0036_));
 sky130_fd_sc_hd__a21bo_1 _1494_ (.A1(_0806_),
    .A2(_0810_),
    .B1_N(_0811_),
    .X(_0815_));
 sky130_fd_sc_hd__xnor2_1 _1495_ (.A(\MOS6502.ADD[7] ),
    .B(_0805_),
    .Y(_0816_));
 sky130_fd_sc_hd__nor2_1 _1496_ (.A(_0815_),
    .B(_0816_),
    .Y(_0817_));
 sky130_fd_sc_hd__a21o_1 _1497_ (.A1(_0815_),
    .A2(_0816_),
    .B1(net67),
    .X(_0818_));
 sky130_fd_sc_hd__o32a_4 _1498_ (.A1(net8),
    .A2(net78),
    .A3(_0247_),
    .B1(_0817_),
    .B2(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__mux2_1 _1499_ (.A0(\MOS6502.AXYS[2][7] ),
    .A1(_0819_),
    .S(_0785_),
    .X(_0037_));
 sky130_fd_sc_hd__and2_4 _1500_ (.A(_0333_),
    .B(_0784_),
    .X(_0820_));
 sky130_fd_sc_hd__mux2_1 _1501_ (.A0(\MOS6502.AXYS[1][0] ),
    .A1(_0786_),
    .S(_0820_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _1502_ (.A0(\MOS6502.AXYS[1][1] ),
    .A1(_0793_),
    .S(_0820_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _1503_ (.A0(\MOS6502.AXYS[1][2] ),
    .A1(_0798_),
    .S(_0820_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _1504_ (.A0(\MOS6502.AXYS[1][3] ),
    .A1(_0802_),
    .S(_0820_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _1505_ (.A0(\MOS6502.AXYS[1][4] ),
    .A1(_0803_),
    .S(_0820_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _1506_ (.A0(\MOS6502.AXYS[1][5] ),
    .A1(_0809_),
    .S(_0820_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _1507_ (.A0(\MOS6502.AXYS[1][6] ),
    .A1(_0814_),
    .S(_0820_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _1508_ (.A0(\MOS6502.AXYS[1][7] ),
    .A1(_0819_),
    .S(_0820_),
    .X(_0045_));
 sky130_fd_sc_hd__a21oi_1 _1509_ (.A1(_0292_),
    .A2(_0304_),
    .B1(\MOS6502.state[5] ),
    .Y(_0821_));
 sky130_fd_sc_hd__or2_2 _1510_ (.A(net65),
    .B(net64),
    .X(_0822_));
 sky130_fd_sc_hd__nand2_1 _1511_ (.A(_0270_),
    .B(_0528_),
    .Y(_0823_));
 sky130_fd_sc_hd__or4_1 _1512_ (.A(_0258_),
    .B(_0293_),
    .C(_0307_),
    .D(_0640_),
    .X(_0824_));
 sky130_fd_sc_hd__or4_1 _1513_ (.A(_0248_),
    .B(_0269_),
    .C(_0288_),
    .D(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__or3_1 _1514_ (.A(_0705_),
    .B(net49),
    .C(_0822_),
    .X(_0826_));
 sky130_fd_sc_hd__or3_1 _1515_ (.A(_0301_),
    .B(_0321_),
    .C(_0472_),
    .X(_0827_));
 sky130_fd_sc_hd__or4_1 _1516_ (.A(_0359_),
    .B(_0825_),
    .C(_0826_),
    .D(_0827_),
    .X(_0125_));
 sky130_fd_sc_hd__or4b_1 _1517_ (.A(_0821_),
    .B(_0823_),
    .C(_0125_),
    .D_N(_0539_),
    .X(_0126_));
 sky130_fd_sc_hd__and3_2 _1518_ (.A(_0254_),
    .B(_0300_),
    .C(_0126_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _1519_ (.A0(\MOS6502.ABL[0] ),
    .A1(net14),
    .S(net38),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _1520_ (.A0(\MOS6502.ABL[1] ),
    .A1(net15),
    .S(net38),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _1521_ (.A0(\MOS6502.ABL[2] ),
    .A1(net16),
    .S(net38),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _1522_ (.A0(\MOS6502.ABL[3] ),
    .A1(net17),
    .S(net38),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _1523_ (.A0(\MOS6502.ABL[4] ),
    .A1(net18),
    .S(net38),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _1524_ (.A0(\MOS6502.ABL[5] ),
    .A1(net19),
    .S(net38),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _1525_ (.A0(\MOS6502.ABL[6] ),
    .A1(net20),
    .S(net38),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _1526_ (.A0(\MOS6502.ABL[7] ),
    .A1(net21),
    .S(net38),
    .X(_0053_));
 sky130_fd_sc_hd__or3_1 _1527_ (.A(\MOS6502.adc_sbc ),
    .B(\MOS6502.compare ),
    .C(\MOS6502.shift ),
    .X(_0128_));
 sky130_fd_sc_hd__or4_1 _1528_ (.A(net79),
    .B(\MOS6502.state[1] ),
    .C(\MOS6502.clc ),
    .D(\MOS6502.sec ),
    .X(_0129_));
 sky130_fd_sc_hd__a2bb2o_1 _1529_ (.A1_N(\MOS6502.write_back ),
    .A2_N(net57),
    .B1(net65),
    .B2(\MOS6502.shift ),
    .X(_0130_));
 sky130_fd_sc_hd__o22a_1 _1530_ (.A1(_0128_),
    .A2(_0129_),
    .B1(_0130_),
    .B2(_0354_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _1531_ (.A0(_0229_),
    .A1(\MOS6502.ADD[0] ),
    .S(net79),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _1532_ (.A0(_0132_),
    .A1(\MOS6502.ALU.CO ),
    .S(_0128_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _1533_ (.A0(net1),
    .A1(_0133_),
    .S(_0355_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _1534_ (.A0(\MOS6502.C ),
    .A1(_0134_),
    .S(_0131_),
    .X(_0054_));
 sky130_fd_sc_hd__o21a_1 _1535_ (.A1(net45),
    .A2(net44),
    .B1(\MOS6502.load_reg ),
    .X(_0135_));
 sky130_fd_sc_hd__or4_1 _1536_ (.A(net79),
    .B(\MOS6502.compare ),
    .C(net57),
    .D(_0135_),
    .X(_0136_));
 sky130_fd_sc_hd__o22a_1 _1537_ (.A1(_0354_),
    .A2(_0822_),
    .B1(_0136_),
    .B2(\MOS6502.bit_ins ),
    .X(_0137_));
 sky130_fd_sc_hd__o21ba_1 _1538_ (.A1(net79),
    .A2(_0354_),
    .B1_N(net65),
    .X(_0138_));
 sky130_fd_sc_hd__or4_1 _1539_ (.A(\MOS6502.ADD[4] ),
    .B(\MOS6502.ADD[5] ),
    .C(\MOS6502.ADD[6] ),
    .D(\MOS6502.ADD[7] ),
    .X(_0139_));
 sky130_fd_sc_hd__or4_1 _1540_ (.A(\MOS6502.ADD[0] ),
    .B(\MOS6502.ADD[1] ),
    .C(\MOS6502.ADD[2] ),
    .D(\MOS6502.ADD[3] ),
    .X(_0140_));
 sky130_fd_sc_hd__nor2_1 _1541_ (.A(_0139_),
    .B(_0140_),
    .Y(_0141_));
 sky130_fd_sc_hd__mux2_1 _1542_ (.A0(\MOS6502.ADD[1] ),
    .A1(net2),
    .S(_0354_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _1543_ (.A0(_0141_),
    .A1(_0142_),
    .S(_0138_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _1544_ (.A0(\MOS6502.Z ),
    .A1(_0143_),
    .S(_0137_),
    .X(_0055_));
 sky130_fd_sc_hd__a211o_1 _1545_ (.A1(\MOS6502.bit_ins ),
    .A2(_0282_),
    .B1(net63),
    .C1(_0354_),
    .X(_0144_));
 sky130_fd_sc_hd__o21a_1 _1546_ (.A1(net65),
    .A2(_0144_),
    .B1(_0136_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _1547_ (.A0(net8),
    .A1(\MOS6502.ADD[7] ),
    .S(_0822_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _1548_ (.A0(\MOS6502.N ),
    .A1(_0146_),
    .S(_0145_),
    .X(_0056_));
 sky130_fd_sc_hd__or4_1 _1549_ (.A(net79),
    .B(\MOS6502.cld ),
    .C(\MOS6502.sed ),
    .D(net57),
    .X(_0147_));
 sky130_fd_sc_hd__o21a_1 _1550_ (.A1(net63),
    .A2(_0354_),
    .B1(_0147_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _1551_ (.A0(_0224_),
    .A1(\MOS6502.ADD[3] ),
    .S(net79),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _1552_ (.A0(net4),
    .A1(_0149_),
    .S(_0355_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _1553_ (.A0(\MOS6502.D ),
    .A1(_0150_),
    .S(_0148_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _1554_ (.A0(\MOS6502.ADD[2] ),
    .A1(_0225_),
    .S(_0286_),
    .X(_0151_));
 sky130_fd_sc_hd__o32a_1 _1555_ (.A1(\MOS6502.cli ),
    .A2(\MOS6502.sei ),
    .A3(_0268_),
    .B1(_0223_),
    .B2(\MOS6502.plp ),
    .X(_0152_));
 sky130_fd_sc_hd__o31a_1 _1556_ (.A1(_0286_),
    .A2(net64),
    .A3(_0354_),
    .B1(_0152_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _1557_ (.A0(net3),
    .A1(_0151_),
    .S(_0355_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _1558_ (.A0(\MOS6502.I ),
    .A1(_0154_),
    .S(_0153_),
    .X(_0155_));
 sky130_fd_sc_hd__or2_1 _1559_ (.A(_0318_),
    .B(_0155_),
    .X(_0058_));
 sky130_fd_sc_hd__nor2_1 _1560_ (.A(net79),
    .B(\MOS6502.clv ),
    .Y(_0156_));
 sky130_fd_sc_hd__o41a_1 _1561_ (.A1(net79),
    .A2(\MOS6502.adc_sbc ),
    .A3(\MOS6502.clv ),
    .A4(net57),
    .B1(_0144_),
    .X(_0157_));
 sky130_fd_sc_hd__xor2_1 _1562_ (.A(\MOS6502.ALU.BI7 ),
    .B(\MOS6502.ALU.AI7 ),
    .X(_0158_));
 sky130_fd_sc_hd__xnor2_1 _1563_ (.A(\MOS6502.ADD[7] ),
    .B(\MOS6502.ALU.CO ),
    .Y(_0159_));
 sky130_fd_sc_hd__xnor2_1 _1564_ (.A(_0158_),
    .B(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__a221o_1 _1565_ (.A1(net79),
    .A2(\MOS6502.ADD[6] ),
    .B1(_0156_),
    .B2(_0160_),
    .C1(net57),
    .X(_0161_));
 sky130_fd_sc_hd__o21a_1 _1566_ (.A1(net7),
    .A2(net63),
    .B1(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _1567_ (.A0(\MOS6502.V ),
    .A1(_0162_),
    .S(_0157_),
    .X(_0059_));
 sky130_fd_sc_hd__or2_4 _1568_ (.A(net11),
    .B(_0300_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _1569_ (.A0(net1),
    .A1(\MOS6502.IRHOLD[0] ),
    .S(_0163_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _1570_ (.A0(net2),
    .A1(\MOS6502.IRHOLD[1] ),
    .S(_0163_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _1571_ (.A0(net3),
    .A1(\MOS6502.IRHOLD[2] ),
    .S(_0163_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _1572_ (.A0(net4),
    .A1(\MOS6502.IRHOLD[3] ),
    .S(_0163_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _1573_ (.A0(net5),
    .A1(\MOS6502.IRHOLD[4] ),
    .S(_0163_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _1574_ (.A0(net6),
    .A1(\MOS6502.IRHOLD[5] ),
    .S(_0163_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _1575_ (.A0(net7),
    .A1(\MOS6502.IRHOLD[6] ),
    .S(_0163_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _1576_ (.A0(net8),
    .A1(\MOS6502.IRHOLD[7] ),
    .S(_0163_),
    .X(_0067_));
 sky130_fd_sc_hd__nand2_1 _1577_ (.A(\MOS6502.IRHOLD_valid ),
    .B(net60),
    .Y(_0164_));
 sky130_fd_sc_hd__a21oi_1 _1578_ (.A1(_0300_),
    .A2(_0164_),
    .B1(net11),
    .Y(_0068_));
 sky130_fd_sc_hd__and3_2 _1579_ (.A(net71),
    .B(_0231_),
    .C(_0235_),
    .X(_0165_));
 sky130_fd_sc_hd__nor2_2 _1580_ (.A(_0627_),
    .B(_0682_),
    .Y(_0166_));
 sky130_fd_sc_hd__nand2_4 _1581_ (.A(\MOS6502.IR[7] ),
    .B(_0236_),
    .Y(_0167_));
 sky130_fd_sc_hd__nor2_1 _1582_ (.A(_0232_),
    .B(\MOS6502.IR[5] ),
    .Y(_0168_));
 sky130_fd_sc_hd__nor2_2 _1583_ (.A(_0233_),
    .B(_0167_),
    .Y(_0169_));
 sky130_fd_sc_hd__a22o_1 _1584_ (.A1(_0165_),
    .A2(_0166_),
    .B1(_0169_),
    .B2(_0634_),
    .X(_0170_));
 sky130_fd_sc_hd__nor2_1 _1585_ (.A(net52),
    .B(_0167_),
    .Y(_0171_));
 sky130_fd_sc_hd__or4_1 _1586_ (.A(_0234_),
    .B(_0601_),
    .C(_0608_),
    .D(_0167_),
    .X(_0172_));
 sky130_fd_sc_hd__and3_1 _1587_ (.A(\MOS6502.IR[7] ),
    .B(_0236_),
    .C(net72),
    .X(_0173_));
 sky130_fd_sc_hd__nand2_2 _1588_ (.A(\MOS6502.IR[5] ),
    .B(_0173_),
    .Y(_0174_));
 sky130_fd_sc_hd__nor2_1 _1589_ (.A(_0682_),
    .B(_0167_),
    .Y(_0175_));
 sky130_fd_sc_hd__a21oi_1 _1590_ (.A1(_0632_),
    .A2(_0174_),
    .B1(_0682_),
    .Y(_0176_));
 sky130_fd_sc_hd__and2_2 _1591_ (.A(net50),
    .B(_0635_),
    .X(_0177_));
 sky130_fd_sc_hd__o221a_1 _1592_ (.A1(_0612_),
    .A2(_0168_),
    .B1(_0174_),
    .B2(_0656_),
    .C1(_0172_),
    .X(_0178_));
 sky130_fd_sc_hd__or4b_1 _1593_ (.A(_0170_),
    .B(_0176_),
    .C(_0177_),
    .D_N(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _1594_ (.A0(\MOS6502.load_reg ),
    .A1(_0179_),
    .S(net61),
    .X(_0069_));
 sky130_fd_sc_hd__a21o_1 _1595_ (.A1(\MOS6502.res ),
    .A2(net60),
    .B1(net11),
    .X(_0070_));
 sky130_fd_sc_hd__nor2_1 _1596_ (.A(net47),
    .B(_0650_),
    .Y(_0180_));
 sky130_fd_sc_hd__a2111o_1 _1597_ (.A1(net72),
    .A2(_0614_),
    .B1(net47),
    .C1(_0167_),
    .D1(net52),
    .X(_0181_));
 sky130_fd_sc_hd__a21bo_1 _1598_ (.A1(_0168_),
    .A2(_0177_),
    .B1_N(_0181_),
    .X(_0182_));
 sky130_fd_sc_hd__a31o_1 _1599_ (.A1(net52),
    .A2(_0601_),
    .A3(_0175_),
    .B1(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__a21o_1 _1600_ (.A1(\MOS6502.dst_reg[0] ),
    .A2(net57),
    .B1(_0637_),
    .X(_0184_));
 sky130_fd_sc_hd__a21o_1 _1601_ (.A1(net62),
    .A2(_0183_),
    .B1(_0184_),
    .X(_0071_));
 sky130_fd_sc_hd__and2_2 _1602_ (.A(net61),
    .B(_0165_),
    .X(_0185_));
 sky130_fd_sc_hd__o21a_1 _1603_ (.A1(_0166_),
    .A2(_0177_),
    .B1(_0165_),
    .X(_0186_));
 sky130_fd_sc_hd__a211o_1 _1604_ (.A1(_0678_),
    .A2(_0171_),
    .B1(_0182_),
    .C1(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _1605_ (.A0(\MOS6502.dst_reg[1] ),
    .A1(_0187_),
    .S(net62),
    .X(_0072_));
 sky130_fd_sc_hd__or2_1 _1606_ (.A(\MOS6502.IR[6] ),
    .B(_0616_),
    .X(_0188_));
 sky130_fd_sc_hd__a21oi_1 _1607_ (.A1(\MOS6502.IR[6] ),
    .A2(net72),
    .B1(net47),
    .Y(_0189_));
 sky130_fd_sc_hd__a31o_1 _1608_ (.A1(_0168_),
    .A2(_0188_),
    .A3(_0189_),
    .B1(net56),
    .X(_0190_));
 sky130_fd_sc_hd__a31o_1 _1609_ (.A1(\MOS6502.IR[5] ),
    .A2(net72),
    .A3(_0175_),
    .B1(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__o21a_1 _1610_ (.A1(\MOS6502.src_reg[0] ),
    .A2(net62),
    .B1(_0191_),
    .X(_0073_));
 sky130_fd_sc_hd__a22o_1 _1611_ (.A1(_0657_),
    .A2(_0169_),
    .B1(_0180_),
    .B2(_0165_),
    .X(_0192_));
 sky130_fd_sc_hd__o32a_1 _1612_ (.A1(_0170_),
    .A2(_0190_),
    .A3(_0192_),
    .B1(net62),
    .B2(\MOS6502.src_reg[1] ),
    .X(_0074_));
 sky130_fd_sc_hd__nor2_2 _1613_ (.A(_0614_),
    .B(_0679_),
    .Y(_0193_));
 sky130_fd_sc_hd__nand2_1 _1614_ (.A(net50),
    .B(_0604_),
    .Y(_0194_));
 sky130_fd_sc_hd__a32o_1 _1615_ (.A1(_0611_),
    .A2(_0614_),
    .A3(_0194_),
    .B1(_0193_),
    .B2(_0173_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _1616_ (.A0(\MOS6502.index_y ),
    .A1(_0195_),
    .S(net62),
    .X(_0075_));
 sky130_fd_sc_hd__o21a_1 _1617_ (.A1(_0611_),
    .A2(_0657_),
    .B1(_0169_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _1618_ (.A0(\MOS6502.store ),
    .A1(_0196_),
    .S(net62),
    .X(_0076_));
 sky130_fd_sc_hd__and2_1 _1619_ (.A(\MOS6502.write_back ),
    .B(net56),
    .X(_0197_));
 sky130_fd_sc_hd__a31o_1 _1620_ (.A1(net61),
    .A2(_0167_),
    .A3(_0193_),
    .B1(_0197_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _1621_ (.A0(\MOS6502.load_only ),
    .A1(_0171_),
    .S(net61),
    .X(_0078_));
 sky130_fd_sc_hd__a21o_1 _1622_ (.A1(\MOS6502.IR[5] ),
    .A2(_0193_),
    .B1(_0177_),
    .X(_0198_));
 sky130_fd_sc_hd__a22o_1 _1623_ (.A1(\MOS6502.inc ),
    .A2(net55),
    .B1(_0185_),
    .B2(_0198_),
    .X(_0079_));
 sky130_fd_sc_hd__nor3_1 _1624_ (.A(net52),
    .B(_0236_),
    .C(_0257_),
    .Y(_0199_));
 sky130_fd_sc_hd__a22o_1 _1625_ (.A1(\MOS6502.adc_sbc ),
    .A2(_0257_),
    .B1(_0611_),
    .B2(_0199_),
    .X(_0080_));
 sky130_fd_sc_hd__and4_1 _1626_ (.A(_0232_),
    .B(net62),
    .C(_0616_),
    .D(_0678_),
    .X(_0200_));
 sky130_fd_sc_hd__a21o_1 _1627_ (.A1(\MOS6502.shift ),
    .A2(net56),
    .B1(_0200_),
    .X(_0081_));
 sky130_fd_sc_hd__and3_1 _1628_ (.A(_0232_),
    .B(_0611_),
    .C(_0199_),
    .X(_0201_));
 sky130_fd_sc_hd__a22o_1 _1629_ (.A1(\MOS6502.adc_bcd ),
    .A2(_0257_),
    .B1(_0201_),
    .B2(\MOS6502.D ),
    .X(_0082_));
 sky130_fd_sc_hd__and3b_1 _1630_ (.A_N(net47),
    .B(_0615_),
    .C(net50),
    .X(_0202_));
 sky130_fd_sc_hd__a21o_1 _1631_ (.A1(net52),
    .A2(_0611_),
    .B1(_0202_),
    .X(_0203_));
 sky130_fd_sc_hd__a22o_1 _1632_ (.A1(\MOS6502.compare ),
    .A2(net55),
    .B1(_0185_),
    .B2(_0203_),
    .X(_0083_));
 sky130_fd_sc_hd__nor2_1 _1633_ (.A(_0628_),
    .B(_0679_),
    .Y(_0204_));
 sky130_fd_sc_hd__mux2_1 _1634_ (.A0(\MOS6502.shift_right ),
    .A1(_0204_),
    .S(net61),
    .X(_0084_));
 sky130_fd_sc_hd__a22o_1 _1635_ (.A1(\MOS6502.rotate ),
    .A2(net57),
    .B1(_0200_),
    .B2(\MOS6502.IR[5] ),
    .X(_0085_));
 sky130_fd_sc_hd__or4_1 _1636_ (.A(\MOS6502.IR[7] ),
    .B(\MOS6502.IR[5] ),
    .C(net56),
    .D(_0612_),
    .X(_0205_));
 sky130_fd_sc_hd__o211a_1 _1637_ (.A1(net52),
    .A2(_0236_),
    .B1(_0611_),
    .C1(_0232_),
    .X(_0206_));
 sky130_fd_sc_hd__o21a_1 _1638_ (.A1(\MOS6502.op[0] ),
    .A2(net61),
    .B1(_0205_),
    .X(_0086_));
 sky130_fd_sc_hd__a21o_1 _1639_ (.A1(net52),
    .A2(_0193_),
    .B1(_0202_),
    .X(_0207_));
 sky130_fd_sc_hd__o31a_1 _1640_ (.A1(_0611_),
    .A2(_0166_),
    .A3(_0207_),
    .B1(_0165_),
    .X(_0208_));
 sky130_fd_sc_hd__nor4_2 _1641_ (.A(net52),
    .B(_0614_),
    .C(net47),
    .D(_0663_),
    .Y(_0209_));
 sky130_fd_sc_hd__a31o_1 _1642_ (.A1(net50),
    .A2(_0635_),
    .A3(_0169_),
    .B1(_0204_),
    .X(_0210_));
 sky130_fd_sc_hd__or4_2 _1643_ (.A(_0206_),
    .B(_0208_),
    .C(_0209_),
    .D(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__nor2_1 _1644_ (.A(net55),
    .B(_0662_),
    .Y(_0212_));
 sky130_fd_sc_hd__a31o_1 _1645_ (.A1(_0232_),
    .A2(_0236_),
    .A3(_0678_),
    .B1(_0211_),
    .X(_0213_));
 sky130_fd_sc_hd__o2bb2a_1 _1646_ (.A1_N(_0211_),
    .A2_N(_0212_),
    .B1(\MOS6502.op[1] ),
    .B2(net61),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _1647_ (.A0(\MOS6502.op[2] ),
    .A1(_0211_),
    .S(net61),
    .X(_0088_));
 sky130_fd_sc_hd__nor2_1 _1648_ (.A(_0231_),
    .B(net55),
    .Y(_0214_));
 sky130_fd_sc_hd__a22o_1 _1649_ (.A1(\MOS6502.op[3] ),
    .A2(net55),
    .B1(_0213_),
    .B2(_0214_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _1650_ (.A0(\MOS6502.bit_ins ),
    .A1(_0209_),
    .S(net61),
    .X(_0090_));
 sky130_fd_sc_hd__a2bb2o_1 _1651_ (.A1_N(_0636_),
    .A2_N(_0174_),
    .B1(\MOS6502.clv ),
    .B2(net55),
    .X(_0091_));
 sky130_fd_sc_hd__and3_2 _1652_ (.A(\MOS6502.IR[5] ),
    .B(net72),
    .C(_0635_),
    .X(_0215_));
 sky130_fd_sc_hd__nor2_1 _1653_ (.A(net56),
    .B(_0628_),
    .Y(_0216_));
 sky130_fd_sc_hd__a22o_1 _1654_ (.A1(\MOS6502.sei ),
    .A2(net56),
    .B1(_0215_),
    .B2(_0216_),
    .X(_0092_));
 sky130_fd_sc_hd__and3_2 _1655_ (.A(net52),
    .B(_0601_),
    .C(_0635_),
    .X(_0217_));
 sky130_fd_sc_hd__a22o_1 _1656_ (.A1(\MOS6502.cli ),
    .A2(net56),
    .B1(_0216_),
    .B2(_0217_),
    .X(_0093_));
 sky130_fd_sc_hd__a22o_1 _1657_ (.A1(\MOS6502.sed ),
    .A2(net55),
    .B1(_0185_),
    .B2(_0215_),
    .X(_0094_));
 sky130_fd_sc_hd__a22o_1 _1658_ (.A1(\MOS6502.cld ),
    .A2(net55),
    .B1(_0185_),
    .B2(_0217_),
    .X(_0095_));
 sky130_fd_sc_hd__a22o_1 _1659_ (.A1(\MOS6502.sec ),
    .A2(net55),
    .B1(_0212_),
    .B2(_0215_),
    .X(_0096_));
 sky130_fd_sc_hd__a22o_1 _1660_ (.A1(\MOS6502.clc ),
    .A2(net55),
    .B1(_0212_),
    .B2(_0217_),
    .X(_0097_));
 sky130_fd_sc_hd__a22o_1 _1661_ (.A1(\MOS6502.php ),
    .A2(net57),
    .B1(_0637_),
    .B2(_0236_),
    .X(_0098_));
 sky130_fd_sc_hd__a22o_1 _1662_ (.A1(\MOS6502.plp ),
    .A2(net58),
    .B1(_0652_),
    .B2(_0236_),
    .X(_0099_));
 sky130_fd_sc_hd__or3b_1 _1663_ (.A(\MOS6502.NMI_edge ),
    .B(\MOS6502.NMI_1 ),
    .C_N(net10),
    .X(_0218_));
 sky130_fd_sc_hd__o21ai_1 _1664_ (.A1(_0221_),
    .A2(_0318_),
    .B1(_0218_),
    .Y(_0100_));
 sky130_fd_sc_hd__mux2_1 _1665_ (.A0(\MOS6502.ABH[0] ),
    .A1(net22),
    .S(net38),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _1666_ (.A0(\MOS6502.ABH[1] ),
    .A1(net23),
    .S(net38),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _1667_ (.A0(\MOS6502.ABH[2] ),
    .A1(net25),
    .S(net39),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _1668_ (.A0(\MOS6502.ABH[3] ),
    .A1(net26),
    .S(net39),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _1669_ (.A0(\MOS6502.ABH[4] ),
    .A1(net27),
    .S(net39),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _1670_ (.A0(\MOS6502.ABH[5] ),
    .A1(net28),
    .S(net39),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _1671_ (.A0(\MOS6502.ABH[6] ),
    .A1(net29),
    .S(net39),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _1672_ (.A0(\MOS6502.ABH[7] ),
    .A1(net30),
    .S(net39),
    .X(_0108_));
 sky130_fd_sc_hd__and3_4 _1673_ (.A(_0326_),
    .B(net44),
    .C(_0784_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _1674_ (.A0(\MOS6502.AXYS[3][0] ),
    .A1(_0786_),
    .S(_0219_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _1675_ (.A0(\MOS6502.AXYS[3][1] ),
    .A1(_0793_),
    .S(_0219_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _1676_ (.A0(\MOS6502.AXYS[3][2] ),
    .A1(_0798_),
    .S(_0219_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _1677_ (.A0(\MOS6502.AXYS[3][3] ),
    .A1(_0802_),
    .S(_0219_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _1678_ (.A0(\MOS6502.AXYS[3][4] ),
    .A1(_0803_),
    .S(_0219_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _1679_ (.A0(\MOS6502.AXYS[3][5] ),
    .A1(_0809_),
    .S(_0219_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _1680_ (.A0(\MOS6502.AXYS[3][6] ),
    .A1(_0814_),
    .S(_0219_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _1681_ (.A0(\MOS6502.AXYS[3][7] ),
    .A1(_0819_),
    .S(_0219_),
    .X(_0116_));
 sky130_fd_sc_hd__and2_4 _1682_ (.A(_0332_),
    .B(_0784_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _1683_ (.A0(\MOS6502.AXYS[0][0] ),
    .A1(_0786_),
    .S(_0220_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _1684_ (.A0(\MOS6502.AXYS[0][1] ),
    .A1(_0793_),
    .S(_0220_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _1685_ (.A0(\MOS6502.AXYS[0][2] ),
    .A1(_0798_),
    .S(_0220_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _1686_ (.A0(\MOS6502.AXYS[0][3] ),
    .A1(_0802_),
    .S(_0220_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _1687_ (.A0(\MOS6502.AXYS[0][4] ),
    .A1(_0803_),
    .S(_0220_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _1688_ (.A0(\MOS6502.AXYS[0][5] ),
    .A1(_0809_),
    .S(_0220_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _1689_ (.A0(\MOS6502.AXYS[0][6] ),
    .A1(_0814_),
    .S(_0220_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _1690_ (.A0(\MOS6502.AXYS[0][7] ),
    .A1(_0819_),
    .S(_0220_),
    .X(_0124_));
 sky130_fd_sc_hd__inv_2 _1691_ (.A(net11),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _1692_ (.A(net11),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _1693_ (.A(net11),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _1694_ (.A(net11),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _1695_ (.A(net11),
    .Y(_0029_));
 sky130_fd_sc_hd__dfrtp_1 _1696_ (.CLK(clknet_4_7_0_clk),
    .D(_0018_),
    .RESET_B(_0024_),
    .Q(\MOS6502.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1697_ (.CLK(clknet_4_7_0_clk),
    .D(_0019_),
    .RESET_B(_0025_),
    .Q(\MOS6502.state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _1698_ (.CLK(clknet_4_7_0_clk),
    .D(_0020_),
    .RESET_B(_0026_),
    .Q(\MOS6502.state[2] ));
 sky130_fd_sc_hd__dfstp_1 _1699_ (.CLK(clknet_4_7_0_clk),
    .D(_0021_),
    .SET_B(_0027_),
    .Q(\MOS6502.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1700_ (.CLK(clknet_4_7_0_clk),
    .D(_0022_),
    .RESET_B(_0028_),
    .Q(\MOS6502.state[4] ));
 sky130_fd_sc_hd__dfrtp_2 _1701_ (.CLK(clknet_4_13_0_clk),
    .D(_0023_),
    .RESET_B(_0029_),
    .Q(\MOS6502.state[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1702_ (.CLK(clknet_4_9_0_clk),
    .D(_0030_),
    .Q(\MOS6502.AXYS[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1703_ (.CLK(clknet_4_8_0_clk),
    .D(_0031_),
    .Q(\MOS6502.AXYS[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1704_ (.CLK(clknet_4_8_0_clk),
    .D(_0032_),
    .Q(\MOS6502.AXYS[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1705_ (.CLK(clknet_4_10_0_clk),
    .D(_0033_),
    .Q(\MOS6502.AXYS[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1706_ (.CLK(clknet_4_10_0_clk),
    .D(_0034_),
    .Q(\MOS6502.AXYS[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1707_ (.CLK(clknet_4_10_0_clk),
    .D(_0035_),
    .Q(\MOS6502.AXYS[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1708_ (.CLK(clknet_4_10_0_clk),
    .D(_0036_),
    .Q(\MOS6502.AXYS[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1709_ (.CLK(clknet_4_9_0_clk),
    .D(_0037_),
    .Q(\MOS6502.AXYS[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1710_ (.CLK(clknet_4_9_0_clk),
    .D(_0038_),
    .Q(\MOS6502.AXYS[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1711_ (.CLK(clknet_4_8_0_clk),
    .D(_0039_),
    .Q(\MOS6502.AXYS[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1712_ (.CLK(clknet_4_8_0_clk),
    .D(_0040_),
    .Q(\MOS6502.AXYS[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1713_ (.CLK(clknet_4_10_0_clk),
    .D(_0041_),
    .Q(\MOS6502.AXYS[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1714_ (.CLK(clknet_4_11_0_clk),
    .D(_0042_),
    .Q(\MOS6502.AXYS[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1715_ (.CLK(clknet_4_11_0_clk),
    .D(_0043_),
    .Q(\MOS6502.AXYS[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1716_ (.CLK(clknet_4_11_0_clk),
    .D(_0044_),
    .Q(\MOS6502.AXYS[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1717_ (.CLK(clknet_4_9_0_clk),
    .D(_0045_),
    .Q(\MOS6502.AXYS[1][7] ));
 sky130_fd_sc_hd__dfxtp_4 _1718_ (.CLK(clknet_4_2_0_clk),
    .D(_0001_),
    .Q(\MOS6502.ALU.CO ));
 sky130_fd_sc_hd__dfxtp_4 _1719_ (.CLK(clknet_4_0_0_clk),
    .D(\MOS6502.ALU.temp[7] ),
    .Q(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1720_ (.CLK(clknet_4_8_0_clk),
    .D(\MOS6502.ALU.temp_HC ),
    .Q(\MOS6502.ALU.HC ));
 sky130_fd_sc_hd__dfxtp_4 _1721_ (.CLK(clknet_4_3_0_clk),
    .D(\MOS6502.ALU.temp[0] ),
    .Q(\MOS6502.ADD[0] ));
 sky130_fd_sc_hd__dfxtp_4 _1722_ (.CLK(clknet_4_2_0_clk),
    .D(\MOS6502.ALU.temp[1] ),
    .Q(\MOS6502.ADD[1] ));
 sky130_fd_sc_hd__dfxtp_4 _1723_ (.CLK(clknet_4_8_0_clk),
    .D(\MOS6502.ALU.temp[2] ),
    .Q(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__dfxtp_4 _1724_ (.CLK(clknet_4_2_0_clk),
    .D(\MOS6502.ALU.temp[3] ),
    .Q(\MOS6502.ADD[3] ));
 sky130_fd_sc_hd__dfxtp_4 _1725_ (.CLK(clknet_4_8_0_clk),
    .D(\MOS6502.ALU.temp[4] ),
    .Q(\MOS6502.ADD[4] ));
 sky130_fd_sc_hd__dfxtp_4 _1726_ (.CLK(clknet_4_2_0_clk),
    .D(\MOS6502.ALU.temp[5] ),
    .Q(\MOS6502.ADD[5] ));
 sky130_fd_sc_hd__dfxtp_4 _1727_ (.CLK(clknet_4_2_0_clk),
    .D(\MOS6502.ALU.temp[6] ),
    .Q(\MOS6502.ADD[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1728_ (.CLK(clknet_4_0_0_clk),
    .D(\MOS6502.AI[7] ),
    .Q(\MOS6502.ALU.AI7 ));
 sky130_fd_sc_hd__dfxtp_1 _1729_ (.CLK(clknet_4_0_0_clk),
    .D(\MOS6502.ALU.temp_BI[7] ),
    .Q(\MOS6502.ALU.BI7 ));
 sky130_fd_sc_hd__dfxtp_2 _1730_ (.CLK(clknet_4_12_0_clk),
    .D(_0002_),
    .Q(\MOS6502.PC[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1731_ (.CLK(clknet_4_11_0_clk),
    .D(_0009_),
    .Q(\MOS6502.PC[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1732_ (.CLK(clknet_4_11_0_clk),
    .D(_0010_),
    .Q(\MOS6502.PC[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1733_ (.CLK(clknet_4_11_0_clk),
    .D(_0011_),
    .Q(\MOS6502.PC[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1734_ (.CLK(clknet_4_14_0_clk),
    .D(_0012_),
    .Q(\MOS6502.PC[4] ));
 sky130_fd_sc_hd__dfxtp_2 _1735_ (.CLK(clknet_4_14_0_clk),
    .D(_0013_),
    .Q(\MOS6502.PC[5] ));
 sky130_fd_sc_hd__dfxtp_2 _1736_ (.CLK(clknet_4_14_0_clk),
    .D(_0014_),
    .Q(\MOS6502.PC[6] ));
 sky130_fd_sc_hd__dfxtp_2 _1737_ (.CLK(clknet_4_12_0_clk),
    .D(_0015_),
    .Q(\MOS6502.PC[7] ));
 sky130_fd_sc_hd__dfxtp_2 _1738_ (.CLK(clknet_4_12_0_clk),
    .D(_0016_),
    .Q(\MOS6502.PC[8] ));
 sky130_fd_sc_hd__dfxtp_2 _1739_ (.CLK(clknet_4_12_0_clk),
    .D(_0017_),
    .Q(\MOS6502.PC[9] ));
 sky130_fd_sc_hd__dfxtp_2 _1740_ (.CLK(clknet_4_13_0_clk),
    .D(_0003_),
    .Q(\MOS6502.PC[10] ));
 sky130_fd_sc_hd__dfxtp_2 _1741_ (.CLK(clknet_4_13_0_clk),
    .D(_0004_),
    .Q(\MOS6502.PC[11] ));
 sky130_fd_sc_hd__dfxtp_2 _1742_ (.CLK(clknet_4_15_0_clk),
    .D(_0005_),
    .Q(\MOS6502.PC[12] ));
 sky130_fd_sc_hd__dfxtp_2 _1743_ (.CLK(clknet_4_15_0_clk),
    .D(_0006_),
    .Q(\MOS6502.PC[13] ));
 sky130_fd_sc_hd__dfxtp_2 _1744_ (.CLK(clknet_4_15_0_clk),
    .D(_0007_),
    .Q(\MOS6502.PC[14] ));
 sky130_fd_sc_hd__dfxtp_2 _1745_ (.CLK(clknet_4_13_0_clk),
    .D(_0008_),
    .Q(\MOS6502.PC[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1746_ (.CLK(clknet_4_11_0_clk),
    .D(_0046_),
    .Q(\MOS6502.ABL[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1747_ (.CLK(clknet_4_11_0_clk),
    .D(_0047_),
    .Q(\MOS6502.ABL[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1748_ (.CLK(clknet_4_14_0_clk),
    .D(_0048_),
    .Q(\MOS6502.ABL[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1749_ (.CLK(clknet_4_14_0_clk),
    .D(_0049_),
    .Q(\MOS6502.ABL[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1750_ (.CLK(clknet_4_14_0_clk),
    .D(_0050_),
    .Q(\MOS6502.ABL[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1751_ (.CLK(clknet_4_14_0_clk),
    .D(_0051_),
    .Q(\MOS6502.ABL[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1752_ (.CLK(clknet_4_14_0_clk),
    .D(_0052_),
    .Q(\MOS6502.ABL[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1753_ (.CLK(clknet_4_14_0_clk),
    .D(_0053_),
    .Q(\MOS6502.ABL[7] ));
 sky130_fd_sc_hd__dfxtp_2 _1754_ (.CLK(clknet_4_3_0_clk),
    .D(_0054_),
    .Q(\MOS6502.C ));
 sky130_fd_sc_hd__dfxtp_1 _1755_ (.CLK(clknet_4_9_0_clk),
    .D(_0000_),
    .Q(\MOS6502.adj_bcd ));
 sky130_fd_sc_hd__dfxtp_1 _1756_ (.CLK(clknet_4_12_0_clk),
    .D(net8),
    .Q(\MOS6502.backwards ));
 sky130_fd_sc_hd__dfxtp_1 _1757_ (.CLK(clknet_4_3_0_clk),
    .D(_0055_),
    .Q(\MOS6502.Z ));
 sky130_fd_sc_hd__dfxtp_1 _1758_ (.CLK(clknet_4_3_0_clk),
    .D(_0056_),
    .Q(\MOS6502.N ));
 sky130_fd_sc_hd__dfxtp_2 _1759_ (.CLK(clknet_4_3_0_clk),
    .D(_0057_),
    .Q(\MOS6502.D ));
 sky130_fd_sc_hd__dfxtp_2 _1760_ (.CLK(clknet_4_6_0_clk),
    .D(_0058_),
    .Q(\MOS6502.I ));
 sky130_fd_sc_hd__dfxtp_1 _1761_ (.CLK(clknet_4_3_0_clk),
    .D(_0059_),
    .Q(\MOS6502.V ));
 sky130_fd_sc_hd__dfxtp_1 _1762_ (.CLK(clknet_4_5_0_clk),
    .D(_0060_),
    .Q(\MOS6502.IRHOLD[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1763_ (.CLK(clknet_4_5_0_clk),
    .D(_0061_),
    .Q(\MOS6502.IRHOLD[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1764_ (.CLK(clknet_4_5_0_clk),
    .D(_0062_),
    .Q(\MOS6502.IRHOLD[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1765_ (.CLK(clknet_4_5_0_clk),
    .D(_0063_),
    .Q(\MOS6502.IRHOLD[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1766_ (.CLK(clknet_4_5_0_clk),
    .D(_0064_),
    .Q(\MOS6502.IRHOLD[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1767_ (.CLK(clknet_4_5_0_clk),
    .D(_0065_),
    .Q(\MOS6502.IRHOLD[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1768_ (.CLK(clknet_4_7_0_clk),
    .D(_0066_),
    .Q(\MOS6502.IRHOLD[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1769_ (.CLK(clknet_4_7_0_clk),
    .D(_0067_),
    .Q(\MOS6502.IRHOLD[7] ));
 sky130_fd_sc_hd__dfxtp_4 _1770_ (.CLK(clknet_4_13_0_clk),
    .D(_0068_),
    .Q(\MOS6502.IRHOLD_valid ));
 sky130_fd_sc_hd__dfxtp_1 _1771_ (.CLK(clknet_4_1_0_clk),
    .D(_0069_),
    .Q(\MOS6502.load_reg ));
 sky130_fd_sc_hd__dfxtp_1 _1772_ (.CLK(clknet_4_13_0_clk),
    .D(_0070_),
    .Q(\MOS6502.res ));
 sky130_fd_sc_hd__dfxtp_1 _1773_ (.CLK(clknet_4_6_0_clk),
    .D(_0071_),
    .Q(\MOS6502.dst_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1774_ (.CLK(clknet_4_1_0_clk),
    .D(_0072_),
    .Q(\MOS6502.dst_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1775_ (.CLK(clknet_4_4_0_clk),
    .D(_0073_),
    .Q(\MOS6502.src_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1776_ (.CLK(clknet_4_4_0_clk),
    .D(_0074_),
    .Q(\MOS6502.src_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1777_ (.CLK(clknet_4_4_0_clk),
    .D(_0075_),
    .Q(\MOS6502.index_y ));
 sky130_fd_sc_hd__dfxtp_2 _1778_ (.CLK(clknet_4_4_0_clk),
    .D(_0076_),
    .Q(\MOS6502.store ));
 sky130_fd_sc_hd__dfxtp_2 _1779_ (.CLK(clknet_4_1_0_clk),
    .D(_0077_),
    .Q(\MOS6502.write_back ));
 sky130_fd_sc_hd__dfxtp_2 _1780_ (.CLK(clknet_4_1_0_clk),
    .D(_0078_),
    .Q(\MOS6502.load_only ));
 sky130_fd_sc_hd__dfxtp_1 _1781_ (.CLK(clknet_4_1_0_clk),
    .D(_0079_),
    .Q(\MOS6502.inc ));
 sky130_fd_sc_hd__dfxtp_1 _1782_ (.CLK(clknet_4_1_0_clk),
    .D(_0080_),
    .Q(\MOS6502.adc_sbc ));
 sky130_fd_sc_hd__dfxtp_1 _1783_ (.CLK(clknet_4_3_0_clk),
    .D(_0081_),
    .Q(\MOS6502.shift ));
 sky130_fd_sc_hd__dfxtp_1 _1784_ (.CLK(clknet_4_2_0_clk),
    .D(_0082_),
    .Q(\MOS6502.adc_bcd ));
 sky130_fd_sc_hd__dfxtp_2 _1785_ (.CLK(clknet_4_1_0_clk),
    .D(_0083_),
    .Q(\MOS6502.compare ));
 sky130_fd_sc_hd__dfxtp_1 _1786_ (.CLK(clknet_4_0_0_clk),
    .D(_0084_),
    .Q(\MOS6502.shift_right ));
 sky130_fd_sc_hd__dfxtp_1 _1787_ (.CLK(clknet_4_6_0_clk),
    .D(_0085_),
    .Q(\MOS6502.rotate ));
 sky130_fd_sc_hd__dfxtp_1 _1788_ (.CLK(clknet_4_2_0_clk),
    .D(_0086_),
    .Q(\MOS6502.op[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1789_ (.CLK(clknet_4_0_0_clk),
    .D(_0087_),
    .Q(\MOS6502.op[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1790_ (.CLK(clknet_4_0_0_clk),
    .D(_0088_),
    .Q(\MOS6502.op[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1791_ (.CLK(clknet_4_0_0_clk),
    .D(_0089_),
    .Q(\MOS6502.op[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1792_ (.CLK(clknet_4_1_0_clk),
    .D(_0090_),
    .Q(\MOS6502.bit_ins ));
 sky130_fd_sc_hd__dfxtp_1 _1793_ (.CLK(clknet_4_1_0_clk),
    .D(_0091_),
    .Q(\MOS6502.clv ));
 sky130_fd_sc_hd__dfxtp_1 _1794_ (.CLK(clknet_4_4_0_clk),
    .D(_0092_),
    .Q(\MOS6502.sei ));
 sky130_fd_sc_hd__dfxtp_1 _1795_ (.CLK(clknet_4_6_0_clk),
    .D(_0093_),
    .Q(\MOS6502.cli ));
 sky130_fd_sc_hd__dfxtp_1 _1796_ (.CLK(clknet_4_1_0_clk),
    .D(_0094_),
    .Q(\MOS6502.sed ));
 sky130_fd_sc_hd__dfxtp_1 _1797_ (.CLK(clknet_4_0_0_clk),
    .D(_0095_),
    .Q(\MOS6502.cld ));
 sky130_fd_sc_hd__dfxtp_1 _1798_ (.CLK(clknet_4_3_0_clk),
    .D(_0096_),
    .Q(\MOS6502.sec ));
 sky130_fd_sc_hd__dfxtp_1 _1799_ (.CLK(clknet_4_1_0_clk),
    .D(_0097_),
    .Q(\MOS6502.clc ));
 sky130_fd_sc_hd__dfxtp_4 _1800_ (.CLK(clknet_4_6_0_clk),
    .D(_0098_),
    .Q(\MOS6502.php ));
 sky130_fd_sc_hd__dfxtp_1 _1801_ (.CLK(clknet_4_6_0_clk),
    .D(_0099_),
    .Q(\MOS6502.plp ));
 sky130_fd_sc_hd__dfxtp_1 _1802_ (.CLK(clknet_4_6_0_clk),
    .D(\MOS6502.IR[5] ),
    .Q(\MOS6502.cond_code[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1803_ (.CLK(clknet_4_3_0_clk),
    .D(\MOS6502.IR[6] ),
    .Q(\MOS6502.cond_code[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1804_ (.CLK(clknet_4_6_0_clk),
    .D(\MOS6502.IR[7] ),
    .Q(\MOS6502.cond_code[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1805_ (.CLK(clknet_4_13_0_clk),
    .D(net10),
    .Q(\MOS6502.NMI_1 ));
 sky130_fd_sc_hd__dfxtp_2 _1806_ (.CLK(clknet_4_13_0_clk),
    .D(_0100_),
    .Q(\MOS6502.NMI_edge ));
 sky130_fd_sc_hd__dfxtp_1 _1807_ (.CLK(clknet_4_12_0_clk),
    .D(_0101_),
    .Q(\MOS6502.ABH[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1808_ (.CLK(clknet_4_14_0_clk),
    .D(_0102_),
    .Q(\MOS6502.ABH[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1809_ (.CLK(clknet_4_15_0_clk),
    .D(_0103_),
    .Q(\MOS6502.ABH[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1810_ (.CLK(clknet_4_15_0_clk),
    .D(_0104_),
    .Q(\MOS6502.ABH[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1811_ (.CLK(clknet_4_15_0_clk),
    .D(_0105_),
    .Q(\MOS6502.ABH[4] ));
 sky130_fd_sc_hd__dfxtp_2 _1812_ (.CLK(clknet_4_15_0_clk),
    .D(_0106_),
    .Q(\MOS6502.ABH[5] ));
 sky130_fd_sc_hd__dfxtp_2 _1813_ (.CLK(clknet_4_15_0_clk),
    .D(_0107_),
    .Q(\MOS6502.ABH[6] ));
 sky130_fd_sc_hd__dfxtp_2 _1814_ (.CLK(clknet_4_15_0_clk),
    .D(_0108_),
    .Q(\MOS6502.ABH[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1815_ (.CLK(clknet_4_9_0_clk),
    .D(_0109_),
    .Q(\MOS6502.AXYS[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1816_ (.CLK(clknet_4_10_0_clk),
    .D(_0110_),
    .Q(\MOS6502.AXYS[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1817_ (.CLK(clknet_4_8_0_clk),
    .D(_0111_),
    .Q(\MOS6502.AXYS[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1818_ (.CLK(clknet_4_10_0_clk),
    .D(_0112_),
    .Q(\MOS6502.AXYS[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1819_ (.CLK(clknet_4_10_0_clk),
    .D(_0113_),
    .Q(\MOS6502.AXYS[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1820_ (.CLK(clknet_4_10_0_clk),
    .D(_0114_),
    .Q(\MOS6502.AXYS[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1821_ (.CLK(clknet_4_10_0_clk),
    .D(_0115_),
    .Q(\MOS6502.AXYS[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1822_ (.CLK(clknet_4_9_0_clk),
    .D(_0116_),
    .Q(\MOS6502.AXYS[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1823_ (.CLK(clknet_4_9_0_clk),
    .D(_0117_),
    .Q(\MOS6502.AXYS[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1824_ (.CLK(clknet_4_8_0_clk),
    .D(_0118_),
    .Q(\MOS6502.AXYS[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1825_ (.CLK(clknet_4_8_0_clk),
    .D(_0119_),
    .Q(\MOS6502.AXYS[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1826_ (.CLK(clknet_4_10_0_clk),
    .D(_0120_),
    .Q(\MOS6502.AXYS[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1827_ (.CLK(clknet_4_11_0_clk),
    .D(_0121_),
    .Q(\MOS6502.AXYS[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1828_ (.CLK(clknet_4_11_0_clk),
    .D(_0122_),
    .Q(\MOS6502.AXYS[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1829_ (.CLK(clknet_4_11_0_clk),
    .D(_0123_),
    .Q(\MOS6502.AXYS[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1830_ (.CLK(clknet_4_9_0_clk),
    .D(_0124_),
    .Q(\MOS6502.AXYS[0][7] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__buf_6 fanout38 (.A(_0127_),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 fanout39 (.A(_0127_),
    .X(net39));
 sky130_fd_sc_hd__buf_4 fanout40 (.A(_0732_),
    .X(net40));
 sky130_fd_sc_hd__buf_2 fanout41 (.A(_0732_),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(_0365_),
    .X(net42));
 sky130_fd_sc_hd__buf_6 fanout43 (.A(_0532_),
    .X(net43));
 sky130_fd_sc_hd__buf_12 fanout44 (.A(_0329_),
    .X(net44));
 sky130_fd_sc_hd__buf_6 fanout45 (.A(_0327_),
    .X(net45));
 sky130_fd_sc_hd__buf_4 fanout46 (.A(_0290_),
    .X(net46));
 sky130_fd_sc_hd__buf_4 fanout47 (.A(_0625_),
    .X(net47));
 sky130_fd_sc_hd__buf_4 fanout48 (.A(_0246_),
    .X(net48));
 sky130_fd_sc_hd__buf_6 fanout49 (.A(_0730_),
    .X(net49));
 sky130_fd_sc_hd__buf_4 fanout50 (.A(_0602_),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_8 fanout51 (.A(_0259_),
    .X(net51));
 sky130_fd_sc_hd__buf_6 fanout52 (.A(_0234_),
    .X(net52));
 sky130_fd_sc_hd__buf_4 fanout53 (.A(_0339_),
    .X(net53));
 sky130_fd_sc_hd__buf_2 fanout54 (.A(_0339_),
    .X(net54));
 sky130_fd_sc_hd__buf_4 fanout55 (.A(net57),
    .X(net55));
 sky130_fd_sc_hd__buf_2 fanout56 (.A(net57),
    .X(net56));
 sky130_fd_sc_hd__buf_4 fanout57 (.A(net60),
    .X(net57));
 sky130_fd_sc_hd__buf_4 fanout58 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__buf_2 fanout59 (.A(net60),
    .X(net59));
 sky130_fd_sc_hd__buf_6 fanout60 (.A(_0314_),
    .X(net60));
 sky130_fd_sc_hd__buf_4 fanout61 (.A(net63),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_8 fanout62 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__buf_4 fanout63 (.A(net64),
    .X(net63));
 sky130_fd_sc_hd__buf_12 fanout64 (.A(_0313_),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_8 fanout65 (.A(_0265_),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_8 fanout66 (.A(_0250_),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 fanout67 (.A(_0250_),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 fanout68 (.A(_0248_),
    .X(net68));
 sky130_fd_sc_hd__buf_6 fanout69 (.A(_0248_),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_16 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__buf_12 fanout71 (.A(_0230_),
    .X(net71));
 sky130_fd_sc_hd__buf_4 fanout72 (.A(_0600_),
    .X(net72));
 sky130_fd_sc_hd__buf_6 fanout73 (.A(_0251_),
    .X(net73));
 sky130_fd_sc_hd__buf_6 fanout74 (.A(_0251_),
    .X(net74));
 sky130_fd_sc_hd__buf_8 fanout75 (.A(net76),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_16 fanout76 (.A(_0242_),
    .X(net76));
 sky130_fd_sc_hd__buf_6 fanout77 (.A(net78),
    .X(net77));
 sky130_fd_sc_hd__buf_6 fanout78 (.A(_0237_),
    .X(net78));
 sky130_fd_sc_hd__buf_4 fanout79 (.A(\MOS6502.plp ),
    .X(net79));
 sky130_fd_sc_hd__buf_4 fanout80 (.A(\MOS6502.state[4] ),
    .X(net80));
 sky130_fd_sc_hd__buf_4 fanout81 (.A(\MOS6502.state[4] ),
    .X(net81));
 sky130_fd_sc_hd__buf_4 fanout82 (.A(net83),
    .X(net82));
 sky130_fd_sc_hd__buf_4 fanout83 (.A(\MOS6502.state[3] ),
    .X(net83));
 sky130_fd_sc_hd__buf_4 fanout84 (.A(net85),
    .X(net84));
 sky130_fd_sc_hd__buf_4 fanout85 (.A(\MOS6502.state[2] ),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_8 fanout86 (.A(\MOS6502.state[1] ),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 fanout87 (.A(\MOS6502.state[1] ),
    .X(net87));
 sky130_fd_sc_hd__buf_4 fanout88 (.A(net89),
    .X(net88));
 sky130_fd_sc_hd__buf_4 fanout89 (.A(\MOS6502.state[0] ),
    .X(net89));
 sky130_fd_sc_hd__buf_8 input1 (.A(io_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(io_in[9]),
    .X(net10));
 sky130_fd_sc_hd__buf_6 input11 (.A(rst),
    .X(net11));
 sky130_fd_sc_hd__buf_8 input2 (.A(io_in[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_6 input3 (.A(io_in[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_8 input4 (.A(io_in[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_6 input5 (.A(io_in[4]),
    .X(net5));
 sky130_fd_sc_hd__buf_6 input6 (.A(io_in[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_8 input7 (.A(io_in[6]),
    .X(net7));
 sky130_fd_sc_hd__buf_6 input8 (.A(io_in[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(io_in[8]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 output12 (.A(net12),
    .X(io_oeb));
 sky130_fd_sc_hd__buf_4 output13 (.A(net13),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_4 output14 (.A(net14),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_4 output15 (.A(net15),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_4 output16 (.A(net16),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_4 output17 (.A(net17),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_4 output18 (.A(net18),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_4 output19 (.A(net19),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_4 output20 (.A(net20),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_4 output21 (.A(net21),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_4 output22 (.A(net22),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_4 output23 (.A(net23),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_4 output24 (.A(net24),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_4 output25 (.A(net25),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_4 output26 (.A(net26),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_4 output27 (.A(net27),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_4 output28 (.A(net28),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_4 output29 (.A(net29),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_4 output30 (.A(net30),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_4 output31 (.A(net31),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_4 output32 (.A(net32),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_4 output33 (.A(net33),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_4 output34 (.A(net34),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_4 output35 (.A(net35),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_4 output36 (.A(net36),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_4 output37 (.A(net37),
    .X(io_out[7]));
 sky130_fd_sc_hd__conb_1 wrapped_6502_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 wrapped_6502_91 (.LO(net91));
 assign io_out[8] = net90;
 assign io_out[9] = net91;
endmodule

