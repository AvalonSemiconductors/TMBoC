magic
tech sky130B
magscale 1 2
timestamp 1677505267
<< nwell >>
rect 1066 41605 43922 42171
rect 1066 40517 43922 41083
rect 1066 39429 43922 39995
rect 1066 38341 43922 38907
rect 1066 37253 43922 37819
rect 1066 36165 43922 36731
rect 1066 35077 43922 35643
rect 1066 33989 43922 34555
rect 1066 32901 43922 33467
rect 1066 31813 43922 32379
rect 1066 30725 43922 31291
rect 1066 29637 43922 30203
rect 1066 28549 43922 29115
rect 1066 27461 43922 28027
rect 1066 26373 43922 26939
rect 1066 25285 43922 25851
rect 1066 24197 43922 24763
rect 1066 23109 43922 23675
rect 1066 22021 43922 22587
rect 1066 20933 43922 21499
rect 1066 19845 43922 20411
rect 1066 18757 43922 19323
rect 1066 17669 43922 18235
rect 1066 16581 43922 17147
rect 1066 15493 43922 16059
rect 1066 14405 43922 14971
rect 1066 13317 43922 13883
rect 1066 12229 43922 12795
rect 1066 11141 43922 11707
rect 1066 10053 43922 10619
rect 1066 8965 43922 9531
rect 1066 7877 43922 8443
rect 1066 6789 43922 7355
rect 1066 5701 43922 6267
rect 1066 4613 43922 5179
rect 1066 3525 43922 4091
rect 1066 2437 43922 3003
<< obsli1 >>
rect 1104 2159 43884 42449
<< obsm1 >>
rect 1104 2128 44054 44124
<< metal2 >>
rect 1278 44200 1390 45000
rect 2842 44200 2954 45000
rect 4406 44200 4518 45000
rect 5970 44200 6082 45000
rect 7534 44200 7646 45000
rect 9098 44200 9210 45000
rect 10662 44200 10774 45000
rect 12226 44200 12338 45000
rect 13790 44200 13902 45000
rect 15354 44200 15466 45000
rect 16918 44200 17030 45000
rect 18482 44200 18594 45000
rect 20046 44200 20158 45000
rect 21610 44200 21722 45000
rect 23174 44200 23286 45000
rect 24738 44200 24850 45000
rect 26302 44200 26414 45000
rect 27866 44200 27978 45000
rect 29430 44200 29542 45000
rect 30994 44200 31106 45000
rect 32558 44200 32670 45000
rect 34122 44200 34234 45000
rect 35686 44200 35798 45000
rect 37250 44200 37362 45000
rect 38814 44200 38926 45000
rect 40378 44200 40490 45000
rect 41942 44200 42054 45000
rect 43506 44200 43618 45000
<< obsm2 >>
rect 1446 44144 2786 44200
rect 3010 44144 4350 44200
rect 4574 44144 5914 44200
rect 6138 44144 7478 44200
rect 7702 44144 9042 44200
rect 9266 44144 10606 44200
rect 10830 44144 12170 44200
rect 12394 44144 13734 44200
rect 13958 44144 15298 44200
rect 15522 44144 16862 44200
rect 17086 44144 18426 44200
rect 18650 44144 19990 44200
rect 20214 44144 21554 44200
rect 21778 44144 23118 44200
rect 23342 44144 24682 44200
rect 24906 44144 26246 44200
rect 26470 44144 27810 44200
rect 28034 44144 29374 44200
rect 29598 44144 30938 44200
rect 31162 44144 32502 44200
rect 32726 44144 34066 44200
rect 34290 44144 35630 44200
rect 35854 44144 37194 44200
rect 37418 44144 38758 44200
rect 38982 44144 40322 44200
rect 40546 44144 41886 44200
rect 42110 44144 43450 44200
rect 43674 44144 44050 44200
rect 1308 2139 44050 44144
<< metal3 >>
rect 44200 42516 45000 42756
rect 44200 38844 45000 39084
rect 44200 35172 45000 35412
rect 44200 31500 45000 31740
rect 44200 27828 45000 28068
rect 44200 24156 45000 24396
rect 44200 20484 45000 20724
rect 44200 16812 45000 17052
rect 44200 13140 45000 13380
rect 44200 9468 45000 9708
rect 44200 5796 45000 6036
rect 44200 2124 45000 2364
<< obsm3 >>
rect 4210 42436 44120 42669
rect 4210 39164 44200 42436
rect 4210 38764 44120 39164
rect 4210 35492 44200 38764
rect 4210 35092 44120 35492
rect 4210 31820 44200 35092
rect 4210 31420 44120 31820
rect 4210 28148 44200 31420
rect 4210 27748 44120 28148
rect 4210 24476 44200 27748
rect 4210 24076 44120 24476
rect 4210 20804 44200 24076
rect 4210 20404 44120 20804
rect 4210 17132 44200 20404
rect 4210 16732 44120 17132
rect 4210 13460 44200 16732
rect 4210 13060 44120 13460
rect 4210 9788 44200 13060
rect 4210 9388 44120 9788
rect 4210 6116 44200 9388
rect 4210 5716 44120 6116
rect 4210 2444 44200 5716
rect 4210 2143 44120 2444
<< metal4 >>
rect 4208 2128 4528 42480
rect 19568 2128 19888 42480
rect 34928 2128 35248 42480
<< obsm4 >>
rect 24531 11323 34848 39949
rect 35328 11323 41341 39949
<< labels >>
rlabel metal3 s 44200 38844 45000 39084 6 clk
port 1 nsew signal input
rlabel metal3 s 44200 2124 45000 2364 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 44200 5796 45000 6036 6 io_in[1]
port 3 nsew signal input
rlabel metal3 s 44200 9468 45000 9708 6 io_in[2]
port 4 nsew signal input
rlabel metal3 s 44200 13140 45000 13380 6 io_in[3]
port 5 nsew signal input
rlabel metal3 s 44200 16812 45000 17052 6 io_in[4]
port 6 nsew signal input
rlabel metal3 s 44200 20484 45000 20724 6 io_in[5]
port 7 nsew signal input
rlabel metal3 s 44200 24156 45000 24396 6 io_in[6]
port 8 nsew signal input
rlabel metal3 s 44200 27828 45000 28068 6 io_in[7]
port 9 nsew signal input
rlabel metal3 s 44200 31500 45000 31740 6 io_in[8]
port 10 nsew signal input
rlabel metal3 s 44200 35172 45000 35412 6 io_in[9]
port 11 nsew signal input
rlabel metal2 s 43506 44200 43618 45000 6 io_oeb
port 12 nsew signal output
rlabel metal2 s 1278 44200 1390 45000 6 io_out[0]
port 13 nsew signal output
rlabel metal2 s 16918 44200 17030 45000 6 io_out[10]
port 14 nsew signal output
rlabel metal2 s 18482 44200 18594 45000 6 io_out[11]
port 15 nsew signal output
rlabel metal2 s 20046 44200 20158 45000 6 io_out[12]
port 16 nsew signal output
rlabel metal2 s 21610 44200 21722 45000 6 io_out[13]
port 17 nsew signal output
rlabel metal2 s 23174 44200 23286 45000 6 io_out[14]
port 18 nsew signal output
rlabel metal2 s 24738 44200 24850 45000 6 io_out[15]
port 19 nsew signal output
rlabel metal2 s 26302 44200 26414 45000 6 io_out[16]
port 20 nsew signal output
rlabel metal2 s 27866 44200 27978 45000 6 io_out[17]
port 21 nsew signal output
rlabel metal2 s 29430 44200 29542 45000 6 io_out[18]
port 22 nsew signal output
rlabel metal2 s 30994 44200 31106 45000 6 io_out[19]
port 23 nsew signal output
rlabel metal2 s 2842 44200 2954 45000 6 io_out[1]
port 24 nsew signal output
rlabel metal2 s 32558 44200 32670 45000 6 io_out[20]
port 25 nsew signal output
rlabel metal2 s 34122 44200 34234 45000 6 io_out[21]
port 26 nsew signal output
rlabel metal2 s 35686 44200 35798 45000 6 io_out[22]
port 27 nsew signal output
rlabel metal2 s 37250 44200 37362 45000 6 io_out[23]
port 28 nsew signal output
rlabel metal2 s 38814 44200 38926 45000 6 io_out[24]
port 29 nsew signal output
rlabel metal2 s 40378 44200 40490 45000 6 io_out[25]
port 30 nsew signal output
rlabel metal2 s 41942 44200 42054 45000 6 io_out[26]
port 31 nsew signal output
rlabel metal2 s 4406 44200 4518 45000 6 io_out[2]
port 32 nsew signal output
rlabel metal2 s 5970 44200 6082 45000 6 io_out[3]
port 33 nsew signal output
rlabel metal2 s 7534 44200 7646 45000 6 io_out[4]
port 34 nsew signal output
rlabel metal2 s 9098 44200 9210 45000 6 io_out[5]
port 35 nsew signal output
rlabel metal2 s 10662 44200 10774 45000 6 io_out[6]
port 36 nsew signal output
rlabel metal2 s 12226 44200 12338 45000 6 io_out[7]
port 37 nsew signal output
rlabel metal2 s 13790 44200 13902 45000 6 io_out[8]
port 38 nsew signal output
rlabel metal2 s 15354 44200 15466 45000 6 io_out[9]
port 39 nsew signal output
rlabel metal3 s 44200 42516 45000 42756 6 rst
port 40 nsew signal input
rlabel metal4 s 4208 2128 4528 42480 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 42480 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 42480 6 vssd1
port 42 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 45000 45000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4531764
string GDS_FILE /media/lucah/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/MOS6502/runs/23_02_27_14_37/results/signoff/wrapped_6502.magic.gds
string GDS_START 862696
<< end >>

